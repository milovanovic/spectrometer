// SPDX-License-Identifier: Apache-2.0

module AXI4StreamWidthAdapater_4_to_1(
  input         clock,
  input         reset,
  output        auto_in_ready,
  input         auto_in_valid,
  input  [7:0]  auto_in_bits_data,
  input         auto_in_bits_last,
  input         auto_out_ready,
  output        auto_out_valid,
  output [31:0] auto_out_bits_data,
  output        auto_out_bits_last
);
  reg [7:0] _T; // @[AXI4StreamWidthAdapter.scala 101:37]
  reg [31:0] _RAND_0;
  reg [7:0] _T_1; // @[AXI4StreamWidthAdapter.scala 101:37]
  reg [31:0] _RAND_1;
  reg [7:0] _T_2; // @[AXI4StreamWidthAdapter.scala 101:37]
  reg [31:0] _RAND_2;
  reg [1:0] _T_3; // @[AXI4StreamWidthAdapter.scala 102:22]
  reg [31:0] _RAND_3;
  wire  _T_4; // @[AXI4StreamWidthAdapter.scala 103:14]
  wire  _T_5; // @[AXI4StreamWidthAdapter.scala 103:38]
  wire [2:0] _T_6; // @[AXI4StreamWidthAdapter.scala 103:60]
  wire [2:0] _T_7; // @[AXI4StreamWidthAdapter.scala 103:33]
  wire [2:0] _GEN_0; // @[AXI4StreamWidthAdapter.scala 103:21]
  wire  _T_9; // @[AXI4StreamWidthAdapter.scala 106:29]
  wire  _T_10; // @[AXI4StreamWidthAdapter.scala 106:22]
  wire  _T_12; // @[AXI4StreamWidthAdapter.scala 106:29]
  wire  _T_13; // @[AXI4StreamWidthAdapter.scala 106:22]
  wire  _T_15; // @[AXI4StreamWidthAdapter.scala 106:29]
  wire  _T_16; // @[AXI4StreamWidthAdapter.scala 106:22]
  wire [23:0] _T_18; // @[Cat.scala 29:58]
  wire  ov0; // @[AXI4StreamWidthAdapter.scala 112:32]
  reg  _T_20; // @[AXI4StreamWidthAdapter.scala 101:37]
  reg [31:0] _RAND_4;
  reg  _T_21; // @[AXI4StreamWidthAdapter.scala 101:37]
  reg [31:0] _RAND_5;
  reg  _T_22; // @[AXI4StreamWidthAdapter.scala 101:37]
  reg [31:0] _RAND_6;
  reg [1:0] _T_23; // @[AXI4StreamWidthAdapter.scala 102:22]
  reg [31:0] _RAND_7;
  wire  _T_25; // @[AXI4StreamWidthAdapter.scala 103:38]
  wire [2:0] _T_26; // @[AXI4StreamWidthAdapter.scala 103:60]
  wire [2:0] _T_27; // @[AXI4StreamWidthAdapter.scala 103:33]
  wire [2:0] _GEN_4; // @[AXI4StreamWidthAdapter.scala 103:21]
  wire  _T_29; // @[AXI4StreamWidthAdapter.scala 106:29]
  wire  _T_30; // @[AXI4StreamWidthAdapter.scala 106:22]
  wire  _T_32; // @[AXI4StreamWidthAdapter.scala 106:29]
  wire  _T_33; // @[AXI4StreamWidthAdapter.scala 106:22]
  wire  _T_35; // @[AXI4StreamWidthAdapter.scala 106:29]
  wire  _T_36; // @[AXI4StreamWidthAdapter.scala 106:22]
  wire [3:0] _T_39; // @[Cat.scala 29:58]
  wire  ov1; // @[AXI4StreamWidthAdapter.scala 112:32]
  reg [1:0] _T_44; // @[AXI4StreamWidthAdapter.scala 102:22]
  reg [31:0] _RAND_8;
  wire  _T_46; // @[AXI4StreamWidthAdapter.scala 103:38]
  wire [2:0] _T_47; // @[AXI4StreamWidthAdapter.scala 103:60]
  wire [2:0] _T_48; // @[AXI4StreamWidthAdapter.scala 103:33]
  wire [2:0] _GEN_8; // @[AXI4StreamWidthAdapter.scala 103:21]
  wire  ov2; // @[AXI4StreamWidthAdapter.scala 112:32]
  reg [1:0] _T_64; // @[AXI4StreamWidthAdapter.scala 102:22]
  reg [31:0] _RAND_9;
  wire  _T_66; // @[AXI4StreamWidthAdapter.scala 103:38]
  wire [2:0] _T_67; // @[AXI4StreamWidthAdapter.scala 103:60]
  wire [2:0] _T_68; // @[AXI4StreamWidthAdapter.scala 103:33]
  wire [2:0] _GEN_12; // @[AXI4StreamWidthAdapter.scala 103:21]
  wire  ov3; // @[AXI4StreamWidthAdapter.scala 112:32]
  reg [1:0] _T_84; // @[AXI4StreamWidthAdapter.scala 102:22]
  reg [31:0] _RAND_10;
  wire  _T_86; // @[AXI4StreamWidthAdapter.scala 103:38]
  wire [2:0] _T_87; // @[AXI4StreamWidthAdapter.scala 103:60]
  wire [2:0] _T_88; // @[AXI4StreamWidthAdapter.scala 103:33]
  wire [2:0] _GEN_16; // @[AXI4StreamWidthAdapter.scala 103:21]
  wire  ov4; // @[AXI4StreamWidthAdapter.scala 112:32]
  wire  _T_101; // @[AXI4StreamWidthAdapter.scala 42:16]
  wire  _T_103; // @[AXI4StreamWidthAdapter.scala 42:11]
  wire  _T_104; // @[AXI4StreamWidthAdapter.scala 42:11]
  wire  _T_105; // @[AXI4StreamWidthAdapter.scala 43:16]
  wire  _T_107; // @[AXI4StreamWidthAdapter.scala 43:11]
  wire  _T_108; // @[AXI4StreamWidthAdapter.scala 43:11]
  wire  _T_109; // @[AXI4StreamWidthAdapter.scala 44:16]
  wire  _T_111; // @[AXI4StreamWidthAdapter.scala 44:11]
  wire  _T_112; // @[AXI4StreamWidthAdapter.scala 44:11]
  wire  _T_113; // @[AXI4StreamWidthAdapter.scala 45:16]
  wire  _T_115; // @[AXI4StreamWidthAdapter.scala 45:11]
  wire  _T_116; // @[AXI4StreamWidthAdapter.scala 45:11]
  assign _T_4 = auto_in_valid & auto_out_ready; // @[AXI4StreamWidthAdapter.scala 103:14]
  assign _T_5 = _T_3 == 2'h3; // @[AXI4StreamWidthAdapter.scala 103:38]
  assign _T_6 = _T_3 + 2'h1; // @[AXI4StreamWidthAdapter.scala 103:60]
  assign _T_7 = _T_5 ? 3'h0 : _T_6; // @[AXI4StreamWidthAdapter.scala 103:33]
  assign _GEN_0 = _T_4 ? _T_7 : {{1'd0}, _T_3}; // @[AXI4StreamWidthAdapter.scala 103:21]
  assign _T_9 = _T_3 == 2'h0; // @[AXI4StreamWidthAdapter.scala 106:29]
  assign _T_10 = _T_4 & _T_9; // @[AXI4StreamWidthAdapter.scala 106:22]
  assign _T_12 = _T_3 == 2'h1; // @[AXI4StreamWidthAdapter.scala 106:29]
  assign _T_13 = _T_4 & _T_12; // @[AXI4StreamWidthAdapter.scala 106:22]
  assign _T_15 = _T_3 == 2'h2; // @[AXI4StreamWidthAdapter.scala 106:29]
  assign _T_16 = _T_4 & _T_15; // @[AXI4StreamWidthAdapter.scala 106:22]
  assign _T_18 = {auto_in_bits_data,_T_2,_T_1}; // @[Cat.scala 29:58]
  assign ov0 = _T_5 & auto_in_valid; // @[AXI4StreamWidthAdapter.scala 112:32]
  assign _T_25 = _T_23 == 2'h3; // @[AXI4StreamWidthAdapter.scala 103:38]
  assign _T_26 = _T_23 + 2'h1; // @[AXI4StreamWidthAdapter.scala 103:60]
  assign _T_27 = _T_25 ? 3'h0 : _T_26; // @[AXI4StreamWidthAdapter.scala 103:33]
  assign _GEN_4 = _T_4 ? _T_27 : {{1'd0}, _T_23}; // @[AXI4StreamWidthAdapter.scala 103:21]
  assign _T_29 = _T_23 == 2'h0; // @[AXI4StreamWidthAdapter.scala 106:29]
  assign _T_30 = _T_4 & _T_29; // @[AXI4StreamWidthAdapter.scala 106:22]
  assign _T_32 = _T_23 == 2'h1; // @[AXI4StreamWidthAdapter.scala 106:29]
  assign _T_33 = _T_4 & _T_32; // @[AXI4StreamWidthAdapter.scala 106:22]
  assign _T_35 = _T_23 == 2'h2; // @[AXI4StreamWidthAdapter.scala 106:29]
  assign _T_36 = _T_4 & _T_35; // @[AXI4StreamWidthAdapter.scala 106:22]
  assign _T_39 = {auto_in_bits_last,_T_22,_T_21,_T_20}; // @[Cat.scala 29:58]
  assign ov1 = _T_25 & auto_in_valid; // @[AXI4StreamWidthAdapter.scala 112:32]
  assign _T_46 = _T_44 == 2'h3; // @[AXI4StreamWidthAdapter.scala 103:38]
  assign _T_47 = _T_44 + 2'h1; // @[AXI4StreamWidthAdapter.scala 103:60]
  assign _T_48 = _T_46 ? 3'h0 : _T_47; // @[AXI4StreamWidthAdapter.scala 103:33]
  assign _GEN_8 = _T_4 ? _T_48 : {{1'd0}, _T_44}; // @[AXI4StreamWidthAdapter.scala 103:21]
  assign ov2 = _T_46 & auto_in_valid; // @[AXI4StreamWidthAdapter.scala 112:32]
  assign _T_66 = _T_64 == 2'h3; // @[AXI4StreamWidthAdapter.scala 103:38]
  assign _T_67 = _T_64 + 2'h1; // @[AXI4StreamWidthAdapter.scala 103:60]
  assign _T_68 = _T_66 ? 3'h0 : _T_67; // @[AXI4StreamWidthAdapter.scala 103:33]
  assign _GEN_12 = _T_4 ? _T_68 : {{1'd0}, _T_64}; // @[AXI4StreamWidthAdapter.scala 103:21]
  assign ov3 = _T_66 & auto_in_valid; // @[AXI4StreamWidthAdapter.scala 112:32]
  assign _T_86 = _T_84 == 2'h3; // @[AXI4StreamWidthAdapter.scala 103:38]
  assign _T_87 = _T_84 + 2'h1; // @[AXI4StreamWidthAdapter.scala 103:60]
  assign _T_88 = _T_86 ? 3'h0 : _T_87; // @[AXI4StreamWidthAdapter.scala 103:33]
  assign _GEN_16 = _T_4 ? _T_88 : {{1'd0}, _T_84}; // @[AXI4StreamWidthAdapter.scala 103:21]
  assign ov4 = _T_86 & auto_in_valid; // @[AXI4StreamWidthAdapter.scala 112:32]
  assign _T_101 = ov0 == ov1; // @[AXI4StreamWidthAdapter.scala 42:16]
  assign _T_103 = _T_101 | reset; // @[AXI4StreamWidthAdapter.scala 42:11]
  assign _T_104 = ~_T_103; // @[AXI4StreamWidthAdapter.scala 42:11]
  assign _T_105 = ov0 == ov2; // @[AXI4StreamWidthAdapter.scala 43:16]
  assign _T_107 = _T_105 | reset; // @[AXI4StreamWidthAdapter.scala 43:11]
  assign _T_108 = ~_T_107; // @[AXI4StreamWidthAdapter.scala 43:11]
  assign _T_109 = ov0 == ov3; // @[AXI4StreamWidthAdapter.scala 44:16]
  assign _T_111 = _T_109 | reset; // @[AXI4StreamWidthAdapter.scala 44:11]
  assign _T_112 = ~_T_111; // @[AXI4StreamWidthAdapter.scala 44:11]
  assign _T_113 = ov0 == ov4; // @[AXI4StreamWidthAdapter.scala 45:16]
  assign _T_115 = _T_113 | reset; // @[AXI4StreamWidthAdapter.scala 45:11]
  assign _T_116 = ~_T_115; // @[AXI4StreamWidthAdapter.scala 45:11]
  assign auto_in_ready = auto_out_ready; // @[LazyModule.scala 173:31]
  assign auto_out_valid = _T_5 & auto_in_valid; // @[LazyModule.scala 173:49]
  assign auto_out_bits_data = {_T_18,_T}; // @[LazyModule.scala 173:49]
  assign auto_out_bits_last = _T_39 != 4'h0; // @[LazyModule.scala 173:49]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T = _RAND_0[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1 = _RAND_1[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_2 = _RAND_2[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_3 = _RAND_3[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_20 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_21 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_22 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_23 = _RAND_7[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_44 = _RAND_8[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_64 = _RAND_9[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_84 = _RAND_10[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (_T_10) begin
      _T <= auto_in_bits_data;
    end
    if (_T_13) begin
      _T_1 <= auto_in_bits_data;
    end
    if (_T_16) begin
      _T_2 <= auto_in_bits_data;
    end
    if (reset) begin
      _T_3 <= 2'h0;
    end else begin
      _T_3 <= _GEN_0[1:0];
    end
    if (_T_30) begin
      _T_20 <= auto_in_bits_last;
    end
    if (_T_33) begin
      _T_21 <= auto_in_bits_last;
    end
    if (_T_36) begin
      _T_22 <= auto_in_bits_last;
    end
    if (reset) begin
      _T_23 <= 2'h0;
    end else begin
      _T_23 <= _GEN_4[1:0];
    end
    if (reset) begin
      _T_44 <= 2'h0;
    end else begin
      _T_44 <= _GEN_8[1:0];
    end
    if (reset) begin
      _T_64 <= 2'h0;
    end else begin
      _T_64 <= _GEN_12[1:0];
    end
    if (reset) begin
      _T_84 <= 2'h0;
    end else begin
      _T_84 <= _GEN_16[1:0];
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_104) begin
          $fwrite(32'h80000002,"Assertion failed\n    at AXI4StreamWidthAdapter.scala:42 assert(ov0 === ov1)\n"); // @[AXI4StreamWidthAdapter.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_104) begin
          $fatal; // @[AXI4StreamWidthAdapter.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_108) begin
          $fwrite(32'h80000002,"Assertion failed\n    at AXI4StreamWidthAdapter.scala:43 assert(ov0 === ov2)\n"); // @[AXI4StreamWidthAdapter.scala 43:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_108) begin
          $fatal; // @[AXI4StreamWidthAdapter.scala 43:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_112) begin
          $fwrite(32'h80000002,"Assertion failed\n    at AXI4StreamWidthAdapter.scala:44 assert(ov0 === ov3)\n"); // @[AXI4StreamWidthAdapter.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_112) begin
          $fatal; // @[AXI4StreamWidthAdapter.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_116) begin
          $fwrite(32'h80000002,"Assertion failed\n    at AXI4StreamWidthAdapter.scala:45 assert(ov0 === ov4)\n"); // @[AXI4StreamWidthAdapter.scala 45:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_116) begin
          $fatal; // @[AXI4StreamWidthAdapter.scala 45:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module Queue(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input         io_enq_bits_read,
  input  [31:0] io_enq_bits_data,
  input         io_enq_bits_extra,
  input         io_deq_ready,
  output        io_deq_valid,
  output        io_deq_bits_read,
  output [31:0] io_deq_bits_data,
  output        io_deq_bits_extra
);
  reg  _T_read [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_0;
  wire  _T_read__T_18_data; // @[Decoupled.scala 209:24]
  wire  _T_read__T_18_addr; // @[Decoupled.scala 209:24]
  wire  _T_read__T_10_data; // @[Decoupled.scala 209:24]
  wire  _T_read__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T_read__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T_read__T_10_en; // @[Decoupled.scala 209:24]
  reg [31:0] _T_data [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_1;
  wire [31:0] _T_data__T_18_data; // @[Decoupled.scala 209:24]
  wire  _T_data__T_18_addr; // @[Decoupled.scala 209:24]
  wire [31:0] _T_data__T_10_data; // @[Decoupled.scala 209:24]
  wire  _T_data__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T_data__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T_data__T_10_en; // @[Decoupled.scala 209:24]
  reg  _T_extra [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_2;
  wire  _T_extra__T_18_data; // @[Decoupled.scala 209:24]
  wire  _T_extra__T_18_addr; // @[Decoupled.scala 209:24]
  wire  _T_extra__T_10_data; // @[Decoupled.scala 209:24]
  wire  _T_extra__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T_extra__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T_extra__T_10_en; // @[Decoupled.scala 209:24]
  reg  value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_3;
  reg  value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_4;
  reg  _T_1; // @[Decoupled.scala 212:35]
  reg [31:0] _RAND_5;
  wire  _T_2; // @[Decoupled.scala 214:41]
  wire  _T_3; // @[Decoupled.scala 215:36]
  wire  _T_4; // @[Decoupled.scala 215:33]
  wire  _T_5; // @[Decoupled.scala 216:32]
  wire  _T_6; // @[Decoupled.scala 40:37]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _T_12; // @[Counter.scala 39:22]
  wire  _T_14; // @[Counter.scala 39:22]
  wire  _T_15; // @[Decoupled.scala 227:16]
  assign _T_read__T_18_addr = value_1;
  assign _T_read__T_18_data = _T_read[_T_read__T_18_addr]; // @[Decoupled.scala 209:24]
  assign _T_read__T_10_data = io_enq_bits_read;
  assign _T_read__T_10_addr = value;
  assign _T_read__T_10_mask = 1'h1;
  assign _T_read__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_data__T_18_addr = value_1;
  assign _T_data__T_18_data = _T_data[_T_data__T_18_addr]; // @[Decoupled.scala 209:24]
  assign _T_data__T_10_data = io_enq_bits_data;
  assign _T_data__T_10_addr = value;
  assign _T_data__T_10_mask = 1'h1;
  assign _T_data__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_extra__T_18_addr = value_1;
  assign _T_extra__T_18_data = _T_extra[_T_extra__T_18_addr]; // @[Decoupled.scala 209:24]
  assign _T_extra__T_10_data = io_enq_bits_extra;
  assign _T_extra__T_10_addr = value;
  assign _T_extra__T_10_mask = 1'h1;
  assign _T_extra__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_2 = value == value_1; // @[Decoupled.scala 214:41]
  assign _T_3 = ~_T_1; // @[Decoupled.scala 215:36]
  assign _T_4 = _T_2 & _T_3; // @[Decoupled.scala 215:33]
  assign _T_5 = _T_2 & _T_1; // @[Decoupled.scala 216:32]
  assign _T_6 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  assign _T_8 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  assign _T_12 = value + 1'h1; // @[Counter.scala 39:22]
  assign _T_14 = value_1 + 1'h1; // @[Counter.scala 39:22]
  assign _T_15 = _T_6 != _T_8; // @[Decoupled.scala 227:16]
  assign io_enq_ready = ~_T_5; // @[Decoupled.scala 232:16]
  assign io_deq_valid = ~_T_4; // @[Decoupled.scala 231:16]
  assign io_deq_bits_read = _T_read__T_18_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_data = _T_data__T_18_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_extra = _T_extra__T_18_data; // @[Decoupled.scala 233:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_read[initvar] = _RAND_0[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_data[initvar] = _RAND_1[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_extra[initvar] = _RAND_2[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  value = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  value_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_1 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T_read__T_10_en & _T_read__T_10_mask) begin
      _T_read[_T_read__T_10_addr] <= _T_read__T_10_data; // @[Decoupled.scala 209:24]
    end
    if(_T_data__T_10_en & _T_data__T_10_mask) begin
      _T_data[_T_data__T_10_addr] <= _T_data__T_10_data; // @[Decoupled.scala 209:24]
    end
    if(_T_extra__T_10_en & _T_extra__T_10_mask) begin
      _T_extra[_T_extra__T_10_addr] <= _T_extra__T_10_data; // @[Decoupled.scala 209:24]
    end
    if (reset) begin
      value <= 1'h0;
    end else if (_T_6) begin
      value <= _T_12;
    end
    if (reset) begin
      value_1 <= 1'h0;
    end else if (_T_8) begin
      value_1 <= _T_14;
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else if (_T_15) begin
      _T_1 <= _T_6;
    end
  end
endmodule
module AXI4Splitter(
  input         clock,
  input         reset,
  output        auto_mem_in_aw_ready,
  input         auto_mem_in_aw_valid,
  input         auto_mem_in_aw_bits_id,
  input  [29:0] auto_mem_in_aw_bits_addr,
  output        auto_mem_in_w_ready,
  input         auto_mem_in_w_valid,
  input  [31:0] auto_mem_in_w_bits_data,
  input  [3:0]  auto_mem_in_w_bits_strb,
  input         auto_mem_in_b_ready,
  output        auto_mem_in_b_valid,
  output        auto_mem_in_b_bits_id,
  output        auto_mem_in_ar_ready,
  input         auto_mem_in_ar_valid,
  input         auto_mem_in_ar_bits_id,
  input  [29:0] auto_mem_in_ar_bits_addr,
  input  [2:0]  auto_mem_in_ar_bits_size,
  input         auto_mem_in_r_ready,
  output        auto_mem_in_r_valid,
  output        auto_mem_in_r_bits_id,
  output [31:0] auto_mem_in_r_bits_data,
  output        auto_stream_in_ready,
  input         auto_stream_in_valid,
  input  [31:0] auto_stream_in_bits_data,
  input         auto_stream_in_bits_last,
  input         auto_stream_out_4_ready,
  output        auto_stream_out_4_valid,
  output [31:0] auto_stream_out_4_bits_data,
  output        auto_stream_out_4_bits_last,
  input         auto_stream_out_3_ready,
  output        auto_stream_out_3_valid,
  output [31:0] auto_stream_out_3_bits_data,
  output        auto_stream_out_3_bits_last,
  input         auto_stream_out_2_ready,
  output        auto_stream_out_2_valid,
  output [31:0] auto_stream_out_2_bits_data,
  output        auto_stream_out_2_bits_last,
  input         auto_stream_out_1_ready,
  output        auto_stream_out_1_valid,
  output [31:0] auto_stream_out_1_bits_data,
  output        auto_stream_out_1_bits_last,
  input         auto_stream_out_0_ready,
  output        auto_stream_out_0_valid,
  output [31:0] auto_stream_out_0_bits_data,
  output        auto_stream_out_0_bits_last
);
  wire  Queue_clock; // @[Decoupled.scala 287:21]
  wire  Queue_reset; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_read; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_enq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_extra; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_read; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_deq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_extra; // @[Decoupled.scala 287:21]
  reg [31:0] ctrlReg; // @[Splitter.scala 27:26]
  reg [31:0] _RAND_0;
  reg [31:0] maskReg; // @[Splitter.scala 28:26]
  reg [31:0] _RAND_1;
  wire  _T_7; // @[RegisterRouter.scala 40:39]
  wire  _T_8; // @[RegisterRouter.scala 40:26]
  wire  _T_9; // @[RegisterRouter.scala 42:29]
  wire  _T_52_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 290:17]
  wire [29:0] _T_16; // @[RegisterRouter.scala 48:19]
  wire [1:0] _T_56; // @[RegisterRouter.scala 59:16]
  wire  _T_58; // @[RegisterRouter.scala 59:16]
  wire  _T_10; // @[RegisterRouter.scala 42:26]
  wire [1:0] _T_19; // @[OneHot.scala 65:12]
  wire [1:0] _T_21; // @[Misc.scala 200:81]
  wire  _T_22; // @[Misc.scala 204:21]
  wire  _T_25; // @[Misc.scala 209:20]
  wire  _T_27; // @[Misc.scala 213:38]
  wire  _T_28; // @[Misc.scala 213:29]
  wire  _T_30; // @[Misc.scala 213:38]
  wire  _T_31; // @[Misc.scala 213:29]
  wire  _T_34; // @[Misc.scala 209:20]
  wire  _T_35; // @[Misc.scala 212:27]
  wire  _T_36; // @[Misc.scala 213:38]
  wire  _T_37; // @[Misc.scala 213:29]
  wire  _T_38; // @[Misc.scala 212:27]
  wire  _T_39; // @[Misc.scala 213:38]
  wire  _T_40; // @[Misc.scala 213:29]
  wire  _T_41; // @[Misc.scala 212:27]
  wire  _T_42; // @[Misc.scala 213:38]
  wire  _T_43; // @[Misc.scala 213:29]
  wire  _T_44; // @[Misc.scala 212:27]
  wire  _T_45; // @[Misc.scala 213:38]
  wire  _T_46; // @[Misc.scala 213:29]
  wire [3:0] _T_49; // @[Cat.scala 29:58]
  wire [3:0] _T_51; // @[RegisterRouter.scala 54:25]
  wire [7:0] _T_70; // @[Bitwise.scala 72:12]
  wire [7:0] _T_72; // @[Bitwise.scala 72:12]
  wire [7:0] _T_74; // @[Bitwise.scala 72:12]
  wire [7:0] _T_76; // @[Bitwise.scala 72:12]
  wire [31:0] _T_79; // @[Cat.scala 29:58]
  wire  _T_98; // @[RegisterRouter.scala 59:16]
  wire  _T_151; // @[RegisterRouter.scala 59:16]
  wire [1:0] _T_145; // @[OneHot.scala 58:35]
  wire  _T_168; // @[RegisterRouter.scala 59:16]
  wire  _T_175; // @[RegisterRouter.scala 59:16]
  wire  _T_176; // @[RegisterRouter.scala 59:16]
  wire  _T_105; // @[RegisterRouter.scala 59:16]
  wire  _T_170; // @[RegisterRouter.scala 59:16]
  wire  _T_171; // @[RegisterRouter.scala 59:16]
  wire  _T_128; // @[RegisterRouter.scala 59:16]
  wire  _GEN_11; // @[MuxLiteral.scala 48:10]
  wire [31:0] _GEN_13; // @[MuxLiteral.scala 48:10]
  wire  _T_226_bits_read; // @[Decoupled.scala 308:19 Decoupled.scala 309:14]
  wire  _T_226_valid; // @[Decoupled.scala 308:19 Decoupled.scala 310:15]
  wire  _T_229; // @[RegisterRouter.scala 65:29]
  wire  _T_232; // @[Splitter.scala 45:34]
  wire  _T_233; // @[Splitter.scala 45:34]
  wire  _T_234; // @[Splitter.scala 45:34]
  wire  readyOR; // @[Splitter.scala 45:34]
  wire  _T_235; // @[Splitter.scala 46:34]
  wire  _T_236; // @[Splitter.scala 46:34]
  wire  _T_237; // @[Splitter.scala 46:34]
  wire  readyAND; // @[Splitter.scala 46:34]
  wire  _T_238; // @[Splitter.scala 49:19]
  wire  _T_239; // @[Splitter.scala 52:24]
  wire  _GEN_14; // @[Splitter.scala 52:33]
  wire  _T_242; // @[Splitter.scala 62:34]
  wire  _T_246; // @[Splitter.scala 62:34]
  wire  _T_250; // @[Splitter.scala 62:34]
  wire  _T_254; // @[Splitter.scala 62:34]
  wire  _T_258; // @[Splitter.scala 62:34]
  Queue Queue ( // @[Decoupled.scala 287:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_read(Queue_io_enq_bits_read),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_extra(Queue_io_enq_bits_extra),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_read(Queue_io_deq_bits_read),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_extra(Queue_io_deq_bits_extra)
  );
  assign _T_7 = auto_mem_in_aw_valid & auto_mem_in_w_valid; // @[RegisterRouter.scala 40:39]
  assign _T_8 = auto_mem_in_ar_valid | _T_7; // @[RegisterRouter.scala 40:26]
  assign _T_9 = ~auto_mem_in_ar_valid; // @[RegisterRouter.scala 42:29]
  assign _T_52_ready = Queue_io_enq_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 290:17]
  assign _T_16 = auto_mem_in_ar_valid ? auto_mem_in_ar_bits_addr : auto_mem_in_aw_bits_addr; // @[RegisterRouter.scala 48:19]
  assign _T_56 = _T_16[3:2] & 2'h2; // @[RegisterRouter.scala 59:16]
  assign _T_58 = _T_56 == 2'h0; // @[RegisterRouter.scala 59:16]
  assign _T_10 = _T_52_ready & _T_9; // @[RegisterRouter.scala 42:26]
  assign _T_19 = 2'h1 << auto_mem_in_ar_bits_size[0]; // @[OneHot.scala 65:12]
  assign _T_21 = _T_19 | 2'h1; // @[Misc.scala 200:81]
  assign _T_22 = auto_mem_in_ar_bits_size >= 3'h2; // @[Misc.scala 204:21]
  assign _T_25 = ~auto_mem_in_ar_bits_addr[1]; // @[Misc.scala 209:20]
  assign _T_27 = _T_21[1] & _T_25; // @[Misc.scala 213:38]
  assign _T_28 = _T_22 | _T_27; // @[Misc.scala 213:29]
  assign _T_30 = _T_21[1] & auto_mem_in_ar_bits_addr[1]; // @[Misc.scala 213:38]
  assign _T_31 = _T_22 | _T_30; // @[Misc.scala 213:29]
  assign _T_34 = ~auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 209:20]
  assign _T_35 = _T_25 & _T_34; // @[Misc.scala 212:27]
  assign _T_36 = _T_21[0] & _T_35; // @[Misc.scala 213:38]
  assign _T_37 = _T_28 | _T_36; // @[Misc.scala 213:29]
  assign _T_38 = _T_25 & auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  assign _T_39 = _T_21[0] & _T_38; // @[Misc.scala 213:38]
  assign _T_40 = _T_28 | _T_39; // @[Misc.scala 213:29]
  assign _T_41 = auto_mem_in_ar_bits_addr[1] & _T_34; // @[Misc.scala 212:27]
  assign _T_42 = _T_21[0] & _T_41; // @[Misc.scala 213:38]
  assign _T_43 = _T_31 | _T_42; // @[Misc.scala 213:29]
  assign _T_44 = auto_mem_in_ar_bits_addr[1] & auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  assign _T_45 = _T_21[0] & _T_44; // @[Misc.scala 213:38]
  assign _T_46 = _T_31 | _T_45; // @[Misc.scala 213:29]
  assign _T_49 = {_T_46,_T_43,_T_40,_T_37}; // @[Cat.scala 29:58]
  assign _T_51 = auto_mem_in_ar_valid ? _T_49 : auto_mem_in_w_bits_strb; // @[RegisterRouter.scala 54:25]
  assign _T_70 = _T_51[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_72 = _T_51[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_74 = _T_51[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_76 = _T_51[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_79 = {_T_76,_T_74,_T_72,_T_70}; // @[Cat.scala 29:58]
  assign _T_98 = _T_79 == 32'hffffffff; // @[RegisterRouter.scala 59:16]
  assign _T_151 = _T_8 & _T_52_ready; // @[RegisterRouter.scala 59:16]
  assign _T_145 = 2'h1 << _T_16[2]; // @[OneHot.scala 58:35]
  assign _T_168 = _T_151 & _T_9; // @[RegisterRouter.scala 59:16]
  assign _T_175 = _T_168 & _T_145[1]; // @[RegisterRouter.scala 59:16]
  assign _T_176 = _T_175 & _T_58; // @[RegisterRouter.scala 59:16]
  assign _T_105 = _T_176 & _T_98; // @[RegisterRouter.scala 59:16]
  assign _T_170 = _T_168 & _T_145[0]; // @[RegisterRouter.scala 59:16]
  assign _T_171 = _T_170 & _T_58; // @[RegisterRouter.scala 59:16]
  assign _T_128 = _T_171 & _T_98; // @[RegisterRouter.scala 59:16]
  assign _GEN_11 = _T_16[2] ? _T_58 : _T_58; // @[MuxLiteral.scala 48:10]
  assign _GEN_13 = _T_16[2] ? maskReg : ctrlReg; // @[MuxLiteral.scala 48:10]
  assign _T_226_bits_read = Queue_io_deq_bits_read; // @[Decoupled.scala 308:19 Decoupled.scala 309:14]
  assign _T_226_valid = Queue_io_deq_valid; // @[Decoupled.scala 308:19 Decoupled.scala 310:15]
  assign _T_229 = ~_T_226_bits_read; // @[RegisterRouter.scala 65:29]
  assign _T_232 = auto_stream_out_0_ready | auto_stream_out_1_ready; // @[Splitter.scala 45:34]
  assign _T_233 = _T_232 | auto_stream_out_2_ready; // @[Splitter.scala 45:34]
  assign _T_234 = _T_233 | auto_stream_out_3_ready; // @[Splitter.scala 45:34]
  assign readyOR = _T_234 | auto_stream_out_4_ready; // @[Splitter.scala 45:34]
  assign _T_235 = auto_stream_out_0_ready & auto_stream_out_1_ready; // @[Splitter.scala 46:34]
  assign _T_236 = _T_235 & auto_stream_out_2_ready; // @[Splitter.scala 46:34]
  assign _T_237 = _T_236 & auto_stream_out_3_ready; // @[Splitter.scala 46:34]
  assign readyAND = _T_237 & auto_stream_out_4_ready; // @[Splitter.scala 46:34]
  assign _T_238 = ctrlReg == 32'h0; // @[Splitter.scala 49:19]
  assign _T_239 = ctrlReg == 32'h1; // @[Splitter.scala 52:24]
  assign _GEN_14 = _T_239 & readyOR; // @[Splitter.scala 52:33]
  assign _T_242 = ~maskReg[0]; // @[Splitter.scala 62:34]
  assign _T_246 = ~maskReg[1]; // @[Splitter.scala 62:34]
  assign _T_250 = ~maskReg[2]; // @[Splitter.scala 62:34]
  assign _T_254 = ~maskReg[3]; // @[Splitter.scala 62:34]
  assign _T_258 = ~maskReg[4]; // @[Splitter.scala 62:34]
  assign auto_mem_in_aw_ready = _T_10 & auto_mem_in_w_valid; // @[LazyModule.scala 173:31]
  assign auto_mem_in_w_ready = _T_10 & auto_mem_in_aw_valid; // @[LazyModule.scala 173:31]
  assign auto_mem_in_b_valid = _T_226_valid & _T_229; // @[LazyModule.scala 173:31]
  assign auto_mem_in_b_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_mem_in_ar_ready = Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_valid = _T_226_valid & _T_226_bits_read; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 173:31]
  assign auto_stream_in_ready = _T_238 ? readyAND : _GEN_14; // @[LazyModule.scala 173:31]
  assign auto_stream_out_4_valid = auto_stream_in_valid & _T_258; // @[LazyModule.scala 173:49]
  assign auto_stream_out_4_bits_data = auto_stream_in_bits_data; // @[LazyModule.scala 173:49]
  assign auto_stream_out_4_bits_last = auto_stream_in_bits_last; // @[LazyModule.scala 173:49]
  assign auto_stream_out_3_valid = auto_stream_in_valid & _T_254; // @[LazyModule.scala 173:49]
  assign auto_stream_out_3_bits_data = auto_stream_in_bits_data; // @[LazyModule.scala 173:49]
  assign auto_stream_out_3_bits_last = auto_stream_in_bits_last; // @[LazyModule.scala 173:49]
  assign auto_stream_out_2_valid = auto_stream_in_valid & _T_250; // @[LazyModule.scala 173:49]
  assign auto_stream_out_2_bits_data = auto_stream_in_bits_data; // @[LazyModule.scala 173:49]
  assign auto_stream_out_2_bits_last = auto_stream_in_bits_last; // @[LazyModule.scala 173:49]
  assign auto_stream_out_1_valid = auto_stream_in_valid & _T_246; // @[LazyModule.scala 173:49]
  assign auto_stream_out_1_bits_data = auto_stream_in_bits_data; // @[LazyModule.scala 173:49]
  assign auto_stream_out_1_bits_last = auto_stream_in_bits_last; // @[LazyModule.scala 173:49]
  assign auto_stream_out_0_valid = auto_stream_in_valid & _T_242; // @[LazyModule.scala 173:49]
  assign auto_stream_out_0_bits_data = auto_stream_in_bits_data; // @[LazyModule.scala 173:49]
  assign auto_stream_out_0_bits_last = auto_stream_in_bits_last; // @[LazyModule.scala 173:49]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_mem_in_ar_valid | _T_7; // @[Decoupled.scala 288:22]
  assign Queue_io_enq_bits_read = auto_mem_in_ar_valid; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_data = _GEN_11 ? _GEN_13 : 32'h0; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_extra = auto_mem_in_ar_valid ? auto_mem_in_ar_bits_id : auto_mem_in_aw_bits_id; // @[Decoupled.scala 289:21]
  assign Queue_io_deq_ready = _T_226_bits_read ? auto_mem_in_r_ready : auto_mem_in_b_ready; // @[Decoupled.scala 311:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ctrlReg = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  maskReg = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      ctrlReg <= 32'h0;
    end else if (_T_128) begin
      ctrlReg <= auto_mem_in_w_bits_data;
    end
    if (reset) begin
      maskReg <= 32'h0;
    end else if (_T_105) begin
      maskReg <= auto_mem_in_w_bits_data;
    end
  end
endmodule
module Queue_1(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input  [7:0] io_enq_bits_data,
  input        io_enq_bits_last,
  input        io_deq_ready,
  output       io_deq_valid,
  output [7:0] io_deq_bits_data,
  output       io_deq_bits_last
);
  reg [7:0] _T_data [0:0]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_0;
  wire [7:0] _T_data__T_14_data; // @[Decoupled.scala 209:24]
  wire  _T_data__T_14_addr; // @[Decoupled.scala 209:24]
  wire [7:0] _T_data__T_10_data; // @[Decoupled.scala 209:24]
  wire  _T_data__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T_data__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T_data__T_10_en; // @[Decoupled.scala 209:24]
  reg  _T_last [0:0]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_1;
  wire  _T_last__T_14_data; // @[Decoupled.scala 209:24]
  wire  _T_last__T_14_addr; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_data; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_en; // @[Decoupled.scala 209:24]
  reg  _T_1; // @[Decoupled.scala 212:35]
  reg [31:0] _RAND_2;
  wire  _T_3; // @[Decoupled.scala 215:36]
  wire  _T_6; // @[Decoupled.scala 40:37]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[Decoupled.scala 240:27]
  wire  _GEN_22; // @[Decoupled.scala 237:18]
  wire  _GEN_21; // @[Decoupled.scala 237:18]
  wire  _T_11; // @[Decoupled.scala 227:16]
  wire  _T_12; // @[Decoupled.scala 231:19]
  assign _T_data__T_14_addr = 1'h0;
  assign _T_data__T_14_data = _T_data[_T_data__T_14_addr]; // @[Decoupled.scala 209:24]
  assign _T_data__T_10_data = io_enq_bits_data;
  assign _T_data__T_10_addr = 1'h0;
  assign _T_data__T_10_mask = 1'h1;
  assign _T_data__T_10_en = _T_3 ? _GEN_13 : _T_6;
  assign _T_last__T_14_addr = 1'h0;
  assign _T_last__T_14_data = _T_last[_T_last__T_14_addr]; // @[Decoupled.scala 209:24]
  assign _T_last__T_10_data = io_enq_bits_last;
  assign _T_last__T_10_addr = 1'h0;
  assign _T_last__T_10_mask = 1'h1;
  assign _T_last__T_10_en = _T_3 ? _GEN_13 : _T_6;
  assign _T_3 = ~_T_1; // @[Decoupled.scala 215:36]
  assign _T_6 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  assign _T_8 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = io_deq_ready ? 1'h0 : _T_6; // @[Decoupled.scala 240:27]
  assign _GEN_22 = _T_3 ? _GEN_13 : _T_6; // @[Decoupled.scala 237:18]
  assign _GEN_21 = _T_3 ? 1'h0 : _T_8; // @[Decoupled.scala 237:18]
  assign _T_11 = _GEN_22 != _GEN_21; // @[Decoupled.scala 227:16]
  assign _T_12 = ~_T_3; // @[Decoupled.scala 231:19]
  assign io_enq_ready = io_deq_ready | _T_3; // @[Decoupled.scala 232:16 Decoupled.scala 245:40]
  assign io_deq_valid = io_enq_valid | _T_12; // @[Decoupled.scala 231:16 Decoupled.scala 236:40]
  assign io_deq_bits_data = _T_3 ? io_enq_bits_data : _T_data__T_14_data; // @[Decoupled.scala 233:15 Decoupled.scala 238:19]
  assign io_deq_bits_last = _T_3 ? io_enq_bits_last : _T_last__T_14_data; // @[Decoupled.scala 233:15 Decoupled.scala 238:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_data[initvar] = _RAND_0[7:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_last[initvar] = _RAND_1[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_1 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T_data__T_10_en & _T_data__T_10_mask) begin
      _T_data[_T_data__T_10_addr] <= _T_data__T_10_data; // @[Decoupled.scala 209:24]
    end
    if(_T_last__T_10_en & _T_last__T_10_mask) begin
      _T_last[_T_last__T_10_addr] <= _T_last__T_10_data; // @[Decoupled.scala 209:24]
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else if (_T_11) begin
      if (_T_3) begin
        if (io_deq_ready) begin
          _T_1 <= 1'h0;
        end else begin
          _T_1 <= _T_6;
        end
      end else begin
        _T_1 <= _T_6;
      end
    end
  end
endmodule
module StreamBuffer(
  input        clock,
  input        reset,
  input        auto_out_out_ready,
  output       auto_out_out_valid,
  output [7:0] auto_out_out_bits_data,
  output       auto_out_out_bits_last,
  output       auto_in_in_ready,
  input        auto_in_in_valid,
  input  [7:0] auto_in_in_bits_data,
  input        auto_in_in_bits_last
);
  wire  Queue_clock; // @[Decoupled.scala 287:21]
  wire  Queue_reset; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 287:21]
  wire [7:0] Queue_io_enq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_last; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 287:21]
  wire [7:0] Queue_io_deq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_last; // @[Decoupled.scala 287:21]
  Queue_1 Queue ( // @[Decoupled.scala 287:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_last(Queue_io_enq_bits_last),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_last(Queue_io_deq_bits_last)
  );
  assign auto_out_out_valid = Queue_io_deq_valid; // @[LazyModule.scala 173:49]
  assign auto_out_out_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_out_bits_last = Queue_io_deq_bits_last; // @[LazyModule.scala 173:49]
  assign auto_in_in_ready = Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_in_in_valid; // @[Decoupled.scala 288:22]
  assign Queue_io_enq_bits_data = auto_in_in_bits_data; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_last = auto_in_in_bits_last; // @[Decoupled.scala 289:21]
  assign Queue_io_deq_ready = auto_out_out_ready; // @[Decoupled.scala 311:15]
endmodule
module QueueCompatibility(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input  [1:0] io_enq_bits,
  input        io_deq_ready,
  output       io_deq_valid,
  output [1:0] io_deq_bits
);
  reg [1:0] _T [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_0;
  wire [1:0] _T__T_18_data; // @[Decoupled.scala 209:24]
  wire  _T__T_18_addr; // @[Decoupled.scala 209:24]
  wire [1:0] _T__T_10_data; // @[Decoupled.scala 209:24]
  wire  _T__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T__T_10_en; // @[Decoupled.scala 209:24]
  reg  value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_1;
  reg  value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_2;
  reg  _T_1; // @[Decoupled.scala 212:35]
  reg [31:0] _RAND_3;
  wire  _T_2; // @[Decoupled.scala 214:41]
  wire  _T_3; // @[Decoupled.scala 215:36]
  wire  _T_4; // @[Decoupled.scala 215:33]
  wire  _T_5; // @[Decoupled.scala 216:32]
  wire  _T_6; // @[Decoupled.scala 40:37]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _T_12; // @[Counter.scala 39:22]
  wire  _GEN_9; // @[Decoupled.scala 240:27]
  wire  _GEN_12; // @[Decoupled.scala 237:18]
  wire  _T_14; // @[Counter.scala 39:22]
  wire  _GEN_11; // @[Decoupled.scala 237:18]
  wire  _T_15; // @[Decoupled.scala 227:16]
  wire  _T_16; // @[Decoupled.scala 231:19]
  assign _T__T_18_addr = value_1;
  assign _T__T_18_data = _T[_T__T_18_addr]; // @[Decoupled.scala 209:24]
  assign _T__T_10_data = io_enq_bits;
  assign _T__T_10_addr = value;
  assign _T__T_10_mask = 1'h1;
  assign _T__T_10_en = _T_4 ? _GEN_9 : _T_6;
  assign _T_2 = value == value_1; // @[Decoupled.scala 214:41]
  assign _T_3 = ~_T_1; // @[Decoupled.scala 215:36]
  assign _T_4 = _T_2 & _T_3; // @[Decoupled.scala 215:33]
  assign _T_5 = _T_2 & _T_1; // @[Decoupled.scala 216:32]
  assign _T_6 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  assign _T_8 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  assign _T_12 = value + 1'h1; // @[Counter.scala 39:22]
  assign _GEN_9 = io_deq_ready ? 1'h0 : _T_6; // @[Decoupled.scala 240:27]
  assign _GEN_12 = _T_4 ? _GEN_9 : _T_6; // @[Decoupled.scala 237:18]
  assign _T_14 = value_1 + 1'h1; // @[Counter.scala 39:22]
  assign _GEN_11 = _T_4 ? 1'h0 : _T_8; // @[Decoupled.scala 237:18]
  assign _T_15 = _GEN_12 != _GEN_11; // @[Decoupled.scala 227:16]
  assign _T_16 = ~_T_4; // @[Decoupled.scala 231:19]
  assign io_enq_ready = ~_T_5; // @[Decoupled.scala 232:16]
  assign io_deq_valid = io_enq_valid | _T_16; // @[Decoupled.scala 231:16 Decoupled.scala 236:40]
  assign io_deq_bits = _T_4 ? io_enq_bits : _T__T_18_data; // @[Decoupled.scala 233:15 Decoupled.scala 238:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T[initvar] = _RAND_0[1:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  value = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  value_1 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_1 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T__T_10_en & _T__T_10_mask) begin
      _T[_T__T_10_addr] <= _T__T_10_data; // @[Decoupled.scala 209:24]
    end
    if (reset) begin
      value <= 1'h0;
    end else if (_GEN_12) begin
      value <= _T_12;
    end
    if (reset) begin
      value_1 <= 1'h0;
    end else if (_GEN_11) begin
      value_1 <= _T_14;
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else if (_T_15) begin
      if (_T_4) begin
        if (io_deq_ready) begin
          _T_1 <= 1'h0;
        end else begin
          _T_1 <= _T_6;
        end
      end else begin
        _T_1 <= _T_6;
      end
    end
  end
endmodule
module AXI4Xbar(
  input         clock,
  input         reset,
  output        auto_in_aw_ready,
  input         auto_in_aw_valid,
  input         auto_in_aw_bits_id,
  input  [29:0] auto_in_aw_bits_addr,
  output        auto_in_w_ready,
  input         auto_in_w_valid,
  input  [31:0] auto_in_w_bits_data,
  input  [3:0]  auto_in_w_bits_strb,
  input         auto_in_w_bits_last,
  input         auto_in_b_ready,
  output        auto_in_b_valid,
  output [1:0]  auto_in_b_bits_resp,
  output        auto_in_ar_ready,
  input         auto_in_ar_valid,
  input         auto_in_ar_bits_id,
  input  [29:0] auto_in_ar_bits_addr,
  input  [2:0]  auto_in_ar_bits_size,
  input         auto_in_r_ready,
  output        auto_in_r_valid,
  output [31:0] auto_in_r_bits_data,
  output [1:0]  auto_in_r_bits_resp,
  output        auto_in_r_bits_last,
  input         auto_out_1_aw_ready,
  output        auto_out_1_aw_valid,
  output        auto_out_1_aw_bits_id,
  output [29:0] auto_out_1_aw_bits_addr,
  input         auto_out_1_w_ready,
  output        auto_out_1_w_valid,
  output [31:0] auto_out_1_w_bits_data,
  output [3:0]  auto_out_1_w_bits_strb,
  output        auto_out_1_b_ready,
  input         auto_out_1_b_valid,
  input         auto_out_1_b_bits_id,
  input         auto_out_1_ar_ready,
  output        auto_out_1_ar_valid,
  output        auto_out_1_ar_bits_id,
  output [29:0] auto_out_1_ar_bits_addr,
  output [2:0]  auto_out_1_ar_bits_size,
  output        auto_out_1_r_ready,
  input         auto_out_1_r_valid,
  input         auto_out_1_r_bits_id,
  input  [31:0] auto_out_1_r_bits_data,
  input         auto_out_0_aw_ready,
  output        auto_out_0_aw_valid,
  output [29:0] auto_out_0_aw_bits_addr,
  input         auto_out_0_w_ready,
  output        auto_out_0_w_valid,
  output [31:0] auto_out_0_w_bits_data,
  output        auto_out_0_b_ready,
  input         auto_out_0_b_valid
);
  wire  awIn_0_clock; // @[Xbar.scala 55:47]
  wire  awIn_0_reset; // @[Xbar.scala 55:47]
  wire  awIn_0_io_enq_ready; // @[Xbar.scala 55:47]
  wire  awIn_0_io_enq_valid; // @[Xbar.scala 55:47]
  wire [1:0] awIn_0_io_enq_bits; // @[Xbar.scala 55:47]
  wire  awIn_0_io_deq_ready; // @[Xbar.scala 55:47]
  wire  awIn_0_io_deq_valid; // @[Xbar.scala 55:47]
  wire [1:0] awIn_0_io_deq_bits; // @[Xbar.scala 55:47]
  wire [30:0] _T_1; // @[Parameters.scala 137:49]
  wire [30:0] _T_3; // @[Parameters.scala 137:52]
  wire  requestARIO_0_0; // @[Parameters.scala 137:67]
  wire [29:0] _T_5; // @[Parameters.scala 137:31]
  wire [30:0] _T_6; // @[Parameters.scala 137:49]
  wire [30:0] _T_8; // @[Parameters.scala 137:52]
  wire  requestARIO_0_1; // @[Parameters.scala 137:67]
  wire [30:0] _T_11; // @[Parameters.scala 137:49]
  wire [30:0] _T_13; // @[Parameters.scala 137:52]
  wire  requestAWIO_0_0; // @[Parameters.scala 137:67]
  wire [29:0] _T_15; // @[Parameters.scala 137:31]
  wire [30:0] _T_16; // @[Parameters.scala 137:49]
  wire [30:0] _T_18; // @[Parameters.scala 137:52]
  wire  requestAWIO_0_1; // @[Parameters.scala 137:67]
  wire  requestROI_1_0; // @[Parameters.scala 47:9]
  wire  requestBOI_1_0; // @[Parameters.scala 47:9]
  wire [1:0] _T_20; // @[Xbar.scala 64:75]
  wire  requestWIO_0_0; // @[Xbar.scala 65:73]
  wire  requestWIO_0_1; // @[Xbar.scala 65:73]
  wire [1:0] _T_27; // @[Xbar.scala 93:45]
  wire  in_0_ar_ready; // @[Mux.scala 27:72]
  reg [2:0] _T_36; // @[Xbar.scala 104:34]
  reg [31:0] _RAND_0;
  wire  _T_55; // @[Xbar.scala 112:22]
  reg  _T_37; // @[Xbar.scala 105:29]
  reg [31:0] _RAND_1;
  wire  _T_54; // @[Xbar.scala 111:75]
  wire  _T_56; // @[Xbar.scala 112:34]
  wire  _T_57; // @[Xbar.scala 112:80]
  wire  _T_59; // @[Xbar.scala 112:48]
  wire  io_in_0_ar_ready; // @[Xbar.scala 130:45]
  wire  _T_31; // @[Decoupled.scala 40:37]
  reg  _T_222; // @[Xbar.scala 242:23]
  reg [31:0] _RAND_2;
  wire  _T_129; // @[Xbar.scala 222:40]
  reg  _T_278_1; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_3;
  wire  _T_285; // @[Mux.scala 27:72]
  wire  in_0_r_valid; // @[Xbar.scala 278:22]
  wire  _T_33; // @[Decoupled.scala 40:37]
  wire [1:0] _T_224; // @[Cat.scala 29:58]
  reg [1:0] _T_231; // @[Arbiter.scala 20:23]
  reg [31:0] _RAND_4;
  wire [1:0] _T_232; // @[Arbiter.scala 21:30]
  wire [1:0] _T_233; // @[Arbiter.scala 21:28]
  wire [3:0] _T_234; // @[Cat.scala 29:58]
  wire [3:0] _GEN_18; // @[package.scala 208:43]
  wire [3:0] _T_236; // @[package.scala 208:43]
  wire [3:0] _T_239; // @[Arbiter.scala 22:66]
  wire [3:0] _GEN_19; // @[Arbiter.scala 22:58]
  wire [3:0] _T_240; // @[Arbiter.scala 22:58]
  wire [1:0] _T_243; // @[Arbiter.scala 23:39]
  wire [1:0] _T_244; // @[Arbiter.scala 23:18]
  wire  _T_257; // @[Xbar.scala 250:63]
  wire  _T_279_1; // @[Xbar.scala 262:23]
  wire [35:0] _T_295; // @[Mux.scala 27:72]
  wire [35:0] _T_296; // @[Mux.scala 27:72]
  wire  in_0_r_bits_last; // @[Mux.scala 27:72]
  wire  _T_35; // @[Xbar.scala 120:45]
  wire [2:0] _GEN_20; // @[Xbar.scala 106:30]
  wire [2:0] _T_39; // @[Xbar.scala 106:30]
  wire [2:0] _GEN_21; // @[Xbar.scala 106:48]
  wire [2:0] _T_41; // @[Xbar.scala 106:48]
  wire  _T_42; // @[Xbar.scala 107:23]
  wire  _T_43; // @[Xbar.scala 107:43]
  wire  _T_44; // @[Xbar.scala 107:34]
  wire  _T_46; // @[Xbar.scala 107:22]
  wire  _T_47; // @[Xbar.scala 107:22]
  wire  _T_48; // @[Xbar.scala 108:23]
  wire  _T_50; // @[Xbar.scala 108:34]
  wire  _T_52; // @[Xbar.scala 108:22]
  wire  _T_53; // @[Xbar.scala 108:22]
  wire  _T_115; // @[Mux.scala 27:72]
  wire  _T_116; // @[Mux.scala 27:72]
  wire  in_0_aw_ready; // @[Mux.scala 27:72]
  reg  _T_90; // @[Xbar.scala 137:30]
  reg [31:0] _RAND_5;
  wire  _T_94; // @[Xbar.scala 139:57]
  wire  _T_95; // @[Xbar.scala 139:45]
  reg [2:0] _T_64; // @[Xbar.scala 104:34]
  reg [31:0] _RAND_6;
  wire  _T_83; // @[Xbar.scala 112:22]
  reg  _T_65; // @[Xbar.scala 105:29]
  reg [31:0] _RAND_7;
  wire  _T_82; // @[Xbar.scala 111:75]
  wire  _T_84; // @[Xbar.scala 112:34]
  wire  _T_85; // @[Xbar.scala 112:80]
  wire  _T_87; // @[Xbar.scala 112:48]
  wire  io_in_0_aw_ready; // @[Xbar.scala 139:82]
  wire  _T_60; // @[Decoupled.scala 40:37]
  reg  _T_304; // @[Xbar.scala 242:23]
  reg [31:0] _RAND_8;
  wire  _T_133; // @[Xbar.scala 222:40]
  wire  _T_305; // @[Xbar.scala 246:36]
  reg  _T_360_0; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_9;
  wire  _T_366; // @[Mux.scala 27:72]
  reg  _T_360_1; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_10;
  wire  _T_367; // @[Mux.scala 27:72]
  wire  _T_368; // @[Mux.scala 27:72]
  wire  in_0_b_valid; // @[Xbar.scala 278:22]
  wire  _T_62; // @[Decoupled.scala 40:37]
  wire [2:0] _GEN_22; // @[Xbar.scala 106:30]
  wire [2:0] _T_67; // @[Xbar.scala 106:30]
  wire [2:0] _GEN_23; // @[Xbar.scala 106:48]
  wire [2:0] _T_69; // @[Xbar.scala 106:48]
  wire  _T_70; // @[Xbar.scala 107:23]
  wire  _T_71; // @[Xbar.scala 107:43]
  wire  _T_72; // @[Xbar.scala 107:34]
  wire  _T_74; // @[Xbar.scala 107:22]
  wire  _T_75; // @[Xbar.scala 107:22]
  wire  _T_76; // @[Xbar.scala 108:23]
  wire  _T_78; // @[Xbar.scala 108:34]
  wire  _T_80; // @[Xbar.scala 108:22]
  wire  _T_81; // @[Xbar.scala 108:22]
  wire  in_0_ar_valid; // @[Xbar.scala 129:45]
  wire  _T_92; // @[Xbar.scala 138:45]
  wire  in_0_aw_valid; // @[Xbar.scala 138:82]
  wire  _T_97; // @[Xbar.scala 140:54]
  wire  _T_99; // @[Decoupled.scala 40:37]
  wire  _GEN_2; // @[Xbar.scala 141:38]
  wire  _T_100; // @[Decoupled.scala 40:37]
  wire  in_0_w_valid; // @[Xbar.scala 145:43]
  wire  _T_122; // @[Mux.scala 27:72]
  wire  _T_123; // @[Mux.scala 27:72]
  wire  in_0_w_ready; // @[Mux.scala 27:72]
  wire  _T_103; // @[Xbar.scala 147:50]
  wire  out_0_ar_valid; // @[Xbar.scala 222:40]
  wire  out_1_ar_valid; // @[Xbar.scala 222:40]
  wire  out_0_aw_valid; // @[Xbar.scala 222:40]
  wire  out_1_aw_valid; // @[Xbar.scala 222:40]
  wire  _T_140; // @[Xbar.scala 256:60]
  wire  _T_146; // @[Xbar.scala 258:23]
  wire  _T_148; // @[Xbar.scala 258:12]
  wire  _T_149; // @[Xbar.scala 258:12]
  wire  _T_161; // @[Xbar.scala 256:60]
  wire  _T_167; // @[Xbar.scala 258:23]
  wire  _T_169; // @[Xbar.scala 258:12]
  wire  _T_170; // @[Xbar.scala 258:12]
  wire  _T_184; // @[Xbar.scala 256:60]
  wire  _T_190; // @[Xbar.scala 258:23]
  wire  _T_192; // @[Xbar.scala 258:12]
  wire  _T_193; // @[Xbar.scala 258:12]
  wire  _T_205; // @[Xbar.scala 256:60]
  wire  _T_211; // @[Xbar.scala 258:23]
  wire  _T_213; // @[Xbar.scala 258:12]
  wire  _T_214; // @[Xbar.scala 258:12]
  wire  _T_245; // @[Arbiter.scala 24:27]
  wire  _T_246; // @[Arbiter.scala 24:18]
  wire [1:0] _T_247; // @[Arbiter.scala 25:29]
  wire [2:0] _T_248; // @[package.scala 199:48]
  wire [1:0] _T_250; // @[package.scala 199:43]
  wire  _T_271; // @[Xbar.scala 258:13]
  wire  _T_273; // @[Xbar.scala 258:23]
  wire  _T_275; // @[Xbar.scala 258:12]
  wire  _T_276; // @[Xbar.scala 258:12]
  wire  _GEN_13; // @[Xbar.scala 266:21]
  wire  _GEN_14; // @[Xbar.scala 267:24]
  wire  _T_281_1; // @[Xbar.scala 270:24]
  wire [1:0] _T_306; // @[Cat.scala 29:58]
  reg [1:0] _T_313; // @[Arbiter.scala 20:23]
  reg [31:0] _RAND_11;
  wire [1:0] _T_314; // @[Arbiter.scala 21:30]
  wire [1:0] _T_315; // @[Arbiter.scala 21:28]
  wire [3:0] _T_316; // @[Cat.scala 29:58]
  wire [3:0] _GEN_24; // @[package.scala 208:43]
  wire [3:0] _T_318; // @[package.scala 208:43]
  wire [3:0] _T_321; // @[Arbiter.scala 22:66]
  wire [3:0] _GEN_25; // @[Arbiter.scala 22:58]
  wire [3:0] _T_322; // @[Arbiter.scala 22:58]
  wire [1:0] _T_325; // @[Arbiter.scala 23:39]
  wire [1:0] _T_326; // @[Arbiter.scala 23:18]
  wire  _T_327; // @[Arbiter.scala 24:27]
  wire  _T_328; // @[Arbiter.scala 24:18]
  wire [1:0] _T_329; // @[Arbiter.scala 25:29]
  wire [2:0] _T_330; // @[package.scala 199:48]
  wire [1:0] _T_332; // @[package.scala 199:43]
  wire  _T_338; // @[Xbar.scala 250:63]
  wire  _T_339; // @[Xbar.scala 250:63]
  wire  _T_342; // @[Xbar.scala 255:50]
  wire  _T_344; // @[Xbar.scala 256:60]
  wire  _T_347; // @[Xbar.scala 256:60]
  wire  _T_348; // @[Xbar.scala 256:57]
  wire  _T_351; // @[Xbar.scala 256:11]
  wire  _T_352; // @[Xbar.scala 256:11]
  wire  _T_353; // @[Xbar.scala 258:13]
  wire  _T_355; // @[Xbar.scala 258:23]
  wire  _T_357; // @[Xbar.scala 258:12]
  wire  _T_358; // @[Xbar.scala 258:12]
  wire  _T_361_1; // @[Xbar.scala 262:23]
  wire  _GEN_16; // @[Xbar.scala 266:21]
  wire  _GEN_17; // @[Xbar.scala 267:24]
  wire  _T_363_0; // @[Xbar.scala 270:24]
  wire  _T_363_1; // @[Xbar.scala 270:24]
  wire [2:0] _T_373; // @[Mux.scala 27:72]
  wire [2:0] _T_374; // @[Mux.scala 27:72]
  QueueCompatibility awIn_0 ( // @[Xbar.scala 55:47]
    .clock(awIn_0_clock),
    .reset(awIn_0_reset),
    .io_enq_ready(awIn_0_io_enq_ready),
    .io_enq_valid(awIn_0_io_enq_valid),
    .io_enq_bits(awIn_0_io_enq_bits),
    .io_deq_ready(awIn_0_io_deq_ready),
    .io_deq_valid(awIn_0_io_deq_valid),
    .io_deq_bits(awIn_0_io_deq_bits)
  );
  assign _T_1 = {1'b0,$signed(auto_in_ar_bits_addr)}; // @[Parameters.scala 137:49]
  assign _T_3 = $signed(_T_1) & 31'sh2000; // @[Parameters.scala 137:52]
  assign requestARIO_0_0 = $signed(_T_3) == 31'sh0; // @[Parameters.scala 137:67]
  assign _T_5 = auto_in_ar_bits_addr ^ 30'h2000; // @[Parameters.scala 137:31]
  assign _T_6 = {1'b0,$signed(_T_5)}; // @[Parameters.scala 137:49]
  assign _T_8 = $signed(_T_6) & 31'sh2000; // @[Parameters.scala 137:52]
  assign requestARIO_0_1 = $signed(_T_8) == 31'sh0; // @[Parameters.scala 137:67]
  assign _T_11 = {1'b0,$signed(auto_in_aw_bits_addr)}; // @[Parameters.scala 137:49]
  assign _T_13 = $signed(_T_11) & 31'sh2000; // @[Parameters.scala 137:52]
  assign requestAWIO_0_0 = $signed(_T_13) == 31'sh0; // @[Parameters.scala 137:67]
  assign _T_15 = auto_in_aw_bits_addr ^ 30'h2000; // @[Parameters.scala 137:31]
  assign _T_16 = {1'b0,$signed(_T_15)}; // @[Parameters.scala 137:49]
  assign _T_18 = $signed(_T_16) & 31'sh2000; // @[Parameters.scala 137:52]
  assign requestAWIO_0_1 = $signed(_T_18) == 31'sh0; // @[Parameters.scala 137:67]
  assign requestROI_1_0 = ~auto_out_1_r_bits_id; // @[Parameters.scala 47:9]
  assign requestBOI_1_0 = ~auto_out_1_b_bits_id; // @[Parameters.scala 47:9]
  assign _T_20 = {requestAWIO_0_1,requestAWIO_0_0}; // @[Xbar.scala 64:75]
  assign requestWIO_0_0 = awIn_0_io_deq_bits[0]; // @[Xbar.scala 65:73]
  assign requestWIO_0_1 = awIn_0_io_deq_bits[1]; // @[Xbar.scala 65:73]
  assign _T_27 = {requestARIO_0_1,requestARIO_0_0}; // @[Xbar.scala 93:45]
  assign in_0_ar_ready = requestARIO_0_1 & auto_out_1_ar_ready; // @[Mux.scala 27:72]
  assign _T_55 = _T_36 == 3'h0; // @[Xbar.scala 112:22]
  assign _T_54 = _T_37 == _T_27[1]; // @[Xbar.scala 111:75]
  assign _T_56 = _T_55 | _T_54; // @[Xbar.scala 112:34]
  assign _T_57 = _T_36 != 3'h7; // @[Xbar.scala 112:80]
  assign _T_59 = _T_56 & _T_57; // @[Xbar.scala 112:48]
  assign io_in_0_ar_ready = in_0_ar_ready & _T_59; // @[Xbar.scala 130:45]
  assign _T_31 = io_in_0_ar_ready & auto_in_ar_valid; // @[Decoupled.scala 40:37]
  assign _T_129 = auto_out_1_r_valid & requestROI_1_0; // @[Xbar.scala 222:40]
  assign _T_285 = _T_278_1 & _T_129; // @[Mux.scala 27:72]
  assign in_0_r_valid = _T_222 ? _T_129 : _T_285; // @[Xbar.scala 278:22]
  assign _T_33 = auto_in_r_ready & in_0_r_valid; // @[Decoupled.scala 40:37]
  assign _T_224 = {_T_129,1'h0}; // @[Cat.scala 29:58]
  assign _T_232 = ~_T_231; // @[Arbiter.scala 21:30]
  assign _T_233 = _T_224 & _T_232; // @[Arbiter.scala 21:28]
  assign _T_234 = {_T_233,_T_129,1'h0}; // @[Cat.scala 29:58]
  assign _GEN_18 = {{1'd0}, _T_234[3:1]}; // @[package.scala 208:43]
  assign _T_236 = _T_234 | _GEN_18; // @[package.scala 208:43]
  assign _T_239 = {_T_231, 2'h0}; // @[Arbiter.scala 22:66]
  assign _GEN_19 = {{1'd0}, _T_236[3:1]}; // @[Arbiter.scala 22:58]
  assign _T_240 = _GEN_19 | _T_239; // @[Arbiter.scala 22:58]
  assign _T_243 = _T_240[3:2] & _T_240[1:0]; // @[Arbiter.scala 23:39]
  assign _T_244 = ~_T_243; // @[Arbiter.scala 23:18]
  assign _T_257 = _T_244[1] & _T_129; // @[Xbar.scala 250:63]
  assign _T_279_1 = _T_222 ? _T_257 : _T_278_1; // @[Xbar.scala 262:23]
  assign _T_295 = {auto_out_1_r_bits_id,auto_out_1_r_bits_data,3'h1}; // @[Mux.scala 27:72]
  assign _T_296 = _T_279_1 ? _T_295 : 36'h0; // @[Mux.scala 27:72]
  assign in_0_r_bits_last = _T_296[0]; // @[Mux.scala 27:72]
  assign _T_35 = _T_33 & in_0_r_bits_last; // @[Xbar.scala 120:45]
  assign _GEN_20 = {{2'd0}, _T_31}; // @[Xbar.scala 106:30]
  assign _T_39 = _T_36 + _GEN_20; // @[Xbar.scala 106:30]
  assign _GEN_21 = {{2'd0}, _T_35}; // @[Xbar.scala 106:48]
  assign _T_41 = _T_39 - _GEN_21; // @[Xbar.scala 106:48]
  assign _T_42 = ~_T_35; // @[Xbar.scala 107:23]
  assign _T_43 = _T_36 != 3'h0; // @[Xbar.scala 107:43]
  assign _T_44 = _T_42 | _T_43; // @[Xbar.scala 107:34]
  assign _T_46 = _T_44 | reset; // @[Xbar.scala 107:22]
  assign _T_47 = ~_T_46; // @[Xbar.scala 107:22]
  assign _T_48 = ~_T_31; // @[Xbar.scala 108:23]
  assign _T_50 = _T_48 | _T_57; // @[Xbar.scala 108:34]
  assign _T_52 = _T_50 | reset; // @[Xbar.scala 108:22]
  assign _T_53 = ~_T_52; // @[Xbar.scala 108:22]
  assign _T_115 = requestAWIO_0_0 & auto_out_0_aw_ready; // @[Mux.scala 27:72]
  assign _T_116 = requestAWIO_0_1 & auto_out_1_aw_ready; // @[Mux.scala 27:72]
  assign in_0_aw_ready = _T_115 | _T_116; // @[Mux.scala 27:72]
  assign _T_94 = _T_90 | awIn_0_io_enq_ready; // @[Xbar.scala 139:57]
  assign _T_95 = in_0_aw_ready & _T_94; // @[Xbar.scala 139:45]
  assign _T_83 = _T_64 == 3'h0; // @[Xbar.scala 112:22]
  assign _T_82 = _T_65 == _T_20[1]; // @[Xbar.scala 111:75]
  assign _T_84 = _T_83 | _T_82; // @[Xbar.scala 112:34]
  assign _T_85 = _T_64 != 3'h7; // @[Xbar.scala 112:80]
  assign _T_87 = _T_84 & _T_85; // @[Xbar.scala 112:48]
  assign io_in_0_aw_ready = _T_95 & _T_87; // @[Xbar.scala 139:82]
  assign _T_60 = io_in_0_aw_ready & auto_in_aw_valid; // @[Decoupled.scala 40:37]
  assign _T_133 = auto_out_1_b_valid & requestBOI_1_0; // @[Xbar.scala 222:40]
  assign _T_305 = auto_out_0_b_valid | _T_133; // @[Xbar.scala 246:36]
  assign _T_366 = _T_360_0 & auto_out_0_b_valid; // @[Mux.scala 27:72]
  assign _T_367 = _T_360_1 & _T_133; // @[Mux.scala 27:72]
  assign _T_368 = _T_366 | _T_367; // @[Mux.scala 27:72]
  assign in_0_b_valid = _T_304 ? _T_305 : _T_368; // @[Xbar.scala 278:22]
  assign _T_62 = auto_in_b_ready & in_0_b_valid; // @[Decoupled.scala 40:37]
  assign _GEN_22 = {{2'd0}, _T_60}; // @[Xbar.scala 106:30]
  assign _T_67 = _T_64 + _GEN_22; // @[Xbar.scala 106:30]
  assign _GEN_23 = {{2'd0}, _T_62}; // @[Xbar.scala 106:48]
  assign _T_69 = _T_67 - _GEN_23; // @[Xbar.scala 106:48]
  assign _T_70 = ~_T_62; // @[Xbar.scala 107:23]
  assign _T_71 = _T_64 != 3'h0; // @[Xbar.scala 107:43]
  assign _T_72 = _T_70 | _T_71; // @[Xbar.scala 107:34]
  assign _T_74 = _T_72 | reset; // @[Xbar.scala 107:22]
  assign _T_75 = ~_T_74; // @[Xbar.scala 107:22]
  assign _T_76 = ~_T_60; // @[Xbar.scala 108:23]
  assign _T_78 = _T_76 | _T_85; // @[Xbar.scala 108:34]
  assign _T_80 = _T_78 | reset; // @[Xbar.scala 108:22]
  assign _T_81 = ~_T_80; // @[Xbar.scala 108:22]
  assign in_0_ar_valid = auto_in_ar_valid & _T_59; // @[Xbar.scala 129:45]
  assign _T_92 = auto_in_aw_valid & _T_94; // @[Xbar.scala 138:45]
  assign in_0_aw_valid = _T_92 & _T_87; // @[Xbar.scala 138:82]
  assign _T_97 = ~_T_90; // @[Xbar.scala 140:54]
  assign _T_99 = awIn_0_io_enq_ready & awIn_0_io_enq_valid; // @[Decoupled.scala 40:37]
  assign _GEN_2 = _T_99 | _T_90; // @[Xbar.scala 141:38]
  assign _T_100 = in_0_aw_ready & in_0_aw_valid; // @[Decoupled.scala 40:37]
  assign in_0_w_valid = auto_in_w_valid & awIn_0_io_deq_valid; // @[Xbar.scala 145:43]
  assign _T_122 = requestWIO_0_0 & auto_out_0_w_ready; // @[Mux.scala 27:72]
  assign _T_123 = requestWIO_0_1 & auto_out_1_w_ready; // @[Mux.scala 27:72]
  assign in_0_w_ready = _T_122 | _T_123; // @[Mux.scala 27:72]
  assign _T_103 = auto_in_w_valid & auto_in_w_bits_last; // @[Xbar.scala 147:50]
  assign out_0_ar_valid = in_0_ar_valid & requestARIO_0_0; // @[Xbar.scala 222:40]
  assign out_1_ar_valid = in_0_ar_valid & requestARIO_0_1; // @[Xbar.scala 222:40]
  assign out_0_aw_valid = in_0_aw_valid & requestAWIO_0_0; // @[Xbar.scala 222:40]
  assign out_1_aw_valid = in_0_aw_valid & requestAWIO_0_1; // @[Xbar.scala 222:40]
  assign _T_140 = ~out_0_aw_valid; // @[Xbar.scala 256:60]
  assign _T_146 = _T_140 | out_0_aw_valid; // @[Xbar.scala 258:23]
  assign _T_148 = _T_146 | reset; // @[Xbar.scala 258:12]
  assign _T_149 = ~_T_148; // @[Xbar.scala 258:12]
  assign _T_161 = ~out_0_ar_valid; // @[Xbar.scala 256:60]
  assign _T_167 = _T_161 | out_0_ar_valid; // @[Xbar.scala 258:23]
  assign _T_169 = _T_167 | reset; // @[Xbar.scala 258:12]
  assign _T_170 = ~_T_169; // @[Xbar.scala 258:12]
  assign _T_184 = ~out_1_aw_valid; // @[Xbar.scala 256:60]
  assign _T_190 = _T_184 | out_1_aw_valid; // @[Xbar.scala 258:23]
  assign _T_192 = _T_190 | reset; // @[Xbar.scala 258:12]
  assign _T_193 = ~_T_192; // @[Xbar.scala 258:12]
  assign _T_205 = ~out_1_ar_valid; // @[Xbar.scala 256:60]
  assign _T_211 = _T_205 | out_1_ar_valid; // @[Xbar.scala 258:23]
  assign _T_213 = _T_211 | reset; // @[Xbar.scala 258:12]
  assign _T_214 = ~_T_213; // @[Xbar.scala 258:12]
  assign _T_245 = _T_224 != 2'h0; // @[Arbiter.scala 24:27]
  assign _T_246 = _T_222 & _T_245; // @[Arbiter.scala 24:18]
  assign _T_247 = _T_244 & _T_224; // @[Arbiter.scala 25:29]
  assign _T_248 = {_T_247, 1'h0}; // @[package.scala 199:48]
  assign _T_250 = _T_247 | _T_248[1:0]; // @[package.scala 199:43]
  assign _T_271 = ~_T_129; // @[Xbar.scala 258:13]
  assign _T_273 = _T_271 | _T_257; // @[Xbar.scala 258:23]
  assign _T_275 = _T_273 | reset; // @[Xbar.scala 258:12]
  assign _T_276 = ~_T_275; // @[Xbar.scala 258:12]
  assign _GEN_13 = _T_129 ? 1'h0 : _T_222; // @[Xbar.scala 266:21]
  assign _GEN_14 = _T_33 | _GEN_13; // @[Xbar.scala 267:24]
  assign _T_281_1 = _T_222 ? _T_244[1] : _T_278_1; // @[Xbar.scala 270:24]
  assign _T_306 = {_T_133,auto_out_0_b_valid}; // @[Cat.scala 29:58]
  assign _T_314 = ~_T_313; // @[Arbiter.scala 21:30]
  assign _T_315 = _T_306 & _T_314; // @[Arbiter.scala 21:28]
  assign _T_316 = {_T_315,_T_133,auto_out_0_b_valid}; // @[Cat.scala 29:58]
  assign _GEN_24 = {{1'd0}, _T_316[3:1]}; // @[package.scala 208:43]
  assign _T_318 = _T_316 | _GEN_24; // @[package.scala 208:43]
  assign _T_321 = {_T_313, 2'h0}; // @[Arbiter.scala 22:66]
  assign _GEN_25 = {{1'd0}, _T_318[3:1]}; // @[Arbiter.scala 22:58]
  assign _T_322 = _GEN_25 | _T_321; // @[Arbiter.scala 22:58]
  assign _T_325 = _T_322[3:2] & _T_322[1:0]; // @[Arbiter.scala 23:39]
  assign _T_326 = ~_T_325; // @[Arbiter.scala 23:18]
  assign _T_327 = _T_306 != 2'h0; // @[Arbiter.scala 24:27]
  assign _T_328 = _T_304 & _T_327; // @[Arbiter.scala 24:18]
  assign _T_329 = _T_326 & _T_306; // @[Arbiter.scala 25:29]
  assign _T_330 = {_T_329, 1'h0}; // @[package.scala 199:48]
  assign _T_332 = _T_329 | _T_330[1:0]; // @[package.scala 199:43]
  assign _T_338 = _T_326[0] & auto_out_0_b_valid; // @[Xbar.scala 250:63]
  assign _T_339 = _T_326[1] & _T_133; // @[Xbar.scala 250:63]
  assign _T_342 = _T_338 | _T_339; // @[Xbar.scala 255:50]
  assign _T_344 = ~_T_338; // @[Xbar.scala 256:60]
  assign _T_347 = ~_T_339; // @[Xbar.scala 256:60]
  assign _T_348 = _T_344 | _T_347; // @[Xbar.scala 256:57]
  assign _T_351 = _T_348 | reset; // @[Xbar.scala 256:11]
  assign _T_352 = ~_T_351; // @[Xbar.scala 256:11]
  assign _T_353 = ~_T_305; // @[Xbar.scala 258:13]
  assign _T_355 = _T_353 | _T_342; // @[Xbar.scala 258:23]
  assign _T_357 = _T_355 | reset; // @[Xbar.scala 258:12]
  assign _T_358 = ~_T_357; // @[Xbar.scala 258:12]
  assign _T_361_1 = _T_304 ? _T_339 : _T_360_1; // @[Xbar.scala 262:23]
  assign _GEN_16 = _T_305 ? 1'h0 : _T_304; // @[Xbar.scala 266:21]
  assign _GEN_17 = _T_62 | _GEN_16; // @[Xbar.scala 267:24]
  assign _T_363_0 = _T_304 ? _T_326[0] : _T_360_0; // @[Xbar.scala 270:24]
  assign _T_363_1 = _T_304 ? _T_326[1] : _T_360_1; // @[Xbar.scala 270:24]
  assign _T_373 = {auto_out_1_b_bits_id,2'h0}; // @[Mux.scala 27:72]
  assign _T_374 = _T_361_1 ? _T_373 : 3'h0; // @[Mux.scala 27:72]
  assign auto_in_aw_ready = _T_95 & _T_87; // @[LazyModule.scala 173:31]
  assign auto_in_w_ready = in_0_w_ready & awIn_0_io_deq_valid; // @[LazyModule.scala 173:31]
  assign auto_in_b_valid = _T_304 ? _T_305 : _T_368; // @[LazyModule.scala 173:31]
  assign auto_in_b_bits_resp = _T_374[1:0]; // @[LazyModule.scala 173:31]
  assign auto_in_ar_ready = in_0_ar_ready & _T_59; // @[LazyModule.scala 173:31]
  assign auto_in_r_valid = _T_222 ? _T_129 : _T_285; // @[LazyModule.scala 173:31]
  assign auto_in_r_bits_data = _T_296[34:3]; // @[LazyModule.scala 173:31]
  assign auto_in_r_bits_resp = _T_296[2:1]; // @[LazyModule.scala 173:31]
  assign auto_in_r_bits_last = _T_296[0]; // @[LazyModule.scala 173:31]
  assign auto_out_1_aw_valid = in_0_aw_valid & requestAWIO_0_1; // @[LazyModule.scala 173:49]
  assign auto_out_1_aw_bits_id = auto_in_aw_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_1_aw_bits_addr = auto_in_aw_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_1_w_valid = in_0_w_valid & requestWIO_0_1; // @[LazyModule.scala 173:49]
  assign auto_out_1_w_bits_data = auto_in_w_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_1_w_bits_strb = auto_in_w_bits_strb; // @[LazyModule.scala 173:49]
  assign auto_out_1_b_ready = auto_in_b_ready & _T_363_1; // @[LazyModule.scala 173:49]
  assign auto_out_1_ar_valid = in_0_ar_valid & requestARIO_0_1; // @[LazyModule.scala 173:49]
  assign auto_out_1_ar_bits_id = auto_in_ar_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_1_ar_bits_addr = auto_in_ar_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_1_ar_bits_size = auto_in_ar_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_1_r_ready = auto_in_r_ready & _T_281_1; // @[LazyModule.scala 173:49]
  assign auto_out_0_aw_valid = in_0_aw_valid & requestAWIO_0_0; // @[LazyModule.scala 173:49]
  assign auto_out_0_aw_bits_addr = auto_in_aw_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_0_w_valid = in_0_w_valid & requestWIO_0_0; // @[LazyModule.scala 173:49]
  assign auto_out_0_w_bits_data = auto_in_w_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_0_b_ready = auto_in_b_ready & _T_363_0; // @[LazyModule.scala 173:49]
  assign awIn_0_clock = clock;
  assign awIn_0_reset = reset;
  assign awIn_0_io_enq_valid = auto_in_aw_valid & _T_97; // @[Xbar.scala 140:30]
  assign awIn_0_io_enq_bits = {requestAWIO_0_1,requestAWIO_0_0}; // @[Xbar.scala 64:57]
  assign awIn_0_io_deq_ready = _T_103 & in_0_w_ready; // @[Xbar.scala 147:30]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_36 = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_37 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_222 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_278_1 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_231 = _RAND_4[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_90 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_64 = _RAND_6[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_65 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_304 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_360_0 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_360_1 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_313 = _RAND_11[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      _T_36 <= 3'h0;
    end else begin
      _T_36 <= _T_41;
    end
    if (_T_31) begin
      _T_37 <= _T_27[1];
    end
    _T_222 <= reset | _GEN_14;
    if (reset) begin
      _T_278_1 <= 1'h0;
    end else if (_T_222) begin
      _T_278_1 <= _T_257;
    end
    if (reset) begin
      _T_231 <= 2'h3;
    end else if (_T_246) begin
      _T_231 <= _T_250;
    end
    if (reset) begin
      _T_90 <= 1'h0;
    end else if (_T_100) begin
      _T_90 <= 1'h0;
    end else begin
      _T_90 <= _GEN_2;
    end
    if (reset) begin
      _T_64 <= 3'h0;
    end else begin
      _T_64 <= _T_69;
    end
    if (_T_60) begin
      _T_65 <= _T_20[1];
    end
    _T_304 <= reset | _GEN_17;
    if (reset) begin
      _T_360_0 <= 1'h0;
    end else if (_T_304) begin
      _T_360_0 <= _T_338;
    end
    if (reset) begin
      _T_360_1 <= 1'h0;
    end else if (_T_304) begin
      _T_360_1 <= _T_339;
    end
    if (reset) begin
      _T_313 <= 2'h3;
    end else if (_T_328) begin
      _T_313 <= _T_332;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_47) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:107 assert (!resp_fire || count =/= UInt(0))\n"); // @[Xbar.scala 107:22]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_47) begin
          $fatal; // @[Xbar.scala 107:22]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_53) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:108 assert (!req_fire  || count =/= UInt(flight))\n"); // @[Xbar.scala 108:22]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_53) begin
          $fatal; // @[Xbar.scala 108:22]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_75) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:107 assert (!resp_fire || count =/= UInt(0))\n"); // @[Xbar.scala 107:22]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_75) begin
          $fatal; // @[Xbar.scala 107:22]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_81) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:108 assert (!req_fire  || count =/= UInt(flight))\n"); // @[Xbar.scala 108:22]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_81) begin
          $fatal; // @[Xbar.scala 108:22]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_149) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_149) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_170) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_170) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_193) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_193) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_214) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_214) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_276) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_276) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_352) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:256 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n"); // @[Xbar.scala 256:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_352) begin
          $fatal; // @[Xbar.scala 256:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_358) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_358) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module PLFGDspBlockMem(
  input         clock,
  input         reset,
  output        auto_mem_in_aw_ready,
  input         auto_mem_in_aw_valid,
  input         auto_mem_in_aw_bits_id,
  input  [29:0] auto_mem_in_aw_bits_addr,
  output        auto_mem_in_w_ready,
  input         auto_mem_in_w_valid,
  input  [31:0] auto_mem_in_w_bits_data,
  input  [3:0]  auto_mem_in_w_bits_strb,
  input         auto_mem_in_w_bits_last,
  input         auto_mem_in_b_ready,
  output        auto_mem_in_b_valid,
  output [1:0]  auto_mem_in_b_bits_resp,
  output        auto_mem_in_ar_ready,
  input         auto_mem_in_ar_valid,
  input         auto_mem_in_ar_bits_id,
  input  [29:0] auto_mem_in_ar_bits_addr,
  input  [2:0]  auto_mem_in_ar_bits_size,
  input         auto_mem_in_r_ready,
  output        auto_mem_in_r_valid,
  output [31:0] auto_mem_in_r_bits_data,
  output [1:0]  auto_mem_in_r_bits_resp,
  output        auto_mem_in_r_bits_last,
  input         auto_stream_out_ready,
  output        auto_stream_out_valid,
  output [31:0] auto_stream_out_bits_data,
  output        auto_stream_out_bits_last
);
  wire  axi4xbar_clock; // @[Xbar.scala 211:30]
  wire  axi4xbar_reset; // @[Xbar.scala 211:30]
  wire  axi4xbar_auto_in_aw_ready; // @[Xbar.scala 211:30]
  wire  axi4xbar_auto_in_aw_valid; // @[Xbar.scala 211:30]
  wire  axi4xbar_auto_in_aw_bits_id; // @[Xbar.scala 211:30]
  wire [29:0] axi4xbar_auto_in_aw_bits_addr; // @[Xbar.scala 211:30]
  wire  axi4xbar_auto_in_w_ready; // @[Xbar.scala 211:30]
  wire  axi4xbar_auto_in_w_valid; // @[Xbar.scala 211:30]
  wire [31:0] axi4xbar_auto_in_w_bits_data; // @[Xbar.scala 211:30]
  wire [3:0] axi4xbar_auto_in_w_bits_strb; // @[Xbar.scala 211:30]
  wire  axi4xbar_auto_in_w_bits_last; // @[Xbar.scala 211:30]
  wire  axi4xbar_auto_in_b_ready; // @[Xbar.scala 211:30]
  wire  axi4xbar_auto_in_b_valid; // @[Xbar.scala 211:30]
  wire [1:0] axi4xbar_auto_in_b_bits_resp; // @[Xbar.scala 211:30]
  wire  axi4xbar_auto_in_ar_ready; // @[Xbar.scala 211:30]
  wire  axi4xbar_auto_in_ar_valid; // @[Xbar.scala 211:30]
  wire  axi4xbar_auto_in_ar_bits_id; // @[Xbar.scala 211:30]
  wire [29:0] axi4xbar_auto_in_ar_bits_addr; // @[Xbar.scala 211:30]
  wire [2:0] axi4xbar_auto_in_ar_bits_size; // @[Xbar.scala 211:30]
  wire  axi4xbar_auto_in_r_ready; // @[Xbar.scala 211:30]
  wire  axi4xbar_auto_in_r_valid; // @[Xbar.scala 211:30]
  wire [31:0] axi4xbar_auto_in_r_bits_data; // @[Xbar.scala 211:30]
  wire [1:0] axi4xbar_auto_in_r_bits_resp; // @[Xbar.scala 211:30]
  wire  axi4xbar_auto_in_r_bits_last; // @[Xbar.scala 211:30]
  wire  axi4xbar_auto_out_1_aw_ready; // @[Xbar.scala 211:30]
  wire  axi4xbar_auto_out_1_aw_valid; // @[Xbar.scala 211:30]
  wire  axi4xbar_auto_out_1_aw_bits_id; // @[Xbar.scala 211:30]
  wire [29:0] axi4xbar_auto_out_1_aw_bits_addr; // @[Xbar.scala 211:30]
  wire  axi4xbar_auto_out_1_w_ready; // @[Xbar.scala 211:30]
  wire  axi4xbar_auto_out_1_w_valid; // @[Xbar.scala 211:30]
  wire [31:0] axi4xbar_auto_out_1_w_bits_data; // @[Xbar.scala 211:30]
  wire [3:0] axi4xbar_auto_out_1_w_bits_strb; // @[Xbar.scala 211:30]
  wire  axi4xbar_auto_out_1_b_ready; // @[Xbar.scala 211:30]
  wire  axi4xbar_auto_out_1_b_valid; // @[Xbar.scala 211:30]
  wire  axi4xbar_auto_out_1_b_bits_id; // @[Xbar.scala 211:30]
  wire  axi4xbar_auto_out_1_ar_ready; // @[Xbar.scala 211:30]
  wire  axi4xbar_auto_out_1_ar_valid; // @[Xbar.scala 211:30]
  wire  axi4xbar_auto_out_1_ar_bits_id; // @[Xbar.scala 211:30]
  wire [29:0] axi4xbar_auto_out_1_ar_bits_addr; // @[Xbar.scala 211:30]
  wire [2:0] axi4xbar_auto_out_1_ar_bits_size; // @[Xbar.scala 211:30]
  wire  axi4xbar_auto_out_1_r_ready; // @[Xbar.scala 211:30]
  wire  axi4xbar_auto_out_1_r_valid; // @[Xbar.scala 211:30]
  wire  axi4xbar_auto_out_1_r_bits_id; // @[Xbar.scala 211:30]
  wire [31:0] axi4xbar_auto_out_1_r_bits_data; // @[Xbar.scala 211:30]
  wire  axi4xbar_auto_out_0_aw_ready; // @[Xbar.scala 211:30]
  wire  axi4xbar_auto_out_0_aw_valid; // @[Xbar.scala 211:30]
  wire [29:0] axi4xbar_auto_out_0_aw_bits_addr; // @[Xbar.scala 211:30]
  wire  axi4xbar_auto_out_0_w_ready; // @[Xbar.scala 211:30]
  wire  axi4xbar_auto_out_0_w_valid; // @[Xbar.scala 211:30]
  wire [31:0] axi4xbar_auto_out_0_w_bits_data; // @[Xbar.scala 211:30]
  wire  axi4xbar_auto_out_0_b_ready; // @[Xbar.scala 211:30]
  wire  axi4xbar_auto_out_0_b_valid; // @[Xbar.scala 211:30]
  reg [25:0] configParamsMem1 [0:15]; // @[PLFGDspBlockMem.scala 110:39]
  reg [31:0] _RAND_0;
  wire [25:0] configParamsMem1__T_64_data; // @[PLFGDspBlockMem.scala 110:39]
  wire [3:0] configParamsMem1__T_64_addr; // @[PLFGDspBlockMem.scala 110:39]
  wire [25:0] configParamsMem1__T_14_data; // @[PLFGDspBlockMem.scala 110:39]
  wire [3:0] configParamsMem1__T_14_addr; // @[PLFGDspBlockMem.scala 110:39]
  wire  configParamsMem1__T_14_mask; // @[PLFGDspBlockMem.scala 110:39]
  wire  configParamsMem1__T_14_en; // @[PLFGDspBlockMem.scala 110:39]
  reg  configParamsMem1__T_64_en_pipe_0;
  reg [31:0] _RAND_1;
  reg [3:0] configParamsMem1__T_64_addr_pipe_0;
  reg [31:0] _RAND_2;
  wire  Queue_clock; // @[Decoupled.scala 287:21]
  wire  Queue_reset; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_read; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_enq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_extra; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_read; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_deq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_extra; // @[Decoupled.scala 287:21]
  reg  w_full1; // @[PLFGDspBlockMem.scala 114:26]
  reg [31:0] _RAND_3;
  wire [29:0] ramIn1_aw_bits_addr; // @[Nodes.scala 370:76 LazyModule.scala 167:31]
  wire  _T_5; // @[PLFGDspBlockMem.scala 119:62]
  wire  ramIn1_b_ready; // @[Nodes.scala 370:76 LazyModule.scala 167:31]
  wire  _T_6; // @[PLFGDspBlockMem.scala 119:59]
  wire  ramIn1_w_valid; // @[Nodes.scala 370:76 LazyModule.scala 167:31]
  wire  ramIn1_aw_ready; // @[PLFGDspBlockMem.scala 119:40]
  wire  ramIn1_aw_valid; // @[Nodes.scala 370:76 LazyModule.scala 167:31]
  wire  _T_11; // @[Decoupled.scala 40:37]
  wire  _GEN_0; // @[PLFGDspBlockMem.scala 121:29]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_1; // @[PLFGDspBlockMem.scala 122:29]
  wire [31:0] ramIn1_w_bits_data; // @[Nodes.scala 370:76 LazyModule.scala 167:31]
  reg  enable; // @[PLFGDspBlockMem.scala 130:25]
  reg [31:0] _RAND_4;
  reg  reset_bit; // @[PLFGDspBlockMem.scala 131:28]
  reg [31:0] _RAND_5;
  reg [1:0] frameNum; // @[PLFGDspBlockMem.scala 132:27]
  reg [31:0] _RAND_6;
  reg [15:0] startingPoint; // @[PLFGDspBlockMem.scala 133:32]
  reg [31:0] _RAND_7;
  reg [7:0] interframeNumOfSamples; // @[PLFGDspBlockMem.scala 134:41]
  reg [31:0] _RAND_8;
  reg [2:0] differentChirpsNum; // @[PLFGDspBlockMem.scala 135:37]
  reg [31:0] _RAND_9;
  reg [15:0] currentVal; // @[PLFGDspBlockMem.scala 138:29]
  reg [31:0] _RAND_10;
  reg [7:0] samplesCounter; // @[PLFGDspBlockMem.scala 139:33]
  reg [31:0] _RAND_11;
  reg [1:0] segmentCounter; // @[PLFGDspBlockMem.scala 140:33]
  reg [31:0] _RAND_12;
  reg [1:0] frameCounter; // @[PLFGDspBlockMem.scala 141:31]
  reg [31:0] _RAND_13;
  reg [5:0] framePauseCounter; // @[PLFGDspBlockMem.scala 142:36]
  reg [31:0] _RAND_14;
  reg  end_; // @[PLFGDspBlockMem.scala 143:22]
  reg [31:0] _RAND_15;
  reg [7:0] samplesCounter2; // @[PLFGDspBlockMem.scala 145:34]
  reg [31:0] _RAND_16;
  reg [1:0] segmentCounter2; // @[PLFGDspBlockMem.scala 146:34]
  reg [31:0] _RAND_17;
  reg [1:0] frameCounter2; // @[PLFGDspBlockMem.scala 147:32]
  reg [31:0] _RAND_18;
  reg  end2; // @[PLFGDspBlockMem.scala 149:23]
  reg [31:0] _RAND_19;
  reg [2:0] repeatedChirpsCounter; // @[PLFGDspBlockMem.scala 151:40]
  reg [31:0] _RAND_20;
  reg [2:0] differentChirpsCounter; // @[PLFGDspBlockMem.scala 152:41]
  reg [31:0] _RAND_21;
  reg [2:0] _T_19; // @[PLFGDspBlockMem.scala 154:49]
  reg [31:0] _RAND_22;
  reg [2:0] repeatedChirpsCounter2; // @[PLFGDspBlockMem.scala 154:41]
  reg [31:0] _RAND_23;
  reg [2:0] _T_20; // @[PLFGDspBlockMem.scala 155:50]
  reg [31:0] _RAND_24;
  reg [2:0] differentChirpsCounter2; // @[PLFGDspBlockMem.scala 155:42]
  reg [31:0] _RAND_25;
  reg [1:0] segmentNums_0; // @[PLFGDspBlockMem.scala 158:30]
  reg [31:0] _RAND_26;
  reg [1:0] segmentNums_1; // @[PLFGDspBlockMem.scala 158:30]
  reg [31:0] _RAND_27;
  reg [1:0] segmentNums_2; // @[PLFGDspBlockMem.scala 158:30]
  reg [31:0] _RAND_28;
  reg [1:0] segmentNums_3; // @[PLFGDspBlockMem.scala 158:30]
  reg [31:0] _RAND_29;
  reg [2:0] repeatedChirpNums_0; // @[PLFGDspBlockMem.scala 159:36]
  reg [31:0] _RAND_30;
  reg [2:0] repeatedChirpNums_1; // @[PLFGDspBlockMem.scala 159:36]
  reg [31:0] _RAND_31;
  reg [2:0] repeatedChirpNums_2; // @[PLFGDspBlockMem.scala 159:36]
  reg [31:0] _RAND_32;
  reg [2:0] repeatedChirpNums_3; // @[PLFGDspBlockMem.scala 159:36]
  reg [31:0] _RAND_33;
  reg [2:0] repeatedChirpNums_4; // @[PLFGDspBlockMem.scala 159:36]
  reg [31:0] _RAND_34;
  reg [2:0] repeatedChirpNums_5; // @[PLFGDspBlockMem.scala 159:36]
  reg [31:0] _RAND_35;
  reg [2:0] repeatedChirpNums_6; // @[PLFGDspBlockMem.scala 159:36]
  reg [31:0] _RAND_36;
  reg [2:0] repeatedChirpNums_7; // @[PLFGDspBlockMem.scala 159:36]
  reg [31:0] _RAND_37;
  reg [1:0] chirpOrdinalNums_0; // @[PLFGDspBlockMem.scala 160:35]
  reg [31:0] _RAND_38;
  reg [1:0] chirpOrdinalNums_1; // @[PLFGDspBlockMem.scala 160:35]
  reg [31:0] _RAND_39;
  reg [1:0] chirpOrdinalNums_2; // @[PLFGDspBlockMem.scala 160:35]
  reg [31:0] _RAND_40;
  reg [1:0] chirpOrdinalNums_3; // @[PLFGDspBlockMem.scala 160:35]
  reg [31:0] _RAND_41;
  reg [1:0] chirpOrdinalNums_4; // @[PLFGDspBlockMem.scala 160:35]
  reg [31:0] _RAND_42;
  reg [1:0] chirpOrdinalNums_5; // @[PLFGDspBlockMem.scala 160:35]
  reg [31:0] _RAND_43;
  reg [1:0] chirpOrdinalNums_6; // @[PLFGDspBlockMem.scala 160:35]
  reg [31:0] _RAND_44;
  reg [1:0] chirpOrdinalNums_7; // @[PLFGDspBlockMem.scala 160:35]
  reg [31:0] _RAND_45;
  wire [25:0] dataFromMem; // @[PLFGDspBlockMem.scala 162:27 PLFGDspBlockMem.scala 163:17]
  wire  _T_66; // @[UIntTypeClass.scala 54:47]
  wire [7:0] _T_70; // @[UIntTypeClass.scala 18:40]
  wire [7:0] numsOfSamples; // @[PLFGDspBlockMem.scala 172:28]
  wire  slopeSigns; // @[PLFGDspBlockMem.scala 174:33]
  wire  segmentResets; // @[PLFGDspBlockMem.scala 175:36]
  wire  _T_2_aw_valid; // @[Nodes.scala 370:76 LazyModule.scala 167:31]
  wire  _T_2_w_valid; // @[Nodes.scala 370:76 LazyModule.scala 167:31]
  wire  _T_72; // @[RegisterRouter.scala 40:39]
  wire  _T_2_ar_valid; // @[Nodes.scala 370:76 LazyModule.scala 167:31]
  wire  _T_73; // @[RegisterRouter.scala 40:26]
  wire  _T_74; // @[RegisterRouter.scala 42:29]
  wire  _T_117_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 290:17]
  wire [29:0] _T_2_ar_bits_addr; // @[Nodes.scala 370:76 LazyModule.scala 167:31]
  wire [29:0] _T_2_aw_bits_addr; // @[Nodes.scala 370:76 LazyModule.scala 167:31]
  wire [29:0] _T_81; // @[RegisterRouter.scala 48:19]
  wire [4:0] _T_825; // @[Cat.scala 29:58]
  wire [5:0] _T_121; // @[RegisterRouter.scala 59:16]
  wire  _T_131; // @[RegisterRouter.scala 59:16]
  wire  _T_75; // @[RegisterRouter.scala 42:26]
  wire  _T_2_ar_bits_id; // @[Nodes.scala 370:76 LazyModule.scala 167:31]
  wire  _T_2_aw_bits_id; // @[Nodes.scala 370:76 LazyModule.scala 167:31]
  wire [2:0] _T_2_ar_bits_size; // @[Nodes.scala 370:76 LazyModule.scala 167:31]
  wire [1:0] _T_84; // @[OneHot.scala 65:12]
  wire [1:0] _T_86; // @[Misc.scala 200:81]
  wire  _T_87; // @[Misc.scala 204:21]
  wire  _T_90; // @[Misc.scala 209:20]
  wire  _T_92; // @[Misc.scala 213:38]
  wire  _T_93; // @[Misc.scala 213:29]
  wire  _T_95; // @[Misc.scala 213:38]
  wire  _T_96; // @[Misc.scala 213:29]
  wire  _T_99; // @[Misc.scala 209:20]
  wire  _T_100; // @[Misc.scala 212:27]
  wire  _T_101; // @[Misc.scala 213:38]
  wire  _T_102; // @[Misc.scala 213:29]
  wire  _T_103; // @[Misc.scala 212:27]
  wire  _T_104; // @[Misc.scala 213:38]
  wire  _T_105; // @[Misc.scala 213:29]
  wire  _T_106; // @[Misc.scala 212:27]
  wire  _T_107; // @[Misc.scala 213:38]
  wire  _T_108; // @[Misc.scala 213:29]
  wire  _T_109; // @[Misc.scala 212:27]
  wire  _T_110; // @[Misc.scala 213:38]
  wire  _T_111; // @[Misc.scala 213:29]
  wire [3:0] _T_114; // @[Cat.scala 29:58]
  wire [3:0] _T_2_w_bits_strb; // @[Nodes.scala 370:76 LazyModule.scala 167:31]
  wire [3:0] _T_116; // @[RegisterRouter.scala 54:25]
  wire [7:0] _T_183; // @[Bitwise.scala 72:12]
  wire [7:0] _T_185; // @[Bitwise.scala 72:12]
  wire [7:0] _T_187; // @[Bitwise.scala 72:12]
  wire [7:0] _T_189; // @[Bitwise.scala 72:12]
  wire [31:0] _T_192; // @[Cat.scala 29:58]
  wire  _T_892; // @[RegisterRouter.scala 59:16]
  wire [31:0] _T_826; // @[OneHot.scala 58:35]
  wire  _T_1059; // @[RegisterRouter.scala 59:16]
  wire  _T_1061; // @[RegisterRouter.scala 59:16]
  wire  _T_1062; // @[RegisterRouter.scala 59:16]
  wire  _T_218; // @[RegisterRouter.scala 59:16]
  wire [31:0] _T_2_w_bits_data; // @[Nodes.scala 370:76 LazyModule.scala 167:31]
  wire  _T_234; // @[RegisterRouter.scala 59:16]
  wire  _T_1086; // @[RegisterRouter.scala 59:16]
  wire  _T_1087; // @[RegisterRouter.scala 59:16]
  wire  _T_241; // @[RegisterRouter.scala 59:16]
  wire  _T_257; // @[RegisterRouter.scala 59:16]
  wire  _T_1111; // @[RegisterRouter.scala 59:16]
  wire  _T_1112; // @[RegisterRouter.scala 59:16]
  wire  _T_264; // @[RegisterRouter.scala 59:16]
  wire  _T_280; // @[RegisterRouter.scala 59:16]
  wire  _T_1181; // @[RegisterRouter.scala 59:16]
  wire  _T_1182; // @[RegisterRouter.scala 59:16]
  wire  _T_287; // @[RegisterRouter.scala 59:16]
  wire  _T_1186; // @[RegisterRouter.scala 59:16]
  wire  _T_1187; // @[RegisterRouter.scala 59:16]
  wire  _T_310; // @[RegisterRouter.scala 59:16]
  wire  _T_1131; // @[RegisterRouter.scala 59:16]
  wire  _T_1132; // @[RegisterRouter.scala 59:16]
  wire  _T_333; // @[RegisterRouter.scala 59:16]
  wire  _T_1161; // @[RegisterRouter.scala 59:16]
  wire  _T_1162; // @[RegisterRouter.scala 59:16]
  wire  _T_356; // @[RegisterRouter.scala 59:16]
  wire  _T_1066; // @[RegisterRouter.scala 59:16]
  wire  _T_1067; // @[RegisterRouter.scala 59:16]
  wire  _T_379; // @[RegisterRouter.scala 59:16]
  wire  _T_1091; // @[RegisterRouter.scala 59:16]
  wire  _T_1092; // @[RegisterRouter.scala 59:16]
  wire  _T_402; // @[RegisterRouter.scala 59:16]
  wire  _T_1166; // @[RegisterRouter.scala 59:16]
  wire  _T_1167; // @[RegisterRouter.scala 59:16]
  wire  _T_425; // @[RegisterRouter.scala 59:16]
  wire  _T_1106; // @[RegisterRouter.scala 59:16]
  wire  _T_1107; // @[RegisterRouter.scala 59:16]
  wire  _T_448; // @[RegisterRouter.scala 59:16]
  wire  _T_1126; // @[RegisterRouter.scala 59:16]
  wire  _T_1127; // @[RegisterRouter.scala 59:16]
  wire  _T_471; // @[RegisterRouter.scala 59:16]
  wire  _T_1071; // @[RegisterRouter.scala 59:16]
  wire  _T_1072; // @[RegisterRouter.scala 59:16]
  wire  _T_494; // @[RegisterRouter.scala 59:16]
  wire  _T_1146; // @[RegisterRouter.scala 59:16]
  wire  _T_1147; // @[RegisterRouter.scala 59:16]
  wire  _T_517; // @[RegisterRouter.scala 59:16]
  wire  _T_1171; // @[RegisterRouter.scala 59:16]
  wire  _T_1172; // @[RegisterRouter.scala 59:16]
  wire  _T_540; // @[RegisterRouter.scala 59:16]
  wire  _T_1121; // @[RegisterRouter.scala 59:16]
  wire  _T_1122; // @[RegisterRouter.scala 59:16]
  wire  _T_563; // @[RegisterRouter.scala 59:16]
  wire  _T_1096; // @[RegisterRouter.scala 59:16]
  wire  _T_1097; // @[RegisterRouter.scala 59:16]
  wire  _T_586; // @[RegisterRouter.scala 59:16]
  wire  _T_602; // @[RegisterRouter.scala 59:16]
  wire  _T_1076; // @[RegisterRouter.scala 59:16]
  wire  _T_1077; // @[RegisterRouter.scala 59:16]
  wire  _T_609; // @[RegisterRouter.scala 59:16]
  wire [9:0] _GEN_24; // @[RegField.scala 134:88]
  wire [9:0] _T_620; // @[RegisterRouter.scala 59:16]
  wire  _T_1151; // @[RegisterRouter.scala 59:16]
  wire  _T_1152; // @[RegisterRouter.scala 59:16]
  wire  _T_632; // @[RegisterRouter.scala 59:16]
  wire  _T_1141; // @[RegisterRouter.scala 59:16]
  wire  _T_1142; // @[RegisterRouter.scala 59:16]
  wire  _T_655; // @[RegisterRouter.scala 59:16]
  wire  _T_1116; // @[RegisterRouter.scala 59:16]
  wire  _T_1117; // @[RegisterRouter.scala 59:16]
  wire  _T_678; // @[RegisterRouter.scala 59:16]
  wire  _T_1176; // @[RegisterRouter.scala 59:16]
  wire  _T_1177; // @[RegisterRouter.scala 59:16]
  wire  _T_701; // @[RegisterRouter.scala 59:16]
  wire  _T_1101; // @[RegisterRouter.scala 59:16]
  wire  _T_1102; // @[RegisterRouter.scala 59:16]
  wire  _T_724; // @[RegisterRouter.scala 59:16]
  wire  _T_1156; // @[RegisterRouter.scala 59:16]
  wire  _T_1157; // @[RegisterRouter.scala 59:16]
  wire  _T_747; // @[RegisterRouter.scala 59:16]
  wire  _T_1081; // @[RegisterRouter.scala 59:16]
  wire  _T_1082; // @[RegisterRouter.scala 59:16]
  wire  _T_770; // @[RegisterRouter.scala 59:16]
  wire  _T_1136; // @[RegisterRouter.scala 59:16]
  wire  _T_1137; // @[RegisterRouter.scala 59:16]
  wire  _T_793; // @[RegisterRouter.scala 59:16]
  wire  _GEN_162; // @[MuxLiteral.scala 48:10]
  wire  _GEN_163; // @[MuxLiteral.scala 48:10]
  wire  _GEN_164; // @[MuxLiteral.scala 48:10]
  wire  _GEN_165; // @[MuxLiteral.scala 48:10]
  wire  _GEN_166; // @[MuxLiteral.scala 48:10]
  wire  _GEN_167; // @[MuxLiteral.scala 48:10]
  wire  _GEN_168; // @[MuxLiteral.scala 48:10]
  wire  _GEN_169; // @[MuxLiteral.scala 48:10]
  wire  _GEN_170; // @[MuxLiteral.scala 48:10]
  wire  _GEN_171; // @[MuxLiteral.scala 48:10]
  wire  _GEN_172; // @[MuxLiteral.scala 48:10]
  wire  _GEN_173; // @[MuxLiteral.scala 48:10]
  wire  _GEN_174; // @[MuxLiteral.scala 48:10]
  wire  _GEN_175; // @[MuxLiteral.scala 48:10]
  wire  _GEN_176; // @[MuxLiteral.scala 48:10]
  wire  _GEN_177; // @[MuxLiteral.scala 48:10]
  wire  _GEN_178; // @[MuxLiteral.scala 48:10]
  wire  _GEN_179; // @[MuxLiteral.scala 48:10]
  wire  _GEN_180; // @[MuxLiteral.scala 48:10]
  wire  _GEN_181; // @[MuxLiteral.scala 48:10]
  wire  _GEN_182; // @[MuxLiteral.scala 48:10]
  wire  _GEN_183; // @[MuxLiteral.scala 48:10]
  wire  _GEN_184; // @[MuxLiteral.scala 48:10]
  wire  _GEN_185; // @[MuxLiteral.scala 48:10]
  wire  _GEN_186; // @[MuxLiteral.scala 48:10]
  wire  _GEN_351; // @[MuxLiteral.scala 48:10]
  wire  _GEN_187; // @[MuxLiteral.scala 48:10]
  wire  _GEN_352; // @[MuxLiteral.scala 48:10]
  wire  _GEN_188; // @[MuxLiteral.scala 48:10]
  wire  _GEN_353; // @[MuxLiteral.scala 48:10]
  wire  _GEN_189; // @[MuxLiteral.scala 48:10]
  wire  _GEN_354; // @[MuxLiteral.scala 48:10]
  wire  _GEN_190; // @[MuxLiteral.scala 48:10]
  wire  _GEN_355; // @[MuxLiteral.scala 48:10]
  wire  _GEN_191; // @[MuxLiteral.scala 48:10]
  wire  _GEN_356; // @[MuxLiteral.scala 48:10]
  wire  _GEN_192; // @[MuxLiteral.scala 48:10]
  wire [15:0] _T_1564_0; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [15:0] _T_1564_1; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [15:0] _GEN_194; // @[MuxLiteral.scala 48:10]
  wire [15:0] _T_1564_2; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [15:0] _GEN_195; // @[MuxLiteral.scala 48:10]
  wire [15:0] _T_1564_3; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [15:0] _GEN_196; // @[MuxLiteral.scala 48:10]
  wire [15:0] _T_1564_4; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [15:0] _GEN_197; // @[MuxLiteral.scala 48:10]
  wire [15:0] _GEN_198; // @[MuxLiteral.scala 48:10]
  wire [15:0] _T_1564_6; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [15:0] _GEN_199; // @[MuxLiteral.scala 48:10]
  wire [15:0] _T_1564_7; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [15:0] _GEN_200; // @[MuxLiteral.scala 48:10]
  wire [15:0] _T_1564_8; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [15:0] _GEN_201; // @[MuxLiteral.scala 48:10]
  wire [15:0] _T_1564_9; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [15:0] _GEN_202; // @[MuxLiteral.scala 48:10]
  wire [15:0] _T_1564_10; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [15:0] _GEN_203; // @[MuxLiteral.scala 48:10]
  wire [15:0] _T_1564_11; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [15:0] _GEN_204; // @[MuxLiteral.scala 48:10]
  wire [15:0] _T_1564_12; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [15:0] _GEN_205; // @[MuxLiteral.scala 48:10]
  wire [15:0] _T_1564_13; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [15:0] _GEN_206; // @[MuxLiteral.scala 48:10]
  wire [15:0] _T_1564_14; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [15:0] _GEN_207; // @[MuxLiteral.scala 48:10]
  wire [15:0] _T_1564_15; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [15:0] _GEN_208; // @[MuxLiteral.scala 48:10]
  wire [15:0] _T_1564_16; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [15:0] _GEN_209; // @[MuxLiteral.scala 48:10]
  wire [15:0] _T_1564_17; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [15:0] _GEN_210; // @[MuxLiteral.scala 48:10]
  wire [15:0] _T_1564_18; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [15:0] _GEN_211; // @[MuxLiteral.scala 48:10]
  wire [15:0] _T_1564_19; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [15:0] _GEN_212; // @[MuxLiteral.scala 48:10]
  wire [15:0] _T_1564_20; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [15:0] _GEN_213; // @[MuxLiteral.scala 48:10]
  wire [15:0] _T_1564_21; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [15:0] _GEN_214; // @[MuxLiteral.scala 48:10]
  wire [15:0] _T_1564_22; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [15:0] _GEN_215; // @[MuxLiteral.scala 48:10]
  wire [15:0] _T_1564_23; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [15:0] _GEN_216; // @[MuxLiteral.scala 48:10]
  wire [15:0] _T_1564_24; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [15:0] _GEN_217; // @[MuxLiteral.scala 48:10]
  wire [15:0] _T_1564_25; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [15:0] _GEN_218; // @[MuxLiteral.scala 48:10]
  wire [15:0] _GEN_219; // @[MuxLiteral.scala 48:10]
  wire [15:0] _GEN_220; // @[MuxLiteral.scala 48:10]
  wire [15:0] _GEN_221; // @[MuxLiteral.scala 48:10]
  wire [15:0] _GEN_222; // @[MuxLiteral.scala 48:10]
  wire [15:0] _GEN_223; // @[MuxLiteral.scala 48:10]
  wire [15:0] _GEN_224; // @[MuxLiteral.scala 48:10]
  wire [15:0] _T_1566; // @[RegisterRouter.scala 59:16]
  wire  _T_1567_bits_read; // @[Decoupled.scala 308:19 Decoupled.scala 309:14]
  wire  _T_2_r_ready; // @[Nodes.scala 370:76 LazyModule.scala 167:31]
  wire  _T_2_b_ready; // @[Nodes.scala 370:76 LazyModule.scala 167:31]
  wire  _T_1567_valid; // @[Decoupled.scala 308:19 Decoupled.scala 310:15]
  wire  _T_1570; // @[RegisterRouter.scala 65:29]
  reg  enable2; // @[PLFGDspBlockMem.scala 218:26]
  reg [31:0] _RAND_46;
  reg [1:0] chirpIndexOld; // @[PLFGDspBlockMem.scala 219:32]
  reg [31:0] _RAND_47;
  reg  started; // @[PLFGDspBlockMem.scala 220:26]
  reg [31:0] _RAND_48;
  wire [1:0] _GEN_226; // @[PLFGDspBlockMem.scala 238:18]
  wire [1:0] _GEN_227; // @[PLFGDspBlockMem.scala 238:18]
  wire [1:0] _GEN_228; // @[PLFGDspBlockMem.scala 238:18]
  wire [1:0] _GEN_229; // @[PLFGDspBlockMem.scala 238:18]
  wire [1:0] _GEN_230; // @[PLFGDspBlockMem.scala 238:18]
  wire [1:0] _GEN_231; // @[PLFGDspBlockMem.scala 238:18]
  wire [1:0] _GEN_232; // @[PLFGDspBlockMem.scala 238:18]
  wire  _T_1573; // @[PLFGDspBlockMem.scala 239:19]
  wire  _T_1574; // @[PLFGDspBlockMem.scala 239:35]
  wire  _T_1575; // @[PLFGDspBlockMem.scala 239:32]
  wire [7:0] _T_1577; // @[PLFGDspBlockMem.scala 241:30]
  wire  _T_1578; // @[PLFGDspBlockMem.scala 241:37]
  wire [1:0] _T_1580; // @[PLFGDspBlockMem.scala 242:32]
  wire [1:0] chirpIndex; // @[PLFGDspBlockMem.scala 224:20]
  wire [1:0] _GEN_234; // @[PLFGDspBlockMem.scala 242:39]
  wire [1:0] _GEN_235; // @[PLFGDspBlockMem.scala 242:39]
  wire [1:0] _GEN_236; // @[PLFGDspBlockMem.scala 242:39]
  wire  _T_1581; // @[PLFGDspBlockMem.scala 242:39]
  wire [2:0] _T_1583; // @[PLFGDspBlockMem.scala 243:41]
  wire [2:0] _GEN_238; // @[PLFGDspBlockMem.scala 243:48]
  wire [2:0] _GEN_239; // @[PLFGDspBlockMem.scala 243:48]
  wire [2:0] _GEN_240; // @[PLFGDspBlockMem.scala 243:48]
  wire [2:0] _GEN_241; // @[PLFGDspBlockMem.scala 243:48]
  wire [2:0] _GEN_242; // @[PLFGDspBlockMem.scala 243:48]
  wire [2:0] _GEN_243; // @[PLFGDspBlockMem.scala 243:48]
  wire [2:0] _GEN_244; // @[PLFGDspBlockMem.scala 243:48]
  wire  _T_1584; // @[PLFGDspBlockMem.scala 243:48]
  wire [2:0] _T_1586; // @[PLFGDspBlockMem.scala 244:44]
  wire  _T_1587; // @[PLFGDspBlockMem.scala 244:51]
  wire  _T_1590; // @[PLFGDspBlockMem.scala 245:31]
  wire [5:0] _T_1592; // @[PLFGDspBlockMem.scala 247:43]
  wire [7:0] _GEN_357; // @[PLFGDspBlockMem.scala 247:50]
  wire  _T_1593; // @[PLFGDspBlockMem.scala 247:50]
  wire [1:0] _T_1597; // @[PLFGDspBlockMem.scala 258:38]
  wire  _T_1598; // @[PLFGDspBlockMem.scala 258:45]
  wire  _GEN_257; // @[PLFGDspBlockMem.scala 258:57]
  wire  _T_1616; // @[PLFGDspBlockMem.scala 298:20]
  wire  _T_1617; // @[PLFGDspBlockMem.scala 298:36]
  wire  _T_1618; // @[PLFGDspBlockMem.scala 298:33]
  wire [7:0] _T_1620; // @[PLFGDspBlockMem.scala 300:31]
  wire  _T_1621; // @[PLFGDspBlockMem.scala 300:38]
  wire [1:0] _T_1623; // @[PLFGDspBlockMem.scala 301:34]
  wire [1:0] _GEN_318; // @[PLFGDspBlockMem.scala 301:41]
  wire [1:0] _GEN_319; // @[PLFGDspBlockMem.scala 301:41]
  wire [1:0] _GEN_320; // @[PLFGDspBlockMem.scala 301:41]
  wire  _T_1626; // @[PLFGDspBlockMem.scala 301:41]
  wire [2:0] _T_1630; // @[PLFGDspBlockMem.scala 303:42]
  wire  _T_1631; // @[PLFGDspBlockMem.scala 303:49]
  wire [2:0] _T_1633; // @[PLFGDspBlockMem.scala 304:45]
  wire  _T_1634; // @[PLFGDspBlockMem.scala 304:52]
  wire  _T_1640; // @[PLFGDspBlockMem.scala 309:38]
  wire  _GEN_321; // @[PLFGDspBlockMem.scala 309:50]
  wire [15:0] _T_1652; // @[PLFGDspBlockMem.scala 326:73]
  wire [15:0] _T_1655; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] _T_1660; // @[FixedPointTypeClass.scala 30:68]
  wire  _T_1675; // @[PLFGDspBlockMem.scala 337:14]
  wire  _GEN_336; // @[PLFGDspBlockMem.scala 298:42]
  wire [15:0] _GEN_342; // @[PLFGDspBlockMem.scala 295:20]
  reg  _T_1679; // @[PLFGDspBlockMem.scala 345:39]
  reg [31:0] _RAND_49;
  wire  _T_1680; // @[PLFGDspBlockMem.scala 345:31]
  wire  _T_1681; // @[PLFGDspBlockMem.scala 345:28]
  reg  lastOutReg; // @[PLFGDspBlockMem.scala 351:29]
  reg [31:0] _RAND_50;
  reg  _T_1682; // @[PLFGDspBlockMem.scala 352:25]
  reg [31:0] _RAND_51;
  wire  _T_1683; // @[PLFGDspBlockMem.scala 352:17]
  wire  lastOut; // @[PLFGDspBlockMem.scala 352:14]
  reg  _T_1685; // @[PLFGDspBlockMem.scala 357:25]
  reg [31:0] _RAND_52;
  wire  _T_1686; // @[PLFGDspBlockMem.scala 357:17]
  wire  _T_1687; // @[PLFGDspBlockMem.scala 357:14]
  reg  _T_1688; // @[PLFGDspBlockMem.scala 359:36]
  reg [31:0] _RAND_53;
  wire  _T_1689; // @[PLFGDspBlockMem.scala 359:26]
  wire  _GEN_345; // @[PLFGDspBlockMem.scala 359:42]
  wire  _GEN_346; // @[PLFGDspBlockMem.scala 357:31]
  wire  _T_1691; // @[PLFGDspBlockMem.scala 362:46]
  wire  _T_1693; // @[PLFGDspBlockMem.scala 365:10]
  wire [2:0] _GEN_359; // @[UIntTypeClass.scala 39:41]
  wire [4:0] _T_1694; // @[UIntTypeClass.scala 39:41]
  wire [4:0] _GEN_360; // @[PLFGDspBlockMem.scala 367:57]
  wire [4:0] _T_1696; // @[PLFGDspBlockMem.scala 367:57]
  AXI4Xbar axi4xbar ( // @[Xbar.scala 211:30]
    .clock(axi4xbar_clock),
    .reset(axi4xbar_reset),
    .auto_in_aw_ready(axi4xbar_auto_in_aw_ready),
    .auto_in_aw_valid(axi4xbar_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4xbar_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4xbar_auto_in_aw_bits_addr),
    .auto_in_w_ready(axi4xbar_auto_in_w_ready),
    .auto_in_w_valid(axi4xbar_auto_in_w_valid),
    .auto_in_w_bits_data(axi4xbar_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi4xbar_auto_in_w_bits_strb),
    .auto_in_w_bits_last(axi4xbar_auto_in_w_bits_last),
    .auto_in_b_ready(axi4xbar_auto_in_b_ready),
    .auto_in_b_valid(axi4xbar_auto_in_b_valid),
    .auto_in_b_bits_resp(axi4xbar_auto_in_b_bits_resp),
    .auto_in_ar_ready(axi4xbar_auto_in_ar_ready),
    .auto_in_ar_valid(axi4xbar_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4xbar_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4xbar_auto_in_ar_bits_addr),
    .auto_in_ar_bits_size(axi4xbar_auto_in_ar_bits_size),
    .auto_in_r_ready(axi4xbar_auto_in_r_ready),
    .auto_in_r_valid(axi4xbar_auto_in_r_valid),
    .auto_in_r_bits_data(axi4xbar_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4xbar_auto_in_r_bits_resp),
    .auto_in_r_bits_last(axi4xbar_auto_in_r_bits_last),
    .auto_out_1_aw_ready(axi4xbar_auto_out_1_aw_ready),
    .auto_out_1_aw_valid(axi4xbar_auto_out_1_aw_valid),
    .auto_out_1_aw_bits_id(axi4xbar_auto_out_1_aw_bits_id),
    .auto_out_1_aw_bits_addr(axi4xbar_auto_out_1_aw_bits_addr),
    .auto_out_1_w_ready(axi4xbar_auto_out_1_w_ready),
    .auto_out_1_w_valid(axi4xbar_auto_out_1_w_valid),
    .auto_out_1_w_bits_data(axi4xbar_auto_out_1_w_bits_data),
    .auto_out_1_w_bits_strb(axi4xbar_auto_out_1_w_bits_strb),
    .auto_out_1_b_ready(axi4xbar_auto_out_1_b_ready),
    .auto_out_1_b_valid(axi4xbar_auto_out_1_b_valid),
    .auto_out_1_b_bits_id(axi4xbar_auto_out_1_b_bits_id),
    .auto_out_1_ar_ready(axi4xbar_auto_out_1_ar_ready),
    .auto_out_1_ar_valid(axi4xbar_auto_out_1_ar_valid),
    .auto_out_1_ar_bits_id(axi4xbar_auto_out_1_ar_bits_id),
    .auto_out_1_ar_bits_addr(axi4xbar_auto_out_1_ar_bits_addr),
    .auto_out_1_ar_bits_size(axi4xbar_auto_out_1_ar_bits_size),
    .auto_out_1_r_ready(axi4xbar_auto_out_1_r_ready),
    .auto_out_1_r_valid(axi4xbar_auto_out_1_r_valid),
    .auto_out_1_r_bits_id(axi4xbar_auto_out_1_r_bits_id),
    .auto_out_1_r_bits_data(axi4xbar_auto_out_1_r_bits_data),
    .auto_out_0_aw_ready(axi4xbar_auto_out_0_aw_ready),
    .auto_out_0_aw_valid(axi4xbar_auto_out_0_aw_valid),
    .auto_out_0_aw_bits_addr(axi4xbar_auto_out_0_aw_bits_addr),
    .auto_out_0_w_ready(axi4xbar_auto_out_0_w_ready),
    .auto_out_0_w_valid(axi4xbar_auto_out_0_w_valid),
    .auto_out_0_w_bits_data(axi4xbar_auto_out_0_w_bits_data),
    .auto_out_0_b_ready(axi4xbar_auto_out_0_b_ready),
    .auto_out_0_b_valid(axi4xbar_auto_out_0_b_valid)
  );
  Queue Queue ( // @[Decoupled.scala 287:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_read(Queue_io_enq_bits_read),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_extra(Queue_io_enq_bits_extra),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_read(Queue_io_deq_bits_read),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_extra(Queue_io_deq_bits_extra)
  );
  assign configParamsMem1__T_64_addr = configParamsMem1__T_64_addr_pipe_0;
  assign configParamsMem1__T_64_data = configParamsMem1[configParamsMem1__T_64_addr]; // @[PLFGDspBlockMem.scala 110:39]
  assign configParamsMem1__T_14_data = ramIn1_w_bits_data[25:0];
  assign configParamsMem1__T_14_addr = ramIn1_aw_bits_addr[5:2];
  assign configParamsMem1__T_14_mask = 1'h1;
  assign configParamsMem1__T_14_en = ramIn1_aw_ready & ramIn1_aw_valid;
  assign ramIn1_aw_bits_addr = axi4xbar_auto_out_0_aw_bits_addr; // @[Nodes.scala 370:76 LazyModule.scala 167:31]
  assign _T_5 = ~w_full1; // @[PLFGDspBlockMem.scala 119:62]
  assign ramIn1_b_ready = axi4xbar_auto_out_0_b_ready; // @[Nodes.scala 370:76 LazyModule.scala 167:31]
  assign _T_6 = ramIn1_b_ready | _T_5; // @[PLFGDspBlockMem.scala 119:59]
  assign ramIn1_w_valid = axi4xbar_auto_out_0_w_valid; // @[Nodes.scala 370:76 LazyModule.scala 167:31]
  assign ramIn1_aw_ready = ramIn1_w_valid & _T_6; // @[PLFGDspBlockMem.scala 119:40]
  assign ramIn1_aw_valid = axi4xbar_auto_out_0_aw_valid; // @[Nodes.scala 370:76 LazyModule.scala 167:31]
  assign _T_11 = ramIn1_b_ready & w_full1; // @[Decoupled.scala 40:37]
  assign _GEN_0 = _T_11 ? 1'h0 : w_full1; // @[PLFGDspBlockMem.scala 121:29]
  assign _T_12 = ramIn1_aw_ready & ramIn1_aw_valid; // @[Decoupled.scala 40:37]
  assign _GEN_1 = _T_12 | _GEN_0; // @[PLFGDspBlockMem.scala 122:29]
  assign ramIn1_w_bits_data = axi4xbar_auto_out_0_w_bits_data; // @[Nodes.scala 370:76 LazyModule.scala 167:31]
  assign dataFromMem = configParamsMem1__T_64_data; // @[PLFGDspBlockMem.scala 162:27 PLFGDspBlockMem.scala 163:17]
  assign _T_66 = dataFromMem[23:16] > 8'h1; // @[UIntTypeClass.scala 54:47]
  assign _T_70 = dataFromMem[23:16] + 8'h1; // @[UIntTypeClass.scala 18:40]
  assign numsOfSamples = _T_66 ? dataFromMem[23:16] : _T_70; // @[PLFGDspBlockMem.scala 172:28]
  assign slopeSigns = dataFromMem[24]; // @[PLFGDspBlockMem.scala 174:33]
  assign segmentResets = dataFromMem[25]; // @[PLFGDspBlockMem.scala 175:36]
  assign _T_2_aw_valid = axi4xbar_auto_out_1_aw_valid; // @[Nodes.scala 370:76 LazyModule.scala 167:31]
  assign _T_2_w_valid = axi4xbar_auto_out_1_w_valid; // @[Nodes.scala 370:76 LazyModule.scala 167:31]
  assign _T_72 = _T_2_aw_valid & _T_2_w_valid; // @[RegisterRouter.scala 40:39]
  assign _T_2_ar_valid = axi4xbar_auto_out_1_ar_valid; // @[Nodes.scala 370:76 LazyModule.scala 167:31]
  assign _T_73 = _T_2_ar_valid | _T_72; // @[RegisterRouter.scala 40:26]
  assign _T_74 = ~_T_2_ar_valid; // @[RegisterRouter.scala 42:29]
  assign _T_117_ready = Queue_io_enq_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 290:17]
  assign _T_2_ar_bits_addr = axi4xbar_auto_out_1_ar_bits_addr; // @[Nodes.scala 370:76 LazyModule.scala 167:31]
  assign _T_2_aw_bits_addr = axi4xbar_auto_out_1_aw_bits_addr; // @[Nodes.scala 370:76 LazyModule.scala 167:31]
  assign _T_81 = _T_2_ar_valid ? _T_2_ar_bits_addr : _T_2_aw_bits_addr; // @[RegisterRouter.scala 48:19]
  assign _T_825 = {_T_81[6],_T_81[5],_T_81[4],_T_81[3],_T_81[2]}; // @[Cat.scala 29:58]
  assign _T_121 = _T_81[7:2] & 6'h20; // @[RegisterRouter.scala 59:16]
  assign _T_131 = _T_121 == 6'h0; // @[RegisterRouter.scala 59:16]
  assign _T_75 = _T_117_ready & _T_74; // @[RegisterRouter.scala 42:26]
  assign _T_2_ar_bits_id = axi4xbar_auto_out_1_ar_bits_id; // @[Nodes.scala 370:76 LazyModule.scala 167:31]
  assign _T_2_aw_bits_id = axi4xbar_auto_out_1_aw_bits_id; // @[Nodes.scala 370:76 LazyModule.scala 167:31]
  assign _T_2_ar_bits_size = axi4xbar_auto_out_1_ar_bits_size; // @[Nodes.scala 370:76 LazyModule.scala 167:31]
  assign _T_84 = 2'h1 << _T_2_ar_bits_size[0]; // @[OneHot.scala 65:12]
  assign _T_86 = _T_84 | 2'h1; // @[Misc.scala 200:81]
  assign _T_87 = _T_2_ar_bits_size >= 3'h2; // @[Misc.scala 204:21]
  assign _T_90 = ~_T_2_ar_bits_addr[1]; // @[Misc.scala 209:20]
  assign _T_92 = _T_86[1] & _T_90; // @[Misc.scala 213:38]
  assign _T_93 = _T_87 | _T_92; // @[Misc.scala 213:29]
  assign _T_95 = _T_86[1] & _T_2_ar_bits_addr[1]; // @[Misc.scala 213:38]
  assign _T_96 = _T_87 | _T_95; // @[Misc.scala 213:29]
  assign _T_99 = ~_T_2_ar_bits_addr[0]; // @[Misc.scala 209:20]
  assign _T_100 = _T_90 & _T_99; // @[Misc.scala 212:27]
  assign _T_101 = _T_86[0] & _T_100; // @[Misc.scala 213:38]
  assign _T_102 = _T_93 | _T_101; // @[Misc.scala 213:29]
  assign _T_103 = _T_90 & _T_2_ar_bits_addr[0]; // @[Misc.scala 212:27]
  assign _T_104 = _T_86[0] & _T_103; // @[Misc.scala 213:38]
  assign _T_105 = _T_93 | _T_104; // @[Misc.scala 213:29]
  assign _T_106 = _T_2_ar_bits_addr[1] & _T_99; // @[Misc.scala 212:27]
  assign _T_107 = _T_86[0] & _T_106; // @[Misc.scala 213:38]
  assign _T_108 = _T_96 | _T_107; // @[Misc.scala 213:29]
  assign _T_109 = _T_2_ar_bits_addr[1] & _T_2_ar_bits_addr[0]; // @[Misc.scala 212:27]
  assign _T_110 = _T_86[0] & _T_109; // @[Misc.scala 213:38]
  assign _T_111 = _T_96 | _T_110; // @[Misc.scala 213:29]
  assign _T_114 = {_T_111,_T_108,_T_105,_T_102}; // @[Cat.scala 29:58]
  assign _T_2_w_bits_strb = axi4xbar_auto_out_1_w_bits_strb; // @[Nodes.scala 370:76 LazyModule.scala 167:31]
  assign _T_116 = _T_2_ar_valid ? _T_114 : _T_2_w_bits_strb; // @[RegisterRouter.scala 54:25]
  assign _T_183 = _T_116[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_185 = _T_116[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_187 = _T_116[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_189 = _T_116[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_192 = {_T_189,_T_187,_T_185,_T_183}; // @[Cat.scala 29:58]
  assign _T_892 = _T_73 & _T_117_ready; // @[RegisterRouter.scala 59:16]
  assign _T_826 = 32'h1 << _T_825; // @[OneHot.scala 58:35]
  assign _T_1059 = _T_892 & _T_74; // @[RegisterRouter.scala 59:16]
  assign _T_1061 = _T_1059 & _T_826[0]; // @[RegisterRouter.scala 59:16]
  assign _T_1062 = _T_1061 & _T_131; // @[RegisterRouter.scala 59:16]
  assign _T_218 = _T_1062 & _T_192[0]; // @[RegisterRouter.scala 59:16]
  assign _T_2_w_bits_data = axi4xbar_auto_out_1_w_bits_data; // @[Nodes.scala 370:76 LazyModule.scala 167:31]
  assign _T_234 = _T_192[15:0] == 16'hffff; // @[RegisterRouter.scala 59:16]
  assign _T_1086 = _T_1059 & _T_826[5]; // @[RegisterRouter.scala 59:16]
  assign _T_1087 = _T_1086 & _T_131; // @[RegisterRouter.scala 59:16]
  assign _T_241 = _T_1087 & _T_234; // @[RegisterRouter.scala 59:16]
  assign _T_257 = _T_192[2:0] == 3'h7; // @[RegisterRouter.scala 59:16]
  assign _T_1111 = _T_1059 & _T_826[10]; // @[RegisterRouter.scala 59:16]
  assign _T_1112 = _T_1111 & _T_131; // @[RegisterRouter.scala 59:16]
  assign _T_264 = _T_1112 & _T_257; // @[RegisterRouter.scala 59:16]
  assign _T_280 = _T_192[1:0] == 2'h3; // @[RegisterRouter.scala 59:16]
  assign _T_1181 = _T_1059 & _T_826[24]; // @[RegisterRouter.scala 59:16]
  assign _T_1182 = _T_1181 & _T_131; // @[RegisterRouter.scala 59:16]
  assign _T_287 = _T_1182 & _T_280; // @[RegisterRouter.scala 59:16]
  assign _T_1186 = _T_1059 & _T_826[25]; // @[RegisterRouter.scala 59:16]
  assign _T_1187 = _T_1186 & _T_131; // @[RegisterRouter.scala 59:16]
  assign _T_310 = _T_1187 & _T_280; // @[RegisterRouter.scala 59:16]
  assign _T_1131 = _T_1059 & _T_826[14]; // @[RegisterRouter.scala 59:16]
  assign _T_1132 = _T_1131 & _T_131; // @[RegisterRouter.scala 59:16]
  assign _T_333 = _T_1132 & _T_257; // @[RegisterRouter.scala 59:16]
  assign _T_1161 = _T_1059 & _T_826[20]; // @[RegisterRouter.scala 59:16]
  assign _T_1162 = _T_1161 & _T_131; // @[RegisterRouter.scala 59:16]
  assign _T_356 = _T_1162 & _T_280; // @[RegisterRouter.scala 59:16]
  assign _T_1066 = _T_1059 & _T_826[1]; // @[RegisterRouter.scala 59:16]
  assign _T_1067 = _T_1066 & _T_131; // @[RegisterRouter.scala 59:16]
  assign _T_379 = _T_1067 & _T_192[0]; // @[RegisterRouter.scala 59:16]
  assign _T_1091 = _T_1059 & _T_826[6]; // @[RegisterRouter.scala 59:16]
  assign _T_1092 = _T_1091 & _T_131; // @[RegisterRouter.scala 59:16]
  assign _T_402 = _T_1092 & _T_280; // @[RegisterRouter.scala 59:16]
  assign _T_1166 = _T_1059 & _T_826[21]; // @[RegisterRouter.scala 59:16]
  assign _T_1167 = _T_1166 & _T_131; // @[RegisterRouter.scala 59:16]
  assign _T_425 = _T_1167 & _T_280; // @[RegisterRouter.scala 59:16]
  assign _T_1106 = _T_1059 & _T_826[9]; // @[RegisterRouter.scala 59:16]
  assign _T_1107 = _T_1106 & _T_131; // @[RegisterRouter.scala 59:16]
  assign _T_448 = _T_1107 & _T_280; // @[RegisterRouter.scala 59:16]
  assign _T_1126 = _T_1059 & _T_826[13]; // @[RegisterRouter.scala 59:16]
  assign _T_1127 = _T_1126 & _T_131; // @[RegisterRouter.scala 59:16]
  assign _T_471 = _T_1127 & _T_257; // @[RegisterRouter.scala 59:16]
  assign _T_1071 = _T_1059 & _T_826[2]; // @[RegisterRouter.scala 59:16]
  assign _T_1072 = _T_1071 & _T_131; // @[RegisterRouter.scala 59:16]
  assign _T_494 = _T_1072 & _T_280; // @[RegisterRouter.scala 59:16]
  assign _T_1146 = _T_1059 & _T_826[17]; // @[RegisterRouter.scala 59:16]
  assign _T_1147 = _T_1146 & _T_131; // @[RegisterRouter.scala 59:16]
  assign _T_517 = _T_1147 & _T_257; // @[RegisterRouter.scala 59:16]
  assign _T_1171 = _T_1059 & _T_826[22]; // @[RegisterRouter.scala 59:16]
  assign _T_1172 = _T_1171 & _T_131; // @[RegisterRouter.scala 59:16]
  assign _T_540 = _T_1172 & _T_280; // @[RegisterRouter.scala 59:16]
  assign _T_1121 = _T_1059 & _T_826[12]; // @[RegisterRouter.scala 59:16]
  assign _T_1122 = _T_1121 & _T_131; // @[RegisterRouter.scala 59:16]
  assign _T_563 = _T_1122 & _T_257; // @[RegisterRouter.scala 59:16]
  assign _T_1096 = _T_1059 & _T_826[7]; // @[RegisterRouter.scala 59:16]
  assign _T_1097 = _T_1096 & _T_131; // @[RegisterRouter.scala 59:16]
  assign _T_586 = _T_1097 & _T_280; // @[RegisterRouter.scala 59:16]
  assign _T_602 = _T_192[9:0] == 10'h3ff; // @[RegisterRouter.scala 59:16]
  assign _T_1076 = _T_1059 & _T_826[3]; // @[RegisterRouter.scala 59:16]
  assign _T_1077 = _T_1076 & _T_131; // @[RegisterRouter.scala 59:16]
  assign _T_609 = _T_1077 & _T_602; // @[RegisterRouter.scala 59:16]
  assign _GEN_24 = _T_609 ? _T_2_w_bits_data[9:0] : {{2'd0}, interframeNumOfSamples}; // @[RegField.scala 134:88]
  assign _T_620 = {{2'd0}, interframeNumOfSamples}; // @[RegisterRouter.scala 59:16]
  assign _T_1151 = _T_1059 & _T_826[18]; // @[RegisterRouter.scala 59:16]
  assign _T_1152 = _T_1151 & _T_131; // @[RegisterRouter.scala 59:16]
  assign _T_632 = _T_1152 & _T_280; // @[RegisterRouter.scala 59:16]
  assign _T_1141 = _T_1059 & _T_826[16]; // @[RegisterRouter.scala 59:16]
  assign _T_1142 = _T_1141 & _T_131; // @[RegisterRouter.scala 59:16]
  assign _T_655 = _T_1142 & _T_257; // @[RegisterRouter.scala 59:16]
  assign _T_1116 = _T_1059 & _T_826[11]; // @[RegisterRouter.scala 59:16]
  assign _T_1117 = _T_1116 & _T_131; // @[RegisterRouter.scala 59:16]
  assign _T_678 = _T_1117 & _T_257; // @[RegisterRouter.scala 59:16]
  assign _T_1176 = _T_1059 & _T_826[23]; // @[RegisterRouter.scala 59:16]
  assign _T_1177 = _T_1176 & _T_131; // @[RegisterRouter.scala 59:16]
  assign _T_701 = _T_1177 & _T_280; // @[RegisterRouter.scala 59:16]
  assign _T_1101 = _T_1059 & _T_826[8]; // @[RegisterRouter.scala 59:16]
  assign _T_1102 = _T_1101 & _T_131; // @[RegisterRouter.scala 59:16]
  assign _T_724 = _T_1102 & _T_280; // @[RegisterRouter.scala 59:16]
  assign _T_1156 = _T_1059 & _T_826[19]; // @[RegisterRouter.scala 59:16]
  assign _T_1157 = _T_1156 & _T_131; // @[RegisterRouter.scala 59:16]
  assign _T_747 = _T_1157 & _T_280; // @[RegisterRouter.scala 59:16]
  assign _T_1081 = _T_1059 & _T_826[4]; // @[RegisterRouter.scala 59:16]
  assign _T_1082 = _T_1081 & _T_131; // @[RegisterRouter.scala 59:16]
  assign _T_770 = _T_1082 & _T_257; // @[RegisterRouter.scala 59:16]
  assign _T_1136 = _T_1059 & _T_826[15]; // @[RegisterRouter.scala 59:16]
  assign _T_1137 = _T_1136 & _T_131; // @[RegisterRouter.scala 59:16]
  assign _T_793 = _T_1137 & _T_257; // @[RegisterRouter.scala 59:16]
  assign _GEN_162 = 5'h1 == _T_825 ? _T_131 : _T_131; // @[MuxLiteral.scala 48:10]
  assign _GEN_163 = 5'h2 == _T_825 ? _T_131 : _GEN_162; // @[MuxLiteral.scala 48:10]
  assign _GEN_164 = 5'h3 == _T_825 ? _T_131 : _GEN_163; // @[MuxLiteral.scala 48:10]
  assign _GEN_165 = 5'h4 == _T_825 ? _T_131 : _GEN_164; // @[MuxLiteral.scala 48:10]
  assign _GEN_166 = 5'h5 == _T_825 ? _T_131 : _GEN_165; // @[MuxLiteral.scala 48:10]
  assign _GEN_167 = 5'h6 == _T_825 ? _T_131 : _GEN_166; // @[MuxLiteral.scala 48:10]
  assign _GEN_168 = 5'h7 == _T_825 ? _T_131 : _GEN_167; // @[MuxLiteral.scala 48:10]
  assign _GEN_169 = 5'h8 == _T_825 ? _T_131 : _GEN_168; // @[MuxLiteral.scala 48:10]
  assign _GEN_170 = 5'h9 == _T_825 ? _T_131 : _GEN_169; // @[MuxLiteral.scala 48:10]
  assign _GEN_171 = 5'ha == _T_825 ? _T_131 : _GEN_170; // @[MuxLiteral.scala 48:10]
  assign _GEN_172 = 5'hb == _T_825 ? _T_131 : _GEN_171; // @[MuxLiteral.scala 48:10]
  assign _GEN_173 = 5'hc == _T_825 ? _T_131 : _GEN_172; // @[MuxLiteral.scala 48:10]
  assign _GEN_174 = 5'hd == _T_825 ? _T_131 : _GEN_173; // @[MuxLiteral.scala 48:10]
  assign _GEN_175 = 5'he == _T_825 ? _T_131 : _GEN_174; // @[MuxLiteral.scala 48:10]
  assign _GEN_176 = 5'hf == _T_825 ? _T_131 : _GEN_175; // @[MuxLiteral.scala 48:10]
  assign _GEN_177 = 5'h10 == _T_825 ? _T_131 : _GEN_176; // @[MuxLiteral.scala 48:10]
  assign _GEN_178 = 5'h11 == _T_825 ? _T_131 : _GEN_177; // @[MuxLiteral.scala 48:10]
  assign _GEN_179 = 5'h12 == _T_825 ? _T_131 : _GEN_178; // @[MuxLiteral.scala 48:10]
  assign _GEN_180 = 5'h13 == _T_825 ? _T_131 : _GEN_179; // @[MuxLiteral.scala 48:10]
  assign _GEN_181 = 5'h14 == _T_825 ? _T_131 : _GEN_180; // @[MuxLiteral.scala 48:10]
  assign _GEN_182 = 5'h15 == _T_825 ? _T_131 : _GEN_181; // @[MuxLiteral.scala 48:10]
  assign _GEN_183 = 5'h16 == _T_825 ? _T_131 : _GEN_182; // @[MuxLiteral.scala 48:10]
  assign _GEN_184 = 5'h17 == _T_825 ? _T_131 : _GEN_183; // @[MuxLiteral.scala 48:10]
  assign _GEN_185 = 5'h18 == _T_825 ? _T_131 : _GEN_184; // @[MuxLiteral.scala 48:10]
  assign _GEN_186 = 5'h19 == _T_825 ? _T_131 : _GEN_185; // @[MuxLiteral.scala 48:10]
  assign _GEN_351 = 5'h1a == _T_825; // @[MuxLiteral.scala 48:10]
  assign _GEN_187 = _GEN_351 | _GEN_186; // @[MuxLiteral.scala 48:10]
  assign _GEN_352 = 5'h1b == _T_825; // @[MuxLiteral.scala 48:10]
  assign _GEN_188 = _GEN_352 | _GEN_187; // @[MuxLiteral.scala 48:10]
  assign _GEN_353 = 5'h1c == _T_825; // @[MuxLiteral.scala 48:10]
  assign _GEN_189 = _GEN_353 | _GEN_188; // @[MuxLiteral.scala 48:10]
  assign _GEN_354 = 5'h1d == _T_825; // @[MuxLiteral.scala 48:10]
  assign _GEN_190 = _GEN_354 | _GEN_189; // @[MuxLiteral.scala 48:10]
  assign _GEN_355 = 5'h1e == _T_825; // @[MuxLiteral.scala 48:10]
  assign _GEN_191 = _GEN_355 | _GEN_190; // @[MuxLiteral.scala 48:10]
  assign _GEN_356 = 5'h1f == _T_825; // @[MuxLiteral.scala 48:10]
  assign _GEN_192 = _GEN_356 | _GEN_191; // @[MuxLiteral.scala 48:10]
  assign _T_1564_0 = {{15'd0}, enable}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  assign _T_1564_1 = {{15'd0}, reset_bit}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  assign _GEN_194 = 5'h1 == _T_825 ? _T_1564_1 : _T_1564_0; // @[MuxLiteral.scala 48:10]
  assign _T_1564_2 = {{14'd0}, frameNum}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  assign _GEN_195 = 5'h2 == _T_825 ? _T_1564_2 : _GEN_194; // @[MuxLiteral.scala 48:10]
  assign _T_1564_3 = {{6'd0}, _T_620}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  assign _GEN_196 = 5'h3 == _T_825 ? _T_1564_3 : _GEN_195; // @[MuxLiteral.scala 48:10]
  assign _T_1564_4 = {{13'd0}, differentChirpsNum}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  assign _GEN_197 = 5'h4 == _T_825 ? _T_1564_4 : _GEN_196; // @[MuxLiteral.scala 48:10]
  assign _GEN_198 = 5'h5 == _T_825 ? startingPoint : _GEN_197; // @[MuxLiteral.scala 48:10]
  assign _T_1564_6 = {{14'd0}, segmentNums_0}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  assign _GEN_199 = 5'h6 == _T_825 ? _T_1564_6 : _GEN_198; // @[MuxLiteral.scala 48:10]
  assign _T_1564_7 = {{14'd0}, segmentNums_1}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  assign _GEN_200 = 5'h7 == _T_825 ? _T_1564_7 : _GEN_199; // @[MuxLiteral.scala 48:10]
  assign _T_1564_8 = {{14'd0}, segmentNums_2}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  assign _GEN_201 = 5'h8 == _T_825 ? _T_1564_8 : _GEN_200; // @[MuxLiteral.scala 48:10]
  assign _T_1564_9 = {{14'd0}, segmentNums_3}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  assign _GEN_202 = 5'h9 == _T_825 ? _T_1564_9 : _GEN_201; // @[MuxLiteral.scala 48:10]
  assign _T_1564_10 = {{13'd0}, repeatedChirpNums_0}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  assign _GEN_203 = 5'ha == _T_825 ? _T_1564_10 : _GEN_202; // @[MuxLiteral.scala 48:10]
  assign _T_1564_11 = {{13'd0}, repeatedChirpNums_1}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  assign _GEN_204 = 5'hb == _T_825 ? _T_1564_11 : _GEN_203; // @[MuxLiteral.scala 48:10]
  assign _T_1564_12 = {{13'd0}, repeatedChirpNums_2}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  assign _GEN_205 = 5'hc == _T_825 ? _T_1564_12 : _GEN_204; // @[MuxLiteral.scala 48:10]
  assign _T_1564_13 = {{13'd0}, repeatedChirpNums_3}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  assign _GEN_206 = 5'hd == _T_825 ? _T_1564_13 : _GEN_205; // @[MuxLiteral.scala 48:10]
  assign _T_1564_14 = {{13'd0}, repeatedChirpNums_4}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  assign _GEN_207 = 5'he == _T_825 ? _T_1564_14 : _GEN_206; // @[MuxLiteral.scala 48:10]
  assign _T_1564_15 = {{13'd0}, repeatedChirpNums_5}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  assign _GEN_208 = 5'hf == _T_825 ? _T_1564_15 : _GEN_207; // @[MuxLiteral.scala 48:10]
  assign _T_1564_16 = {{13'd0}, repeatedChirpNums_6}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  assign _GEN_209 = 5'h10 == _T_825 ? _T_1564_16 : _GEN_208; // @[MuxLiteral.scala 48:10]
  assign _T_1564_17 = {{13'd0}, repeatedChirpNums_7}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  assign _GEN_210 = 5'h11 == _T_825 ? _T_1564_17 : _GEN_209; // @[MuxLiteral.scala 48:10]
  assign _T_1564_18 = {{14'd0}, chirpOrdinalNums_0}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  assign _GEN_211 = 5'h12 == _T_825 ? _T_1564_18 : _GEN_210; // @[MuxLiteral.scala 48:10]
  assign _T_1564_19 = {{14'd0}, chirpOrdinalNums_1}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  assign _GEN_212 = 5'h13 == _T_825 ? _T_1564_19 : _GEN_211; // @[MuxLiteral.scala 48:10]
  assign _T_1564_20 = {{14'd0}, chirpOrdinalNums_2}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  assign _GEN_213 = 5'h14 == _T_825 ? _T_1564_20 : _GEN_212; // @[MuxLiteral.scala 48:10]
  assign _T_1564_21 = {{14'd0}, chirpOrdinalNums_3}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  assign _GEN_214 = 5'h15 == _T_825 ? _T_1564_21 : _GEN_213; // @[MuxLiteral.scala 48:10]
  assign _T_1564_22 = {{14'd0}, chirpOrdinalNums_4}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  assign _GEN_215 = 5'h16 == _T_825 ? _T_1564_22 : _GEN_214; // @[MuxLiteral.scala 48:10]
  assign _T_1564_23 = {{14'd0}, chirpOrdinalNums_5}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  assign _GEN_216 = 5'h17 == _T_825 ? _T_1564_23 : _GEN_215; // @[MuxLiteral.scala 48:10]
  assign _T_1564_24 = {{14'd0}, chirpOrdinalNums_6}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  assign _GEN_217 = 5'h18 == _T_825 ? _T_1564_24 : _GEN_216; // @[MuxLiteral.scala 48:10]
  assign _T_1564_25 = {{14'd0}, chirpOrdinalNums_7}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  assign _GEN_218 = 5'h19 == _T_825 ? _T_1564_25 : _GEN_217; // @[MuxLiteral.scala 48:10]
  assign _GEN_219 = 5'h1a == _T_825 ? 16'h0 : _GEN_218; // @[MuxLiteral.scala 48:10]
  assign _GEN_220 = 5'h1b == _T_825 ? 16'h0 : _GEN_219; // @[MuxLiteral.scala 48:10]
  assign _GEN_221 = 5'h1c == _T_825 ? 16'h0 : _GEN_220; // @[MuxLiteral.scala 48:10]
  assign _GEN_222 = 5'h1d == _T_825 ? 16'h0 : _GEN_221; // @[MuxLiteral.scala 48:10]
  assign _GEN_223 = 5'h1e == _T_825 ? 16'h0 : _GEN_222; // @[MuxLiteral.scala 48:10]
  assign _GEN_224 = 5'h1f == _T_825 ? 16'h0 : _GEN_223; // @[MuxLiteral.scala 48:10]
  assign _T_1566 = _GEN_192 ? _GEN_224 : 16'h0; // @[RegisterRouter.scala 59:16]
  assign _T_1567_bits_read = Queue_io_deq_bits_read; // @[Decoupled.scala 308:19 Decoupled.scala 309:14]
  assign _T_2_r_ready = axi4xbar_auto_out_1_r_ready; // @[Nodes.scala 370:76 LazyModule.scala 167:31]
  assign _T_2_b_ready = axi4xbar_auto_out_1_b_ready; // @[Nodes.scala 370:76 LazyModule.scala 167:31]
  assign _T_1567_valid = Queue_io_deq_valid; // @[Decoupled.scala 308:19 Decoupled.scala 310:15]
  assign _T_1570 = ~_T_1567_bits_read; // @[RegisterRouter.scala 65:29]
  assign _GEN_226 = 3'h1 == differentChirpsCounter ? chirpOrdinalNums_1 : chirpOrdinalNums_0; // @[PLFGDspBlockMem.scala 238:18]
  assign _GEN_227 = 3'h2 == differentChirpsCounter ? chirpOrdinalNums_2 : _GEN_226; // @[PLFGDspBlockMem.scala 238:18]
  assign _GEN_228 = 3'h3 == differentChirpsCounter ? chirpOrdinalNums_3 : _GEN_227; // @[PLFGDspBlockMem.scala 238:18]
  assign _GEN_229 = 3'h4 == differentChirpsCounter ? chirpOrdinalNums_4 : _GEN_228; // @[PLFGDspBlockMem.scala 238:18]
  assign _GEN_230 = 3'h5 == differentChirpsCounter ? chirpOrdinalNums_5 : _GEN_229; // @[PLFGDspBlockMem.scala 238:18]
  assign _GEN_231 = 3'h6 == differentChirpsCounter ? chirpOrdinalNums_6 : _GEN_230; // @[PLFGDspBlockMem.scala 238:18]
  assign _GEN_232 = 3'h7 == differentChirpsCounter ? chirpOrdinalNums_7 : _GEN_231; // @[PLFGDspBlockMem.scala 238:18]
  assign _T_1573 = enable & auto_stream_out_ready; // @[PLFGDspBlockMem.scala 239:19]
  assign _T_1574 = ~end_; // @[PLFGDspBlockMem.scala 239:35]
  assign _T_1575 = _T_1573 & _T_1574; // @[PLFGDspBlockMem.scala 239:32]
  assign _T_1577 = samplesCounter + 8'h1; // @[PLFGDspBlockMem.scala 241:30]
  assign _T_1578 = _T_1577 >= numsOfSamples; // @[PLFGDspBlockMem.scala 241:37]
  assign _T_1580 = segmentCounter + 2'h1; // @[PLFGDspBlockMem.scala 242:32]
  assign chirpIndex = reset_bit ? 2'h0 : _GEN_232; // @[PLFGDspBlockMem.scala 224:20]
  assign _GEN_234 = 2'h1 == chirpIndex ? segmentNums_1 : segmentNums_0; // @[PLFGDspBlockMem.scala 242:39]
  assign _GEN_235 = 2'h2 == chirpIndex ? segmentNums_2 : _GEN_234; // @[PLFGDspBlockMem.scala 242:39]
  assign _GEN_236 = 2'h3 == chirpIndex ? segmentNums_3 : _GEN_235; // @[PLFGDspBlockMem.scala 242:39]
  assign _T_1581 = _T_1580 >= _GEN_236; // @[PLFGDspBlockMem.scala 242:39]
  assign _T_1583 = repeatedChirpsCounter + 3'h1; // @[PLFGDspBlockMem.scala 243:41]
  assign _GEN_238 = 3'h1 == differentChirpsCounter ? repeatedChirpNums_1 : repeatedChirpNums_0; // @[PLFGDspBlockMem.scala 243:48]
  assign _GEN_239 = 3'h2 == differentChirpsCounter ? repeatedChirpNums_2 : _GEN_238; // @[PLFGDspBlockMem.scala 243:48]
  assign _GEN_240 = 3'h3 == differentChirpsCounter ? repeatedChirpNums_3 : _GEN_239; // @[PLFGDspBlockMem.scala 243:48]
  assign _GEN_241 = 3'h4 == differentChirpsCounter ? repeatedChirpNums_4 : _GEN_240; // @[PLFGDspBlockMem.scala 243:48]
  assign _GEN_242 = 3'h5 == differentChirpsCounter ? repeatedChirpNums_5 : _GEN_241; // @[PLFGDspBlockMem.scala 243:48]
  assign _GEN_243 = 3'h6 == differentChirpsCounter ? repeatedChirpNums_6 : _GEN_242; // @[PLFGDspBlockMem.scala 243:48]
  assign _GEN_244 = 3'h7 == differentChirpsCounter ? repeatedChirpNums_7 : _GEN_243; // @[PLFGDspBlockMem.scala 243:48]
  assign _T_1584 = _T_1583 >= _GEN_244; // @[PLFGDspBlockMem.scala 243:48]
  assign _T_1586 = differentChirpsCounter + 3'h1; // @[PLFGDspBlockMem.scala 244:44]
  assign _T_1587 = _T_1586 >= differentChirpsNum; // @[PLFGDspBlockMem.scala 244:51]
  assign _T_1590 = frameNum == 2'h0; // @[PLFGDspBlockMem.scala 245:31]
  assign _T_1592 = framePauseCounter + 6'h1; // @[PLFGDspBlockMem.scala 247:43]
  assign _GEN_357 = {{2'd0}, _T_1592}; // @[PLFGDspBlockMem.scala 247:50]
  assign _T_1593 = _GEN_357 >= interframeNumOfSamples; // @[PLFGDspBlockMem.scala 247:50]
  assign _T_1597 = frameCounter + 2'h1; // @[PLFGDspBlockMem.scala 258:38]
  assign _T_1598 = _T_1597 >= frameNum; // @[PLFGDspBlockMem.scala 258:45]
  assign _GEN_257 = _T_1598 | end_; // @[PLFGDspBlockMem.scala 258:57]
  assign _T_1616 = enable2 & auto_stream_out_ready; // @[PLFGDspBlockMem.scala 298:20]
  assign _T_1617 = ~end2; // @[PLFGDspBlockMem.scala 298:36]
  assign _T_1618 = _T_1616 & _T_1617; // @[PLFGDspBlockMem.scala 298:33]
  assign _T_1620 = samplesCounter2 + 8'h1; // @[PLFGDspBlockMem.scala 300:31]
  assign _T_1621 = _T_1620 >= numsOfSamples; // @[PLFGDspBlockMem.scala 300:38]
  assign _T_1623 = segmentCounter2 + 2'h1; // @[PLFGDspBlockMem.scala 301:34]
  assign _GEN_318 = 2'h1 == chirpIndexOld ? segmentNums_1 : segmentNums_0; // @[PLFGDspBlockMem.scala 301:41]
  assign _GEN_319 = 2'h2 == chirpIndexOld ? segmentNums_2 : _GEN_318; // @[PLFGDspBlockMem.scala 301:41]
  assign _GEN_320 = 2'h3 == chirpIndexOld ? segmentNums_3 : _GEN_319; // @[PLFGDspBlockMem.scala 301:41]
  assign _T_1626 = _T_1623 >= _GEN_320; // @[PLFGDspBlockMem.scala 301:41]
  assign _T_1630 = repeatedChirpsCounter2 + 3'h1; // @[PLFGDspBlockMem.scala 303:42]
  assign _T_1631 = _T_1630 >= _GEN_244; // @[PLFGDspBlockMem.scala 303:49]
  assign _T_1633 = differentChirpsCounter2 + 3'h1; // @[PLFGDspBlockMem.scala 304:45]
  assign _T_1634 = _T_1633 >= differentChirpsNum; // @[PLFGDspBlockMem.scala 304:52]
  assign _T_1640 = frameCounter2 >= frameNum; // @[PLFGDspBlockMem.scala 309:38]
  assign _GEN_321 = _T_1640 | end2; // @[PLFGDspBlockMem.scala 309:50]
  assign _T_1652 = dataFromMem[15:0]; // @[PLFGDspBlockMem.scala 326:73]
  assign _T_1655 = $signed(currentVal) + $signed(_T_1652); // @[FixedPointTypeClass.scala 20:58]
  assign _T_1660 = $signed(currentVal) - $signed(_T_1652); // @[FixedPointTypeClass.scala 30:68]
  assign _T_1675 = ~started; // @[PLFGDspBlockMem.scala 337:14]
  assign _GEN_336 = _T_1618 | started; // @[PLFGDspBlockMem.scala 298:42]
  assign _GEN_342 = reset_bit ? startingPoint : currentVal; // @[PLFGDspBlockMem.scala 295:20]
  assign _T_1680 = ~_T_1679; // @[PLFGDspBlockMem.scala 345:31]
  assign _T_1681 = enable2 & _T_1680; // @[PLFGDspBlockMem.scala 345:28]
  assign _T_1683 = ~_T_1682; // @[PLFGDspBlockMem.scala 352:17]
  assign lastOut = end_ & _T_1683; // @[PLFGDspBlockMem.scala 352:14]
  assign _T_1686 = ~_T_1685; // @[PLFGDspBlockMem.scala 357:17]
  assign _T_1687 = end_ & _T_1686; // @[PLFGDspBlockMem.scala 357:14]
  assign _T_1689 = auto_stream_out_ready & _T_1688; // @[PLFGDspBlockMem.scala 359:26]
  assign _GEN_345 = _T_1689 ? 1'h0 : lastOutReg; // @[PLFGDspBlockMem.scala 359:42]
  assign _GEN_346 = _T_1687 | _GEN_345; // @[PLFGDspBlockMem.scala 357:31]
  assign _T_1691 = lastOut | lastOutReg; // @[PLFGDspBlockMem.scala 362:46]
  assign _T_1693 = ~reset_bit; // @[PLFGDspBlockMem.scala 365:10]
  assign _GEN_359 = {{1'd0}, chirpIndex}; // @[UIntTypeClass.scala 39:41]
  assign _T_1694 = _GEN_359 * 3'h4; // @[UIntTypeClass.scala 39:41]
  assign _GEN_360 = {{3'd0}, segmentCounter}; // @[PLFGDspBlockMem.scala 367:57]
  assign _T_1696 = _T_1694 + _GEN_360; // @[PLFGDspBlockMem.scala 367:57]
  assign auto_mem_in_aw_ready = axi4xbar_auto_in_aw_ready; // @[LazyModule.scala 173:31]
  assign auto_mem_in_w_ready = axi4xbar_auto_in_w_ready; // @[LazyModule.scala 173:31]
  assign auto_mem_in_b_valid = axi4xbar_auto_in_b_valid; // @[LazyModule.scala 173:31]
  assign auto_mem_in_b_bits_resp = axi4xbar_auto_in_b_bits_resp; // @[LazyModule.scala 173:31]
  assign auto_mem_in_ar_ready = axi4xbar_auto_in_ar_ready; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_valid = axi4xbar_auto_in_r_valid; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_bits_data = axi4xbar_auto_in_r_bits_data; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_bits_resp = axi4xbar_auto_in_r_bits_resp; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_bits_last = axi4xbar_auto_in_r_bits_last; // @[LazyModule.scala 173:31]
  assign auto_stream_out_valid = auto_stream_out_ready ? _T_1681 : auto_stream_out_ready; // @[LazyModule.scala 173:49]
  assign auto_stream_out_bits_data = {{16'd0}, _GEN_342}; // @[LazyModule.scala 173:49]
  assign auto_stream_out_bits_last = auto_stream_out_ready & _T_1691; // @[LazyModule.scala 173:49]
  assign axi4xbar_clock = clock;
  assign axi4xbar_reset = reset;
  assign axi4xbar_auto_in_aw_valid = auto_mem_in_aw_valid; // @[LazyModule.scala 167:57]
  assign axi4xbar_auto_in_aw_bits_id = auto_mem_in_aw_bits_id; // @[LazyModule.scala 167:57]
  assign axi4xbar_auto_in_aw_bits_addr = auto_mem_in_aw_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4xbar_auto_in_w_valid = auto_mem_in_w_valid; // @[LazyModule.scala 167:57]
  assign axi4xbar_auto_in_w_bits_data = auto_mem_in_w_bits_data; // @[LazyModule.scala 167:57]
  assign axi4xbar_auto_in_w_bits_strb = auto_mem_in_w_bits_strb; // @[LazyModule.scala 167:57]
  assign axi4xbar_auto_in_w_bits_last = auto_mem_in_w_bits_last; // @[LazyModule.scala 167:57]
  assign axi4xbar_auto_in_b_ready = auto_mem_in_b_ready; // @[LazyModule.scala 167:57]
  assign axi4xbar_auto_in_ar_valid = auto_mem_in_ar_valid; // @[LazyModule.scala 167:57]
  assign axi4xbar_auto_in_ar_bits_id = auto_mem_in_ar_bits_id; // @[LazyModule.scala 167:57]
  assign axi4xbar_auto_in_ar_bits_addr = auto_mem_in_ar_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4xbar_auto_in_ar_bits_size = auto_mem_in_ar_bits_size; // @[LazyModule.scala 167:57]
  assign axi4xbar_auto_in_r_ready = auto_mem_in_r_ready; // @[LazyModule.scala 167:57]
  assign axi4xbar_auto_out_1_aw_ready = _T_75 & _T_2_w_valid; // @[LazyModule.scala 167:31]
  assign axi4xbar_auto_out_1_w_ready = _T_75 & _T_2_aw_valid; // @[LazyModule.scala 167:31]
  assign axi4xbar_auto_out_1_b_valid = _T_1567_valid & _T_1570; // @[LazyModule.scala 167:31]
  assign axi4xbar_auto_out_1_b_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 167:31]
  assign axi4xbar_auto_out_1_ar_ready = Queue_io_enq_ready; // @[LazyModule.scala 167:31]
  assign axi4xbar_auto_out_1_r_valid = _T_1567_valid & _T_1567_bits_read; // @[LazyModule.scala 167:31]
  assign axi4xbar_auto_out_1_r_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 167:31]
  assign axi4xbar_auto_out_1_r_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 167:31]
  assign axi4xbar_auto_out_0_aw_ready = ramIn1_w_valid & _T_6; // @[LazyModule.scala 167:31]
  assign axi4xbar_auto_out_0_w_ready = ramIn1_aw_valid & _T_6; // @[LazyModule.scala 167:31]
  assign axi4xbar_auto_out_0_b_valid = w_full1; // @[LazyModule.scala 167:31]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = _T_2_ar_valid | _T_72; // @[Decoupled.scala 288:22]
  assign Queue_io_enq_bits_read = axi4xbar_auto_out_1_ar_valid; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_data = {{16'd0}, _T_1566}; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_extra = _T_2_ar_valid ? _T_2_ar_bits_id : _T_2_aw_bits_id; // @[Decoupled.scala 289:21]
  assign Queue_io_deq_ready = _T_1567_bits_read ? _T_2_r_ready : _T_2_b_ready; // @[Decoupled.scala 311:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    configParamsMem1[initvar] = _RAND_0[25:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  configParamsMem1__T_64_en_pipe_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  configParamsMem1__T_64_addr_pipe_0 = _RAND_2[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  w_full1 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  enable = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  reset_bit = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  frameNum = _RAND_6[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  startingPoint = _RAND_7[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  interframeNumOfSamples = _RAND_8[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  differentChirpsNum = _RAND_9[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  currentVal = _RAND_10[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  samplesCounter = _RAND_11[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  segmentCounter = _RAND_12[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  frameCounter = _RAND_13[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  framePauseCounter = _RAND_14[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  end_ = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  samplesCounter2 = _RAND_16[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  segmentCounter2 = _RAND_17[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  frameCounter2 = _RAND_18[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  end2 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  repeatedChirpsCounter = _RAND_20[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  differentChirpsCounter = _RAND_21[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_19 = _RAND_22[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  repeatedChirpsCounter2 = _RAND_23[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_20 = _RAND_24[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  differentChirpsCounter2 = _RAND_25[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  segmentNums_0 = _RAND_26[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  segmentNums_1 = _RAND_27[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  segmentNums_2 = _RAND_28[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  segmentNums_3 = _RAND_29[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  repeatedChirpNums_0 = _RAND_30[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  repeatedChirpNums_1 = _RAND_31[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  repeatedChirpNums_2 = _RAND_32[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  repeatedChirpNums_3 = _RAND_33[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  repeatedChirpNums_4 = _RAND_34[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  repeatedChirpNums_5 = _RAND_35[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  repeatedChirpNums_6 = _RAND_36[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  repeatedChirpNums_7 = _RAND_37[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  chirpOrdinalNums_0 = _RAND_38[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  chirpOrdinalNums_1 = _RAND_39[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  chirpOrdinalNums_2 = _RAND_40[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  chirpOrdinalNums_3 = _RAND_41[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  chirpOrdinalNums_4 = _RAND_42[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  chirpOrdinalNums_5 = _RAND_43[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  chirpOrdinalNums_6 = _RAND_44[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  chirpOrdinalNums_7 = _RAND_45[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  enable2 = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  chirpIndexOld = _RAND_47[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  started = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  _T_1679 = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  lastOutReg = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  _T_1682 = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  _T_1685 = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  _T_1688 = _RAND_53[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(configParamsMem1__T_14_en & configParamsMem1__T_14_mask) begin
      configParamsMem1[configParamsMem1__T_14_addr] <= configParamsMem1__T_14_data; // @[PLFGDspBlockMem.scala 110:39]
    end
    configParamsMem1__T_64_en_pipe_0 <= 1'h1;
    if (_T_1693) begin
      if (enable) begin
        configParamsMem1__T_64_addr_pipe_0 <= _T_1696[3:0];
      end else begin
        configParamsMem1__T_64_addr_pipe_0 <= 4'h0;
      end
    end else begin
      configParamsMem1__T_64_addr_pipe_0 <= 4'h0;
    end
    if (reset) begin
      w_full1 <= 1'h0;
    end else begin
      w_full1 <= _GEN_1;
    end
    if (reset) begin
      enable <= 1'h0;
    end else if (_T_218) begin
      enable <= _T_2_w_bits_data[0];
    end
    if (reset) begin
      reset_bit <= 1'h0;
    end else if (_T_379) begin
      reset_bit <= _T_2_w_bits_data[0];
    end
    if (reset) begin
      frameNum <= 2'h1;
    end else if (_T_494) begin
      frameNum <= _T_2_w_bits_data[1:0];
    end
    if (reset) begin
      startingPoint <= 16'h0;
    end else if (_T_241) begin
      startingPoint <= _T_2_w_bits_data[15:0];
    end
    if (reset) begin
      interframeNumOfSamples <= 8'h0;
    end else begin
      interframeNumOfSamples <= _GEN_24[7:0];
    end
    if (reset) begin
      differentChirpsNum <= 3'h1;
    end else if (_T_770) begin
      differentChirpsNum <= _T_2_w_bits_data[2:0];
    end
    if (reset) begin
      currentVal <= startingPoint;
    end else if (reset_bit) begin
      currentVal <= startingPoint;
    end else if (_T_1618) begin
      if (_T_1621) begin
        if (_T_1626) begin
          if (_T_1631) begin
            if (_T_1634) begin
              if (_T_1590) begin
                currentVal <= startingPoint;
              end else if (_T_1640) begin
                currentVal <= startingPoint;
              end else begin
                currentVal <= startingPoint;
              end
            end else begin
              currentVal <= startingPoint;
            end
          end else begin
            currentVal <= startingPoint;
          end
        end else if (segmentResets) begin
          currentVal <= startingPoint;
        end else if (slopeSigns) begin
          currentVal <= _T_1655;
        end else begin
          currentVal <= _T_1660;
        end
      end else if (segmentResets) begin
        currentVal <= startingPoint;
      end else if (slopeSigns) begin
        currentVal <= _T_1655;
      end else begin
        currentVal <= _T_1660;
      end
    end else if (_T_1675) begin
      currentVal <= startingPoint;
    end
    if (reset) begin
      samplesCounter <= 8'h0;
    end else if (reset_bit) begin
      samplesCounter <= 8'h0;
    end else if (_T_1575) begin
      if (_T_1578) begin
        if (_T_1581) begin
          if (_T_1584) begin
            if (_T_1587) begin
              if (_T_1590) begin
                if (_T_1593) begin
                  samplesCounter <= 8'h0;
                end
              end else if (!(_T_1598)) begin
                if (_T_1593) begin
                  samplesCounter <= 8'h0;
                end
              end
            end else begin
              samplesCounter <= 8'h0;
            end
          end else begin
            samplesCounter <= 8'h0;
          end
        end else begin
          samplesCounter <= 8'h0;
        end
      end else begin
        samplesCounter <= _T_1577;
      end
    end
    if (reset) begin
      segmentCounter <= 2'h0;
    end else if (reset_bit) begin
      segmentCounter <= 2'h0;
    end else if (_T_1575) begin
      if (_T_1578) begin
        if (_T_1581) begin
          if (_T_1584) begin
            if (_T_1587) begin
              if (_T_1590) begin
                if (_T_1593) begin
                  segmentCounter <= 2'h0;
                end
              end else if (!(_T_1598)) begin
                if (_T_1593) begin
                  segmentCounter <= 2'h0;
                end
              end
            end else begin
              segmentCounter <= 2'h0;
            end
          end else begin
            segmentCounter <= 2'h0;
          end
        end else begin
          segmentCounter <= _T_1580;
        end
      end
    end
    if (reset) begin
      frameCounter <= 2'h0;
    end else if (reset_bit) begin
      frameCounter <= 2'h0;
    end else if (_T_1575) begin
      if (_T_1578) begin
        if (_T_1581) begin
          if (_T_1584) begin
            if (_T_1587) begin
              if (_T_1590) begin
                if (_T_1593) begin
                  frameCounter <= 2'h0;
                end
              end else if (!(_T_1598)) begin
                if (_T_1593) begin
                  frameCounter <= _T_1597;
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      framePauseCounter <= 6'h0;
    end else if (reset_bit) begin
      framePauseCounter <= 6'h0;
    end else if (_T_1575) begin
      if (_T_1578) begin
        if (_T_1581) begin
          if (_T_1584) begin
            if (_T_1587) begin
              if (_T_1590) begin
                if (_T_1593) begin
                  framePauseCounter <= 6'h0;
                end else begin
                  framePauseCounter <= _T_1592;
                end
              end else if (!(_T_1598)) begin
                if (_T_1593) begin
                  framePauseCounter <= 6'h0;
                end else begin
                  framePauseCounter <= _T_1592;
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      end_ <= 1'h0;
    end else if (!(reset_bit)) begin
      if (_T_1575) begin
        if (_T_1578) begin
          if (_T_1581) begin
            if (_T_1584) begin
              if (_T_1587) begin
                if (_T_1590) begin
                  end_ <= 1'h0;
                end else begin
                  end_ <= _GEN_257;
                end
              end
            end
          end
        end
      end
    end
    samplesCounter2 <= samplesCounter;
    segmentCounter2 <= segmentCounter;
    frameCounter2 <= frameCounter;
    if (reset) begin
      end2 <= 1'h0;
    end else if (!(reset_bit)) begin
      if (_T_1618) begin
        if (_T_1621) begin
          if (_T_1626) begin
            if (_T_1631) begin
              if (_T_1634) begin
                if (_T_1590) begin
                  end2 <= 1'h0;
                end else begin
                  end2 <= _GEN_321;
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      repeatedChirpsCounter <= 3'h0;
    end else if (reset_bit) begin
      repeatedChirpsCounter <= 3'h0;
    end else if (_T_1575) begin
      if (_T_1578) begin
        if (_T_1581) begin
          if (_T_1584) begin
            if (_T_1587) begin
              if (_T_1590) begin
                if (_T_1593) begin
                  repeatedChirpsCounter <= 3'h0;
                end
              end else if (!(_T_1598)) begin
                if (_T_1593) begin
                  repeatedChirpsCounter <= 3'h0;
                end
              end
            end else begin
              repeatedChirpsCounter <= 3'h0;
            end
          end else begin
            repeatedChirpsCounter <= _T_1583;
          end
        end
      end
    end
    if (reset) begin
      differentChirpsCounter <= 3'h0;
    end else if (reset_bit) begin
      differentChirpsCounter <= 3'h0;
    end else if (_T_1575) begin
      if (_T_1578) begin
        if (_T_1581) begin
          if (_T_1584) begin
            if (_T_1587) begin
              if (_T_1590) begin
                if (_T_1593) begin
                  differentChirpsCounter <= 3'h0;
                end
              end else if (!(_T_1598)) begin
                if (_T_1593) begin
                  differentChirpsCounter <= 3'h0;
                end
              end
            end else begin
              differentChirpsCounter <= _T_1586;
            end
          end
        end
      end
    end
    _T_19 <= repeatedChirpsCounter;
    repeatedChirpsCounter2 <= _T_19;
    _T_20 <= differentChirpsCounter;
    differentChirpsCounter2 <= _T_20;
    if (reset) begin
      segmentNums_0 <= 2'h0;
    end else if (_T_402) begin
      segmentNums_0 <= _T_2_w_bits_data[1:0];
    end
    if (reset) begin
      segmentNums_1 <= 2'h0;
    end else if (_T_586) begin
      segmentNums_1 <= _T_2_w_bits_data[1:0];
    end
    if (reset) begin
      segmentNums_2 <= 2'h0;
    end else if (_T_724) begin
      segmentNums_2 <= _T_2_w_bits_data[1:0];
    end
    if (reset) begin
      segmentNums_3 <= 2'h0;
    end else if (_T_448) begin
      segmentNums_3 <= _T_2_w_bits_data[1:0];
    end
    if (reset) begin
      repeatedChirpNums_0 <= 3'h0;
    end else if (_T_264) begin
      repeatedChirpNums_0 <= _T_2_w_bits_data[2:0];
    end
    if (reset) begin
      repeatedChirpNums_1 <= 3'h0;
    end else if (_T_678) begin
      repeatedChirpNums_1 <= _T_2_w_bits_data[2:0];
    end
    if (reset) begin
      repeatedChirpNums_2 <= 3'h0;
    end else if (_T_563) begin
      repeatedChirpNums_2 <= _T_2_w_bits_data[2:0];
    end
    if (reset) begin
      repeatedChirpNums_3 <= 3'h0;
    end else if (_T_471) begin
      repeatedChirpNums_3 <= _T_2_w_bits_data[2:0];
    end
    if (reset) begin
      repeatedChirpNums_4 <= 3'h0;
    end else if (_T_333) begin
      repeatedChirpNums_4 <= _T_2_w_bits_data[2:0];
    end
    if (reset) begin
      repeatedChirpNums_5 <= 3'h0;
    end else if (_T_793) begin
      repeatedChirpNums_5 <= _T_2_w_bits_data[2:0];
    end
    if (reset) begin
      repeatedChirpNums_6 <= 3'h0;
    end else if (_T_655) begin
      repeatedChirpNums_6 <= _T_2_w_bits_data[2:0];
    end
    if (reset) begin
      repeatedChirpNums_7 <= 3'h0;
    end else if (_T_517) begin
      repeatedChirpNums_7 <= _T_2_w_bits_data[2:0];
    end
    if (reset) begin
      chirpOrdinalNums_0 <= 2'h0;
    end else if (_T_632) begin
      chirpOrdinalNums_0 <= _T_2_w_bits_data[1:0];
    end
    if (reset) begin
      chirpOrdinalNums_1 <= 2'h0;
    end else if (_T_747) begin
      chirpOrdinalNums_1 <= _T_2_w_bits_data[1:0];
    end
    if (reset) begin
      chirpOrdinalNums_2 <= 2'h0;
    end else if (_T_356) begin
      chirpOrdinalNums_2 <= _T_2_w_bits_data[1:0];
    end
    if (reset) begin
      chirpOrdinalNums_3 <= 2'h0;
    end else if (_T_425) begin
      chirpOrdinalNums_3 <= _T_2_w_bits_data[1:0];
    end
    if (reset) begin
      chirpOrdinalNums_4 <= 2'h0;
    end else if (_T_540) begin
      chirpOrdinalNums_4 <= _T_2_w_bits_data[1:0];
    end
    if (reset) begin
      chirpOrdinalNums_5 <= 2'h0;
    end else if (_T_701) begin
      chirpOrdinalNums_5 <= _T_2_w_bits_data[1:0];
    end
    if (reset) begin
      chirpOrdinalNums_6 <= 2'h0;
    end else if (_T_287) begin
      chirpOrdinalNums_6 <= _T_2_w_bits_data[1:0];
    end
    if (reset) begin
      chirpOrdinalNums_7 <= 2'h0;
    end else if (_T_310) begin
      chirpOrdinalNums_7 <= _T_2_w_bits_data[1:0];
    end
    enable2 <= enable;
    if (reset_bit) begin
      chirpIndexOld <= 2'h0;
    end else if (3'h7 == differentChirpsCounter) begin
      chirpIndexOld <= chirpOrdinalNums_7;
    end else if (3'h6 == differentChirpsCounter) begin
      chirpIndexOld <= chirpOrdinalNums_6;
    end else if (3'h5 == differentChirpsCounter) begin
      chirpIndexOld <= chirpOrdinalNums_5;
    end else if (3'h4 == differentChirpsCounter) begin
      chirpIndexOld <= chirpOrdinalNums_4;
    end else if (3'h3 == differentChirpsCounter) begin
      chirpIndexOld <= chirpOrdinalNums_3;
    end else if (3'h2 == differentChirpsCounter) begin
      chirpIndexOld <= chirpOrdinalNums_2;
    end else if (3'h1 == differentChirpsCounter) begin
      chirpIndexOld <= chirpOrdinalNums_1;
    end else begin
      chirpIndexOld <= chirpOrdinalNums_0;
    end
    if (reset) begin
      started <= 1'h0;
    end else if (!(reset_bit)) begin
      started <= _GEN_336;
    end
    _T_1679 <= end_;
    if (reset) begin
      lastOutReg <= 1'h0;
    end else begin
      lastOutReg <= _GEN_346;
    end
    _T_1682 <= end_;
    _T_1685 <= end_;
    _T_1688 <= end_;
  end
endmodule
module AXI4Splitter_1(
  input         clock,
  input         reset,
  output        auto_mem_in_aw_ready,
  input         auto_mem_in_aw_valid,
  input         auto_mem_in_aw_bits_id,
  input  [29:0] auto_mem_in_aw_bits_addr,
  output        auto_mem_in_w_ready,
  input         auto_mem_in_w_valid,
  input  [31:0] auto_mem_in_w_bits_data,
  input  [3:0]  auto_mem_in_w_bits_strb,
  input         auto_mem_in_b_ready,
  output        auto_mem_in_b_valid,
  output        auto_mem_in_b_bits_id,
  output        auto_mem_in_ar_ready,
  input         auto_mem_in_ar_valid,
  input         auto_mem_in_ar_bits_id,
  input  [29:0] auto_mem_in_ar_bits_addr,
  input  [2:0]  auto_mem_in_ar_bits_size,
  input         auto_mem_in_r_ready,
  output        auto_mem_in_r_valid,
  output        auto_mem_in_r_bits_id,
  output [31:0] auto_mem_in_r_bits_data,
  output        auto_stream_in_ready,
  input         auto_stream_in_valid,
  input  [31:0] auto_stream_in_bits_data,
  input         auto_stream_in_bits_last,
  input         auto_stream_out_1_ready,
  output        auto_stream_out_1_valid,
  output [31:0] auto_stream_out_1_bits_data,
  output        auto_stream_out_1_bits_last,
  input         auto_stream_out_0_ready,
  output        auto_stream_out_0_valid,
  output [31:0] auto_stream_out_0_bits_data,
  output        auto_stream_out_0_bits_last
);
  wire  Queue_clock; // @[Decoupled.scala 287:21]
  wire  Queue_reset; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_read; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_enq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_extra; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_read; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_deq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_extra; // @[Decoupled.scala 287:21]
  reg [31:0] ctrlReg; // @[Splitter.scala 27:26]
  reg [31:0] _RAND_0;
  reg [31:0] maskReg; // @[Splitter.scala 28:26]
  reg [31:0] _RAND_1;
  wire  _T_4; // @[RegisterRouter.scala 40:39]
  wire  _T_5; // @[RegisterRouter.scala 40:26]
  wire  _T_6; // @[RegisterRouter.scala 42:29]
  wire  _T_49_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 290:17]
  wire [29:0] _T_13; // @[RegisterRouter.scala 48:19]
  wire [1:0] _T_53; // @[RegisterRouter.scala 59:16]
  wire  _T_55; // @[RegisterRouter.scala 59:16]
  wire  _T_7; // @[RegisterRouter.scala 42:26]
  wire [1:0] _T_16; // @[OneHot.scala 65:12]
  wire [1:0] _T_18; // @[Misc.scala 200:81]
  wire  _T_19; // @[Misc.scala 204:21]
  wire  _T_22; // @[Misc.scala 209:20]
  wire  _T_24; // @[Misc.scala 213:38]
  wire  _T_25; // @[Misc.scala 213:29]
  wire  _T_27; // @[Misc.scala 213:38]
  wire  _T_28; // @[Misc.scala 213:29]
  wire  _T_31; // @[Misc.scala 209:20]
  wire  _T_32; // @[Misc.scala 212:27]
  wire  _T_33; // @[Misc.scala 213:38]
  wire  _T_34; // @[Misc.scala 213:29]
  wire  _T_35; // @[Misc.scala 212:27]
  wire  _T_36; // @[Misc.scala 213:38]
  wire  _T_37; // @[Misc.scala 213:29]
  wire  _T_38; // @[Misc.scala 212:27]
  wire  _T_39; // @[Misc.scala 213:38]
  wire  _T_40; // @[Misc.scala 213:29]
  wire  _T_41; // @[Misc.scala 212:27]
  wire  _T_42; // @[Misc.scala 213:38]
  wire  _T_43; // @[Misc.scala 213:29]
  wire [3:0] _T_46; // @[Cat.scala 29:58]
  wire [3:0] _T_48; // @[RegisterRouter.scala 54:25]
  wire [7:0] _T_67; // @[Bitwise.scala 72:12]
  wire [7:0] _T_69; // @[Bitwise.scala 72:12]
  wire [7:0] _T_71; // @[Bitwise.scala 72:12]
  wire [7:0] _T_73; // @[Bitwise.scala 72:12]
  wire [31:0] _T_76; // @[Cat.scala 29:58]
  wire  _T_95; // @[RegisterRouter.scala 59:16]
  wire  _T_148; // @[RegisterRouter.scala 59:16]
  wire [1:0] _T_142; // @[OneHot.scala 58:35]
  wire  _T_165; // @[RegisterRouter.scala 59:16]
  wire  _T_172; // @[RegisterRouter.scala 59:16]
  wire  _T_173; // @[RegisterRouter.scala 59:16]
  wire  _T_102; // @[RegisterRouter.scala 59:16]
  wire  _T_167; // @[RegisterRouter.scala 59:16]
  wire  _T_168; // @[RegisterRouter.scala 59:16]
  wire  _T_125; // @[RegisterRouter.scala 59:16]
  wire  _GEN_11; // @[MuxLiteral.scala 48:10]
  wire [31:0] _GEN_13; // @[MuxLiteral.scala 48:10]
  wire  _T_223_bits_read; // @[Decoupled.scala 308:19 Decoupled.scala 309:14]
  wire  _T_223_valid; // @[Decoupled.scala 308:19 Decoupled.scala 310:15]
  wire  _T_226; // @[RegisterRouter.scala 65:29]
  wire  readyOR; // @[Splitter.scala 45:34]
  wire  readyAND; // @[Splitter.scala 46:34]
  wire  _T_229; // @[Splitter.scala 49:19]
  wire  _T_230; // @[Splitter.scala 52:24]
  wire  _GEN_14; // @[Splitter.scala 52:33]
  wire  _T_233; // @[Splitter.scala 62:34]
  wire  _T_237; // @[Splitter.scala 62:34]
  Queue Queue ( // @[Decoupled.scala 287:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_read(Queue_io_enq_bits_read),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_extra(Queue_io_enq_bits_extra),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_read(Queue_io_deq_bits_read),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_extra(Queue_io_deq_bits_extra)
  );
  assign _T_4 = auto_mem_in_aw_valid & auto_mem_in_w_valid; // @[RegisterRouter.scala 40:39]
  assign _T_5 = auto_mem_in_ar_valid | _T_4; // @[RegisterRouter.scala 40:26]
  assign _T_6 = ~auto_mem_in_ar_valid; // @[RegisterRouter.scala 42:29]
  assign _T_49_ready = Queue_io_enq_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 290:17]
  assign _T_13 = auto_mem_in_ar_valid ? auto_mem_in_ar_bits_addr : auto_mem_in_aw_bits_addr; // @[RegisterRouter.scala 48:19]
  assign _T_53 = _T_13[3:2] & 2'h2; // @[RegisterRouter.scala 59:16]
  assign _T_55 = _T_53 == 2'h0; // @[RegisterRouter.scala 59:16]
  assign _T_7 = _T_49_ready & _T_6; // @[RegisterRouter.scala 42:26]
  assign _T_16 = 2'h1 << auto_mem_in_ar_bits_size[0]; // @[OneHot.scala 65:12]
  assign _T_18 = _T_16 | 2'h1; // @[Misc.scala 200:81]
  assign _T_19 = auto_mem_in_ar_bits_size >= 3'h2; // @[Misc.scala 204:21]
  assign _T_22 = ~auto_mem_in_ar_bits_addr[1]; // @[Misc.scala 209:20]
  assign _T_24 = _T_18[1] & _T_22; // @[Misc.scala 213:38]
  assign _T_25 = _T_19 | _T_24; // @[Misc.scala 213:29]
  assign _T_27 = _T_18[1] & auto_mem_in_ar_bits_addr[1]; // @[Misc.scala 213:38]
  assign _T_28 = _T_19 | _T_27; // @[Misc.scala 213:29]
  assign _T_31 = ~auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 209:20]
  assign _T_32 = _T_22 & _T_31; // @[Misc.scala 212:27]
  assign _T_33 = _T_18[0] & _T_32; // @[Misc.scala 213:38]
  assign _T_34 = _T_25 | _T_33; // @[Misc.scala 213:29]
  assign _T_35 = _T_22 & auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  assign _T_36 = _T_18[0] & _T_35; // @[Misc.scala 213:38]
  assign _T_37 = _T_25 | _T_36; // @[Misc.scala 213:29]
  assign _T_38 = auto_mem_in_ar_bits_addr[1] & _T_31; // @[Misc.scala 212:27]
  assign _T_39 = _T_18[0] & _T_38; // @[Misc.scala 213:38]
  assign _T_40 = _T_28 | _T_39; // @[Misc.scala 213:29]
  assign _T_41 = auto_mem_in_ar_bits_addr[1] & auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  assign _T_42 = _T_18[0] & _T_41; // @[Misc.scala 213:38]
  assign _T_43 = _T_28 | _T_42; // @[Misc.scala 213:29]
  assign _T_46 = {_T_43,_T_40,_T_37,_T_34}; // @[Cat.scala 29:58]
  assign _T_48 = auto_mem_in_ar_valid ? _T_46 : auto_mem_in_w_bits_strb; // @[RegisterRouter.scala 54:25]
  assign _T_67 = _T_48[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_69 = _T_48[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_71 = _T_48[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_73 = _T_48[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_76 = {_T_73,_T_71,_T_69,_T_67}; // @[Cat.scala 29:58]
  assign _T_95 = _T_76 == 32'hffffffff; // @[RegisterRouter.scala 59:16]
  assign _T_148 = _T_5 & _T_49_ready; // @[RegisterRouter.scala 59:16]
  assign _T_142 = 2'h1 << _T_13[2]; // @[OneHot.scala 58:35]
  assign _T_165 = _T_148 & _T_6; // @[RegisterRouter.scala 59:16]
  assign _T_172 = _T_165 & _T_142[1]; // @[RegisterRouter.scala 59:16]
  assign _T_173 = _T_172 & _T_55; // @[RegisterRouter.scala 59:16]
  assign _T_102 = _T_173 & _T_95; // @[RegisterRouter.scala 59:16]
  assign _T_167 = _T_165 & _T_142[0]; // @[RegisterRouter.scala 59:16]
  assign _T_168 = _T_167 & _T_55; // @[RegisterRouter.scala 59:16]
  assign _T_125 = _T_168 & _T_95; // @[RegisterRouter.scala 59:16]
  assign _GEN_11 = _T_13[2] ? _T_55 : _T_55; // @[MuxLiteral.scala 48:10]
  assign _GEN_13 = _T_13[2] ? maskReg : ctrlReg; // @[MuxLiteral.scala 48:10]
  assign _T_223_bits_read = Queue_io_deq_bits_read; // @[Decoupled.scala 308:19 Decoupled.scala 309:14]
  assign _T_223_valid = Queue_io_deq_valid; // @[Decoupled.scala 308:19 Decoupled.scala 310:15]
  assign _T_226 = ~_T_223_bits_read; // @[RegisterRouter.scala 65:29]
  assign readyOR = auto_stream_out_0_ready | auto_stream_out_1_ready; // @[Splitter.scala 45:34]
  assign readyAND = auto_stream_out_0_ready & auto_stream_out_1_ready; // @[Splitter.scala 46:34]
  assign _T_229 = ctrlReg == 32'h0; // @[Splitter.scala 49:19]
  assign _T_230 = ctrlReg == 32'h1; // @[Splitter.scala 52:24]
  assign _GEN_14 = _T_230 & readyOR; // @[Splitter.scala 52:33]
  assign _T_233 = ~maskReg[0]; // @[Splitter.scala 62:34]
  assign _T_237 = ~maskReg[1]; // @[Splitter.scala 62:34]
  assign auto_mem_in_aw_ready = _T_7 & auto_mem_in_w_valid; // @[LazyModule.scala 173:31]
  assign auto_mem_in_w_ready = _T_7 & auto_mem_in_aw_valid; // @[LazyModule.scala 173:31]
  assign auto_mem_in_b_valid = _T_223_valid & _T_226; // @[LazyModule.scala 173:31]
  assign auto_mem_in_b_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_mem_in_ar_ready = Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_valid = _T_223_valid & _T_223_bits_read; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 173:31]
  assign auto_stream_in_ready = _T_229 ? readyAND : _GEN_14; // @[LazyModule.scala 173:31]
  assign auto_stream_out_1_valid = auto_stream_in_valid & _T_237; // @[LazyModule.scala 173:49]
  assign auto_stream_out_1_bits_data = auto_stream_in_bits_data; // @[LazyModule.scala 173:49]
  assign auto_stream_out_1_bits_last = auto_stream_in_bits_last; // @[LazyModule.scala 173:49]
  assign auto_stream_out_0_valid = auto_stream_in_valid & _T_233; // @[LazyModule.scala 173:49]
  assign auto_stream_out_0_bits_data = auto_stream_in_bits_data; // @[LazyModule.scala 173:49]
  assign auto_stream_out_0_bits_last = auto_stream_in_bits_last; // @[LazyModule.scala 173:49]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_mem_in_ar_valid | _T_4; // @[Decoupled.scala 288:22]
  assign Queue_io_enq_bits_read = auto_mem_in_ar_valid; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_data = _GEN_11 ? _GEN_13 : 32'h0; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_extra = auto_mem_in_ar_valid ? auto_mem_in_ar_bits_id : auto_mem_in_aw_bits_id; // @[Decoupled.scala 289:21]
  assign Queue_io_deq_ready = _T_223_bits_read ? auto_mem_in_r_ready : auto_mem_in_b_ready; // @[Decoupled.scala 311:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ctrlReg = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  maskReg = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      ctrlReg <= 32'h0;
    end else if (_T_125) begin
      ctrlReg <= auto_mem_in_w_bits_data;
    end
    if (reset) begin
      maskReg <= 32'h0;
    end else if (_T_102) begin
      maskReg <= auto_mem_in_w_bits_data;
    end
  end
endmodule
module AXI4StreamMux(
  input         clock,
  input         reset,
  output        auto_register_in_aw_ready,
  input         auto_register_in_aw_valid,
  input         auto_register_in_aw_bits_id,
  input  [29:0] auto_register_in_aw_bits_addr,
  output        auto_register_in_w_ready,
  input         auto_register_in_w_valid,
  input  [31:0] auto_register_in_w_bits_data,
  input  [3:0]  auto_register_in_w_bits_strb,
  input         auto_register_in_b_ready,
  output        auto_register_in_b_valid,
  output        auto_register_in_b_bits_id,
  output        auto_register_in_ar_ready,
  input         auto_register_in_ar_valid,
  input         auto_register_in_ar_bits_id,
  input  [29:0] auto_register_in_ar_bits_addr,
  input  [2:0]  auto_register_in_ar_bits_size,
  input         auto_register_in_r_ready,
  output        auto_register_in_r_valid,
  output        auto_register_in_r_bits_id,
  output [31:0] auto_register_in_r_bits_data,
  output        auto_stream_in_2_ready,
  input         auto_stream_in_2_valid,
  input  [31:0] auto_stream_in_2_bits_data,
  input         auto_stream_in_2_bits_last,
  output        auto_stream_in_1_ready,
  input         auto_stream_in_1_valid,
  input  [31:0] auto_stream_in_1_bits_data,
  input         auto_stream_in_1_bits_last,
  output        auto_stream_in_0_ready,
  input         auto_stream_in_0_valid,
  input  [31:0] auto_stream_in_0_bits_data,
  input         auto_stream_in_0_bits_last,
  input         auto_stream_out_0_ready,
  output        auto_stream_out_0_valid,
  output [31:0] auto_stream_out_0_bits_data,
  output        auto_stream_out_0_bits_last
);
  wire  Queue_clock; // @[Decoupled.scala 287:21]
  wire  Queue_reset; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_read; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_enq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_extra; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_read; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_deq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_extra; // @[Decoupled.scala 287:21]
  reg [2:0] sels_0; // @[Mux.scala 32:23]
  reg [31:0] _RAND_0;
  reg [2:0] sels_1; // @[Mux.scala 32:23]
  reg [31:0] _RAND_1;
  wire  _T_3; // @[Mux.scala 45:28]
  wire  _GEN_7; // @[Mux.scala 45:41]
  wire  _GEN_8; // @[Mux.scala 45:41]
  wire  _T_4; // @[Mux.scala 45:28]
  wire  _GEN_12; // @[Mux.scala 45:41]
  wire [31:0] _GEN_15; // @[Mux.scala 45:41]
  wire  _GEN_16; // @[Mux.scala 45:41]
  wire  _GEN_17; // @[Mux.scala 45:41]
  wire  _T_5; // @[Mux.scala 45:28]
  wire  _GEN_21; // @[Mux.scala 45:41]
  wire [31:0] _GEN_24; // @[Mux.scala 45:41]
  wire  _GEN_25; // @[Mux.scala 45:41]
  wire  _GEN_26; // @[Mux.scala 45:41]
  wire  _T_6; // @[Mux.scala 45:28]
  wire  _GEN_30; // @[Mux.scala 45:41]
  wire [31:0] _GEN_33; // @[Mux.scala 45:41]
  wire  _GEN_34; // @[Mux.scala 45:41]
  wire  _T_7; // @[Mux.scala 45:28]
  wire  _T_8; // @[Mux.scala 40:46]
  wire [2:0] _T_10; // @[Mux.scala 41:29]
  wire  _T_11; // @[Mux.scala 45:28]
  wire  _T_12; // @[Mux.scala 45:28]
  wire  _T_13; // @[Mux.scala 45:28]
  wire  _T_17; // @[RegisterRouter.scala 40:39]
  wire  _T_18; // @[RegisterRouter.scala 40:26]
  wire  _T_19; // @[RegisterRouter.scala 42:29]
  wire  _T_62_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 290:17]
  wire [29:0] _T_26; // @[RegisterRouter.scala 48:19]
  wire [1:0] _T_66; // @[RegisterRouter.scala 59:16]
  wire  _T_68; // @[RegisterRouter.scala 59:16]
  wire  _T_20; // @[RegisterRouter.scala 42:26]
  wire [1:0] _T_29; // @[OneHot.scala 65:12]
  wire [1:0] _T_31; // @[Misc.scala 200:81]
  wire  _T_32; // @[Misc.scala 204:21]
  wire  _T_35; // @[Misc.scala 209:20]
  wire  _T_37; // @[Misc.scala 213:38]
  wire  _T_38; // @[Misc.scala 213:29]
  wire  _T_40; // @[Misc.scala 213:38]
  wire  _T_41; // @[Misc.scala 213:29]
  wire  _T_44; // @[Misc.scala 209:20]
  wire  _T_45; // @[Misc.scala 212:27]
  wire  _T_46; // @[Misc.scala 213:38]
  wire  _T_47; // @[Misc.scala 213:29]
  wire  _T_48; // @[Misc.scala 212:27]
  wire  _T_49; // @[Misc.scala 213:38]
  wire  _T_50; // @[Misc.scala 213:29]
  wire  _T_51; // @[Misc.scala 212:27]
  wire  _T_52; // @[Misc.scala 213:38]
  wire  _T_53; // @[Misc.scala 213:29]
  wire  _T_54; // @[Misc.scala 212:27]
  wire  _T_55; // @[Misc.scala 213:38]
  wire  _T_56; // @[Misc.scala 213:29]
  wire [3:0] _T_59; // @[Cat.scala 29:58]
  wire [3:0] _T_61; // @[RegisterRouter.scala 54:25]
  wire [7:0] _T_80; // @[Bitwise.scala 72:12]
  wire [7:0] _T_82; // @[Bitwise.scala 72:12]
  wire [7:0] _T_84; // @[Bitwise.scala 72:12]
  wire [7:0] _T_86; // @[Bitwise.scala 72:12]
  wire [31:0] _T_89; // @[Cat.scala 29:58]
  wire  _T_108; // @[RegisterRouter.scala 59:16]
  wire  _T_161; // @[RegisterRouter.scala 59:16]
  wire [1:0] _T_155; // @[OneHot.scala 58:35]
  wire  _T_178; // @[RegisterRouter.scala 59:16]
  wire  _T_185; // @[RegisterRouter.scala 59:16]
  wire  _T_186; // @[RegisterRouter.scala 59:16]
  wire  _T_115; // @[RegisterRouter.scala 59:16]
  wire  _T_180; // @[RegisterRouter.scala 59:16]
  wire  _T_181; // @[RegisterRouter.scala 59:16]
  wire  _T_138; // @[RegisterRouter.scala 59:16]
  wire  _GEN_101; // @[MuxLiteral.scala 48:10]
  wire [2:0] _GEN_103; // @[MuxLiteral.scala 48:10]
  wire [2:0] _T_235; // @[RegisterRouter.scala 59:16]
  wire  _T_236_bits_read; // @[Decoupled.scala 308:19 Decoupled.scala 309:14]
  wire  _T_236_valid; // @[Decoupled.scala 308:19 Decoupled.scala 310:15]
  wire  _T_239; // @[RegisterRouter.scala 65:29]
  Queue Queue ( // @[Decoupled.scala 287:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_read(Queue_io_enq_bits_read),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_extra(Queue_io_enq_bits_extra),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_read(Queue_io_deq_bits_read),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_extra(Queue_io_deq_bits_extra)
  );
  assign _T_3 = sels_0 == 3'h0; // @[Mux.scala 45:28]
  assign _GEN_7 = _T_3 & auto_stream_in_0_valid; // @[Mux.scala 45:41]
  assign _GEN_8 = _T_3 & auto_stream_out_0_ready; // @[Mux.scala 45:41]
  assign _T_4 = sels_0 == 3'h1; // @[Mux.scala 45:28]
  assign _GEN_12 = _T_4 ? auto_stream_in_1_bits_last : auto_stream_in_0_bits_last; // @[Mux.scala 45:41]
  assign _GEN_15 = _T_4 ? auto_stream_in_1_bits_data : auto_stream_in_0_bits_data; // @[Mux.scala 45:41]
  assign _GEN_16 = _T_4 ? auto_stream_in_1_valid : _GEN_7; // @[Mux.scala 45:41]
  assign _GEN_17 = _T_4 & auto_stream_out_0_ready; // @[Mux.scala 45:41]
  assign _T_5 = sels_0 == 3'h2; // @[Mux.scala 45:28]
  assign _GEN_21 = _T_5 ? auto_stream_in_2_bits_last : _GEN_12; // @[Mux.scala 45:41]
  assign _GEN_24 = _T_5 ? auto_stream_in_2_bits_data : _GEN_15; // @[Mux.scala 45:41]
  assign _GEN_25 = _T_5 ? auto_stream_in_2_valid : _GEN_16; // @[Mux.scala 45:41]
  assign _GEN_26 = _T_5 & auto_stream_out_0_ready; // @[Mux.scala 45:41]
  assign _T_6 = sels_0 == 3'h3; // @[Mux.scala 45:28]
  assign _GEN_30 = _T_6 ? 1'h0 : _GEN_21; // @[Mux.scala 45:41]
  assign _GEN_33 = _T_6 ? 32'hffffffff : _GEN_24; // @[Mux.scala 45:41]
  assign _GEN_34 = _T_6 | _GEN_25; // @[Mux.scala 45:41]
  assign _T_7 = sels_0 == 3'h4; // @[Mux.scala 45:28]
  assign _T_8 = sels_0 == sels_1; // @[Mux.scala 40:46]
  assign _T_10 = _T_8 ? 3'h5 : sels_1; // @[Mux.scala 41:29]
  assign _T_11 = _T_10 == 3'h0; // @[Mux.scala 45:28]
  assign _T_12 = _T_10 == 3'h1; // @[Mux.scala 45:28]
  assign _T_13 = _T_10 == 3'h2; // @[Mux.scala 45:28]
  assign _T_17 = auto_register_in_aw_valid & auto_register_in_w_valid; // @[RegisterRouter.scala 40:39]
  assign _T_18 = auto_register_in_ar_valid | _T_17; // @[RegisterRouter.scala 40:26]
  assign _T_19 = ~auto_register_in_ar_valid; // @[RegisterRouter.scala 42:29]
  assign _T_62_ready = Queue_io_enq_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 290:17]
  assign _T_26 = auto_register_in_ar_valid ? auto_register_in_ar_bits_addr : auto_register_in_aw_bits_addr; // @[RegisterRouter.scala 48:19]
  assign _T_66 = _T_26[3:2] & 2'h2; // @[RegisterRouter.scala 59:16]
  assign _T_68 = _T_66 == 2'h0; // @[RegisterRouter.scala 59:16]
  assign _T_20 = _T_62_ready & _T_19; // @[RegisterRouter.scala 42:26]
  assign _T_29 = 2'h1 << auto_register_in_ar_bits_size[0]; // @[OneHot.scala 65:12]
  assign _T_31 = _T_29 | 2'h1; // @[Misc.scala 200:81]
  assign _T_32 = auto_register_in_ar_bits_size >= 3'h2; // @[Misc.scala 204:21]
  assign _T_35 = ~auto_register_in_ar_bits_addr[1]; // @[Misc.scala 209:20]
  assign _T_37 = _T_31[1] & _T_35; // @[Misc.scala 213:38]
  assign _T_38 = _T_32 | _T_37; // @[Misc.scala 213:29]
  assign _T_40 = _T_31[1] & auto_register_in_ar_bits_addr[1]; // @[Misc.scala 213:38]
  assign _T_41 = _T_32 | _T_40; // @[Misc.scala 213:29]
  assign _T_44 = ~auto_register_in_ar_bits_addr[0]; // @[Misc.scala 209:20]
  assign _T_45 = _T_35 & _T_44; // @[Misc.scala 212:27]
  assign _T_46 = _T_31[0] & _T_45; // @[Misc.scala 213:38]
  assign _T_47 = _T_38 | _T_46; // @[Misc.scala 213:29]
  assign _T_48 = _T_35 & auto_register_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  assign _T_49 = _T_31[0] & _T_48; // @[Misc.scala 213:38]
  assign _T_50 = _T_38 | _T_49; // @[Misc.scala 213:29]
  assign _T_51 = auto_register_in_ar_bits_addr[1] & _T_44; // @[Misc.scala 212:27]
  assign _T_52 = _T_31[0] & _T_51; // @[Misc.scala 213:38]
  assign _T_53 = _T_41 | _T_52; // @[Misc.scala 213:29]
  assign _T_54 = auto_register_in_ar_bits_addr[1] & auto_register_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  assign _T_55 = _T_31[0] & _T_54; // @[Misc.scala 213:38]
  assign _T_56 = _T_41 | _T_55; // @[Misc.scala 213:29]
  assign _T_59 = {_T_56,_T_53,_T_50,_T_47}; // @[Cat.scala 29:58]
  assign _T_61 = auto_register_in_ar_valid ? _T_59 : auto_register_in_w_bits_strb; // @[RegisterRouter.scala 54:25]
  assign _T_80 = _T_61[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_82 = _T_61[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_84 = _T_61[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_86 = _T_61[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_89 = {_T_86,_T_84,_T_82,_T_80}; // @[Cat.scala 29:58]
  assign _T_108 = _T_89[2:0] == 3'h7; // @[RegisterRouter.scala 59:16]
  assign _T_161 = _T_18 & _T_62_ready; // @[RegisterRouter.scala 59:16]
  assign _T_155 = 2'h1 << _T_26[2]; // @[OneHot.scala 58:35]
  assign _T_178 = _T_161 & _T_19; // @[RegisterRouter.scala 59:16]
  assign _T_185 = _T_178 & _T_155[1]; // @[RegisterRouter.scala 59:16]
  assign _T_186 = _T_185 & _T_68; // @[RegisterRouter.scala 59:16]
  assign _T_115 = _T_186 & _T_108; // @[RegisterRouter.scala 59:16]
  assign _T_180 = _T_178 & _T_155[0]; // @[RegisterRouter.scala 59:16]
  assign _T_181 = _T_180 & _T_68; // @[RegisterRouter.scala 59:16]
  assign _T_138 = _T_181 & _T_108; // @[RegisterRouter.scala 59:16]
  assign _GEN_101 = _T_26[2] ? _T_68 : _T_68; // @[MuxLiteral.scala 48:10]
  assign _GEN_103 = _T_26[2] ? sels_1 : sels_0; // @[MuxLiteral.scala 48:10]
  assign _T_235 = _GEN_101 ? _GEN_103 : 3'h0; // @[RegisterRouter.scala 59:16]
  assign _T_236_bits_read = Queue_io_deq_bits_read; // @[Decoupled.scala 308:19 Decoupled.scala 309:14]
  assign _T_236_valid = Queue_io_deq_valid; // @[Decoupled.scala 308:19 Decoupled.scala 310:15]
  assign _T_239 = ~_T_236_bits_read; // @[RegisterRouter.scala 65:29]
  assign auto_register_in_aw_ready = _T_20 & auto_register_in_w_valid; // @[LazyModule.scala 173:31]
  assign auto_register_in_w_ready = _T_20 & auto_register_in_aw_valid; // @[LazyModule.scala 173:31]
  assign auto_register_in_b_valid = _T_236_valid & _T_239; // @[LazyModule.scala 173:31]
  assign auto_register_in_b_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_register_in_ar_ready = Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_register_in_r_valid = _T_236_valid & _T_236_bits_read; // @[LazyModule.scala 173:31]
  assign auto_register_in_r_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_register_in_r_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 173:31]
  assign auto_stream_in_2_ready = _T_13 | _GEN_26; // @[LazyModule.scala 173:31]
  assign auto_stream_in_1_ready = _T_12 | _GEN_17; // @[LazyModule.scala 173:31]
  assign auto_stream_in_0_ready = _T_11 | _GEN_8; // @[LazyModule.scala 173:31]
  assign auto_stream_out_0_valid = _T_7 | _GEN_34; // @[LazyModule.scala 173:49]
  assign auto_stream_out_0_bits_data = _T_7 ? 32'h0 : _GEN_33; // @[LazyModule.scala 173:49]
  assign auto_stream_out_0_bits_last = _T_7 ? 1'h0 : _GEN_30; // @[LazyModule.scala 173:49]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_register_in_ar_valid | _T_17; // @[Decoupled.scala 288:22]
  assign Queue_io_enq_bits_read = auto_register_in_ar_valid; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_data = {{29'd0}, _T_235}; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_extra = auto_register_in_ar_valid ? auto_register_in_ar_bits_id : auto_register_in_aw_bits_id; // @[Decoupled.scala 289:21]
  assign Queue_io_deq_ready = _T_236_bits_read ? auto_register_in_r_ready : auto_register_in_b_ready; // @[Decoupled.scala 311:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  sels_0 = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  sels_1 = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      sels_0 <= 3'h5;
    end else if (_T_138) begin
      sels_0 <= auto_register_in_w_bits_data[2:0];
    end
    if (reset) begin
      sels_1 <= 3'h5;
    end else if (_T_115) begin
      sels_1 <= auto_register_in_w_bits_data[2:0];
    end
  end
endmodule
module AXI4StreamMux_1(
  input         clock,
  input         reset,
  output        auto_register_in_aw_ready,
  input         auto_register_in_aw_valid,
  input         auto_register_in_aw_bits_id,
  input  [29:0] auto_register_in_aw_bits_addr,
  output        auto_register_in_w_ready,
  input         auto_register_in_w_valid,
  input  [31:0] auto_register_in_w_bits_data,
  input  [3:0]  auto_register_in_w_bits_strb,
  input         auto_register_in_b_ready,
  output        auto_register_in_b_valid,
  output        auto_register_in_b_bits_id,
  output        auto_register_in_ar_ready,
  input         auto_register_in_ar_valid,
  input         auto_register_in_ar_bits_id,
  input  [29:0] auto_register_in_ar_bits_addr,
  input  [2:0]  auto_register_in_ar_bits_size,
  input         auto_register_in_r_ready,
  output        auto_register_in_r_valid,
  output        auto_register_in_r_bits_id,
  output [31:0] auto_register_in_r_bits_data,
  output        auto_stream_in_ready,
  input         auto_stream_in_valid,
  input  [31:0] auto_stream_in_bits_data,
  input         auto_stream_in_bits_last,
  input         auto_stream_out_1_ready,
  output        auto_stream_out_1_valid,
  output [31:0] auto_stream_out_1_bits_data,
  output        auto_stream_out_1_bits_last
);
  wire  Queue_clock; // @[Decoupled.scala 287:21]
  wire  Queue_reset; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_read; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_enq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_extra; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_read; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_deq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_extra; // @[Decoupled.scala 287:21]
  reg  sels_0; // @[Mux.scala 32:23]
  reg [31:0] _RAND_0;
  reg  sels_1; // @[Mux.scala 32:23]
  reg [31:0] _RAND_1;
  wire  _T_3; // @[Mux.scala 45:28]
  wire  _T_4; // @[Mux.scala 40:46]
  wire  _T_6; // @[Mux.scala 41:29]
  wire  _T_7; // @[Mux.scala 45:28]
  wire  _T_9; // @[RegisterRouter.scala 40:39]
  wire  _T_10; // @[RegisterRouter.scala 40:26]
  wire  _T_11; // @[RegisterRouter.scala 42:29]
  wire  _T_54_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 290:17]
  wire [29:0] _T_18; // @[RegisterRouter.scala 48:19]
  wire [1:0] _T_58; // @[RegisterRouter.scala 59:16]
  wire  _T_60; // @[RegisterRouter.scala 59:16]
  wire  _T_12; // @[RegisterRouter.scala 42:26]
  wire [1:0] _T_21; // @[OneHot.scala 65:12]
  wire [1:0] _T_23; // @[Misc.scala 200:81]
  wire  _T_24; // @[Misc.scala 204:21]
  wire  _T_27; // @[Misc.scala 209:20]
  wire  _T_29; // @[Misc.scala 213:38]
  wire  _T_30; // @[Misc.scala 213:29]
  wire  _T_32; // @[Misc.scala 213:38]
  wire  _T_33; // @[Misc.scala 213:29]
  wire  _T_36; // @[Misc.scala 209:20]
  wire  _T_37; // @[Misc.scala 212:27]
  wire  _T_38; // @[Misc.scala 213:38]
  wire  _T_39; // @[Misc.scala 213:29]
  wire  _T_40; // @[Misc.scala 212:27]
  wire  _T_41; // @[Misc.scala 213:38]
  wire  _T_42; // @[Misc.scala 213:29]
  wire  _T_43; // @[Misc.scala 212:27]
  wire  _T_44; // @[Misc.scala 213:38]
  wire  _T_45; // @[Misc.scala 213:29]
  wire  _T_46; // @[Misc.scala 212:27]
  wire  _T_47; // @[Misc.scala 213:38]
  wire  _T_48; // @[Misc.scala 213:29]
  wire [3:0] _T_51; // @[Cat.scala 29:58]
  wire [3:0] _T_53; // @[RegisterRouter.scala 54:25]
  wire [7:0] _T_72; // @[Bitwise.scala 72:12]
  wire [7:0] _T_74; // @[Bitwise.scala 72:12]
  wire [7:0] _T_76; // @[Bitwise.scala 72:12]
  wire [7:0] _T_78; // @[Bitwise.scala 72:12]
  wire [31:0] _T_81; // @[Cat.scala 29:58]
  wire  _T_153; // @[RegisterRouter.scala 59:16]
  wire [1:0] _T_147; // @[OneHot.scala 58:35]
  wire  _T_170; // @[RegisterRouter.scala 59:16]
  wire  _T_177; // @[RegisterRouter.scala 59:16]
  wire  _T_178; // @[RegisterRouter.scala 59:16]
  wire  _T_107; // @[RegisterRouter.scala 59:16]
  wire  _GEN_18; // @[RegField.scala 134:88]
  wire  _T_172; // @[RegisterRouter.scala 59:16]
  wire  _T_173; // @[RegisterRouter.scala 59:16]
  wire  _T_130; // @[RegisterRouter.scala 59:16]
  wire  _GEN_19; // @[RegField.scala 134:88]
  wire  _GEN_29; // @[MuxLiteral.scala 48:10]
  wire  _GEN_31; // @[MuxLiteral.scala 48:10]
  wire  _T_227; // @[RegisterRouter.scala 59:16]
  wire  _T_228_bits_read; // @[Decoupled.scala 308:19 Decoupled.scala 309:14]
  wire  _T_228_valid; // @[Decoupled.scala 308:19 Decoupled.scala 310:15]
  wire  _T_231; // @[RegisterRouter.scala 65:29]
  Queue Queue ( // @[Decoupled.scala 287:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_read(Queue_io_enq_bits_read),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_extra(Queue_io_enq_bits_extra),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_read(Queue_io_deq_bits_read),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_extra(Queue_io_deq_bits_extra)
  );
  assign _T_3 = ~sels_0; // @[Mux.scala 45:28]
  assign _T_4 = sels_0 == sels_1; // @[Mux.scala 40:46]
  assign _T_6 = _T_4 | sels_1; // @[Mux.scala 41:29]
  assign _T_7 = ~_T_6; // @[Mux.scala 45:28]
  assign _T_9 = auto_register_in_aw_valid & auto_register_in_w_valid; // @[RegisterRouter.scala 40:39]
  assign _T_10 = auto_register_in_ar_valid | _T_9; // @[RegisterRouter.scala 40:26]
  assign _T_11 = ~auto_register_in_ar_valid; // @[RegisterRouter.scala 42:29]
  assign _T_54_ready = Queue_io_enq_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 290:17]
  assign _T_18 = auto_register_in_ar_valid ? auto_register_in_ar_bits_addr : auto_register_in_aw_bits_addr; // @[RegisterRouter.scala 48:19]
  assign _T_58 = _T_18[3:2] & 2'h2; // @[RegisterRouter.scala 59:16]
  assign _T_60 = _T_58 == 2'h0; // @[RegisterRouter.scala 59:16]
  assign _T_12 = _T_54_ready & _T_11; // @[RegisterRouter.scala 42:26]
  assign _T_21 = 2'h1 << auto_register_in_ar_bits_size[0]; // @[OneHot.scala 65:12]
  assign _T_23 = _T_21 | 2'h1; // @[Misc.scala 200:81]
  assign _T_24 = auto_register_in_ar_bits_size >= 3'h2; // @[Misc.scala 204:21]
  assign _T_27 = ~auto_register_in_ar_bits_addr[1]; // @[Misc.scala 209:20]
  assign _T_29 = _T_23[1] & _T_27; // @[Misc.scala 213:38]
  assign _T_30 = _T_24 | _T_29; // @[Misc.scala 213:29]
  assign _T_32 = _T_23[1] & auto_register_in_ar_bits_addr[1]; // @[Misc.scala 213:38]
  assign _T_33 = _T_24 | _T_32; // @[Misc.scala 213:29]
  assign _T_36 = ~auto_register_in_ar_bits_addr[0]; // @[Misc.scala 209:20]
  assign _T_37 = _T_27 & _T_36; // @[Misc.scala 212:27]
  assign _T_38 = _T_23[0] & _T_37; // @[Misc.scala 213:38]
  assign _T_39 = _T_30 | _T_38; // @[Misc.scala 213:29]
  assign _T_40 = _T_27 & auto_register_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  assign _T_41 = _T_23[0] & _T_40; // @[Misc.scala 213:38]
  assign _T_42 = _T_30 | _T_41; // @[Misc.scala 213:29]
  assign _T_43 = auto_register_in_ar_bits_addr[1] & _T_36; // @[Misc.scala 212:27]
  assign _T_44 = _T_23[0] & _T_43; // @[Misc.scala 213:38]
  assign _T_45 = _T_33 | _T_44; // @[Misc.scala 213:29]
  assign _T_46 = auto_register_in_ar_bits_addr[1] & auto_register_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  assign _T_47 = _T_23[0] & _T_46; // @[Misc.scala 213:38]
  assign _T_48 = _T_33 | _T_47; // @[Misc.scala 213:29]
  assign _T_51 = {_T_48,_T_45,_T_42,_T_39}; // @[Cat.scala 29:58]
  assign _T_53 = auto_register_in_ar_valid ? _T_51 : auto_register_in_w_bits_strb; // @[RegisterRouter.scala 54:25]
  assign _T_72 = _T_53[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_74 = _T_53[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_76 = _T_53[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_78 = _T_53[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_81 = {_T_78,_T_76,_T_74,_T_72}; // @[Cat.scala 29:58]
  assign _T_153 = _T_10 & _T_54_ready; // @[RegisterRouter.scala 59:16]
  assign _T_147 = 2'h1 << _T_18[2]; // @[OneHot.scala 58:35]
  assign _T_170 = _T_153 & _T_11; // @[RegisterRouter.scala 59:16]
  assign _T_177 = _T_170 & _T_147[1]; // @[RegisterRouter.scala 59:16]
  assign _T_178 = _T_177 & _T_60; // @[RegisterRouter.scala 59:16]
  assign _T_107 = _T_178 & _T_81[0]; // @[RegisterRouter.scala 59:16]
  assign _GEN_18 = _T_107 ? auto_register_in_w_bits_data[0] : sels_1; // @[RegField.scala 134:88]
  assign _T_172 = _T_170 & _T_147[0]; // @[RegisterRouter.scala 59:16]
  assign _T_173 = _T_172 & _T_60; // @[RegisterRouter.scala 59:16]
  assign _T_130 = _T_173 & _T_81[0]; // @[RegisterRouter.scala 59:16]
  assign _GEN_19 = _T_130 ? auto_register_in_w_bits_data[0] : sels_0; // @[RegField.scala 134:88]
  assign _GEN_29 = _T_18[2] ? _T_60 : _T_60; // @[MuxLiteral.scala 48:10]
  assign _GEN_31 = _T_18[2] ? sels_1 : sels_0; // @[MuxLiteral.scala 48:10]
  assign _T_227 = _GEN_29 & _GEN_31; // @[RegisterRouter.scala 59:16]
  assign _T_228_bits_read = Queue_io_deq_bits_read; // @[Decoupled.scala 308:19 Decoupled.scala 309:14]
  assign _T_228_valid = Queue_io_deq_valid; // @[Decoupled.scala 308:19 Decoupled.scala 310:15]
  assign _T_231 = ~_T_228_bits_read; // @[RegisterRouter.scala 65:29]
  assign auto_register_in_aw_ready = _T_12 & auto_register_in_w_valid; // @[LazyModule.scala 173:31]
  assign auto_register_in_w_ready = _T_12 & auto_register_in_aw_valid; // @[LazyModule.scala 173:31]
  assign auto_register_in_b_valid = _T_228_valid & _T_231; // @[LazyModule.scala 173:31]
  assign auto_register_in_b_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_register_in_ar_ready = Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_register_in_r_valid = _T_228_valid & _T_228_bits_read; // @[LazyModule.scala 173:31]
  assign auto_register_in_r_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_register_in_r_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 173:31]
  assign auto_stream_in_ready = _T_7 ? auto_stream_out_1_ready : _T_3; // @[LazyModule.scala 173:31]
  assign auto_stream_out_1_valid = _T_7 & auto_stream_in_valid; // @[LazyModule.scala 173:49]
  assign auto_stream_out_1_bits_data = auto_stream_in_bits_data; // @[LazyModule.scala 173:49]
  assign auto_stream_out_1_bits_last = auto_stream_in_bits_last; // @[LazyModule.scala 173:49]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_register_in_ar_valid | _T_9; // @[Decoupled.scala 288:22]
  assign Queue_io_enq_bits_read = auto_register_in_ar_valid; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_data = {{31'd0}, _T_227}; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_extra = auto_register_in_ar_valid ? auto_register_in_ar_bits_id : auto_register_in_aw_bits_id; // @[Decoupled.scala 289:21]
  assign Queue_io_deq_ready = _T_228_bits_read ? auto_register_in_r_ready : auto_register_in_b_ready; // @[Decoupled.scala 311:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  sels_0 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  sels_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    sels_0 <= reset | _GEN_19;
    sels_1 <= reset | _GEN_18;
  end
endmodule
module NCOTableStandardMode(
  input  [8:0]  io_phase,
  output [15:0] io_sinOut,
  output [15:0] io_cosOut
);
  wire [1:0] msbs; // @[NCOTable.scala 123:15]
  wire [6:0] addr; // @[NCOTable.scala 131:15]
  wire  _T_24; // @[Conditional.scala 37:30]
  wire [6:0] _T_26; // @[NCOTable.scala 173:9]
  wire  _T_33; // @[Conditional.scala 37:30]
  wire  _T_42; // @[Conditional.scala 37:30]
  wire  _T_51; // @[Conditional.scala 37:30]
  wire [6:0] _GEN_1; // @[Conditional.scala 39:67]
  wire [6:0] _GEN_7; // @[Conditional.scala 39:67]
  wire [6:0] _GEN_15; // @[Conditional.scala 39:67]
  wire [6:0] cosAddr; // @[Conditional.scala 40:58]
  wire  _T_27; // @[NCOTable.scala 199:27]
  wire  _T_28; // @[NCOTable.scala 199:43]
  wire  _T_29; // @[NCOTable.scala 199:35]
  wire [6:0] _GEN_0; // @[Conditional.scala 39:67]
  wire [6:0] _GEN_6; // @[Conditional.scala 39:67]
  wire [6:0] _GEN_14; // @[Conditional.scala 39:67]
  wire [6:0] sinAddr; // @[Conditional.scala 40:58]
  wire  _T_36; // @[NCOTable.scala 209:27]
  wire  _T_38; // @[NCOTable.scala 209:35]
  wire  _GEN_4; // @[Conditional.scala 39:67]
  wire  _GEN_8; // @[Conditional.scala 39:67]
  wire  _GEN_10; // @[Conditional.scala 39:67]
  wire  _GEN_12; // @[Conditional.scala 39:67]
  wire  _GEN_16; // @[Conditional.scala 39:67]
  wire  _GEN_17; // @[Conditional.scala 39:67]
  wire  _GEN_18; // @[Conditional.scala 39:67]
  wire  _GEN_20; // @[Conditional.scala 39:67]
  wire  sinNegative2; // @[Conditional.scala 40:58]
  wire  cosNegative2; // @[Conditional.scala 40:58]
  wire  _GEN_26; // @[Conditional.scala 40:58]
  wire  _GEN_28; // @[Conditional.scala 40:58]
  wire [15:0] _GEN_31; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_32; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_33; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_34; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_35; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_36; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_37; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_38; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_39; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_40; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_41; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_42; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_43; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_44; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_45; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_46; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_47; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_48; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_49; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_50; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_51; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_52; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_53; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_54; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_55; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_56; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_57; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_58; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_59; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_60; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_61; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_62; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_63; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_64; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_65; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_66; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_67; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_68; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_69; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_70; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_71; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_72; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_73; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_74; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_75; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_76; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_77; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_78; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_79; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_80; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_81; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_82; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_83; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_84; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_85; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_86; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_87; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_88; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_89; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_90; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_91; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_92; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_93; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_94; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_95; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_96; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_97; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_98; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_99; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_100; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_101; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_102; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_103; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_104; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_105; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_106; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_107; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_108; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_109; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_110; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_111; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_112; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_113; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_114; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_115; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_116; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_117; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_118; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_119; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_120; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_121; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_122; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_123; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_124; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_125; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_126; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_127; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_128; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_129; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_130; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_131; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_132; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_133; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_134; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_135; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_136; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_137; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_138; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_139; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_140; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_141; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_142; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_143; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_144; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_145; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_146; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_147; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_148; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_149; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_150; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_151; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_152; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_153; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_154; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_155; // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_156; // @[NCOTable.scala 260:64]
  wire [15:0] _T_65; // @[NCOTable.scala 260:64]
  wire [15:0] sinTableOut; // @[NCOTable.scala 260:23]
  wire [15:0] _GEN_159; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_160; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_161; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_162; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_163; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_164; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_165; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_166; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_167; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_168; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_169; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_170; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_171; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_172; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_173; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_174; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_175; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_176; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_177; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_178; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_179; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_180; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_181; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_182; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_183; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_184; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_185; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_186; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_187; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_188; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_189; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_190; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_191; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_192; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_193; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_194; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_195; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_196; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_197; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_198; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_199; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_200; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_201; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_202; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_203; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_204; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_205; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_206; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_207; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_208; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_209; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_210; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_211; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_212; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_213; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_214; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_215; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_216; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_217; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_218; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_219; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_220; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_221; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_222; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_223; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_224; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_225; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_226; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_227; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_228; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_229; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_230; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_231; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_232; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_233; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_234; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_235; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_236; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_237; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_238; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_239; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_240; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_241; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_242; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_243; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_244; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_245; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_246; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_247; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_248; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_249; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_250; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_251; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_252; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_253; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_254; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_255; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_256; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_257; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_258; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_259; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_260; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_261; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_262; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_263; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_264; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_265; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_266; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_267; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_268; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_269; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_270; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_271; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_272; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_273; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_274; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_275; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_276; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_277; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_278; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_279; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_280; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_281; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_282; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_283; // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_284; // @[NCOTable.scala 261:64]
  wire [15:0] _T_71; // @[NCOTable.scala 261:64]
  wire [15:0] cosTableOut; // @[NCOTable.scala 261:23]
  wire [15:0] _T_75; // @[FixedPointTypeClass.scala 39:43]
  wire [15:0] _T_78; // @[FixedPointTypeClass.scala 39:43]
  assign msbs = io_phase[8:7]; // @[NCOTable.scala 123:15]
  assign addr = io_phase[6:0]; // @[NCOTable.scala 131:15]
  assign _T_24 = 2'h0 == msbs; // @[Conditional.scala 37:30]
  assign _T_26 = 7'h0 - addr; // @[NCOTable.scala 173:9]
  assign _T_33 = 2'h1 == msbs; // @[Conditional.scala 37:30]
  assign _T_42 = 2'h2 == msbs; // @[Conditional.scala 37:30]
  assign _T_51 = 2'h3 == msbs; // @[Conditional.scala 37:30]
  assign _GEN_1 = _T_51 ? addr : 7'h0; // @[Conditional.scala 39:67]
  assign _GEN_7 = _T_42 ? _T_26 : _GEN_1; // @[Conditional.scala 39:67]
  assign _GEN_15 = _T_33 ? addr : _GEN_7; // @[Conditional.scala 39:67]
  assign cosAddr = _T_24 ? _T_26 : _GEN_15; // @[Conditional.scala 40:58]
  assign _T_27 = cosAddr == 7'h0; // @[NCOTable.scala 199:27]
  assign _T_28 = addr == 7'h0; // @[NCOTable.scala 199:43]
  assign _T_29 = _T_27 & _T_28; // @[NCOTable.scala 199:35]
  assign _GEN_0 = _T_51 ? _T_26 : 7'h0; // @[Conditional.scala 39:67]
  assign _GEN_6 = _T_42 ? addr : _GEN_0; // @[Conditional.scala 39:67]
  assign _GEN_14 = _T_33 ? _T_26 : _GEN_6; // @[Conditional.scala 39:67]
  assign sinAddr = _T_24 ? addr : _GEN_14; // @[Conditional.scala 40:58]
  assign _T_36 = sinAddr == 7'h0; // @[NCOTable.scala 209:27]
  assign _T_38 = _T_36 & _T_28; // @[NCOTable.scala 209:35]
  assign _GEN_4 = _T_51 & _T_38; // @[Conditional.scala 39:67]
  assign _GEN_8 = _T_42 | _T_51; // @[Conditional.scala 39:67]
  assign _GEN_10 = _T_42 & _T_29; // @[Conditional.scala 39:67]
  assign _GEN_12 = _T_42 ? 1'h0 : _GEN_4; // @[Conditional.scala 39:67]
  assign _GEN_16 = _T_33 ? 1'h0 : _GEN_8; // @[Conditional.scala 39:67]
  assign _GEN_17 = _T_33 | _T_42; // @[Conditional.scala 39:67]
  assign _GEN_18 = _T_33 ? _T_38 : _GEN_12; // @[Conditional.scala 39:67]
  assign _GEN_20 = _T_33 ? 1'h0 : _GEN_10; // @[Conditional.scala 39:67]
  assign sinNegative2 = _T_24 ? 1'h0 : _GEN_16; // @[Conditional.scala 40:58]
  assign cosNegative2 = _T_24 ? 1'h0 : _GEN_17; // @[Conditional.scala 40:58]
  assign _GEN_26 = _T_24 ? _T_29 : _GEN_20; // @[Conditional.scala 40:58]
  assign _GEN_28 = _T_24 ? 1'h0 : _GEN_18; // @[Conditional.scala 40:58]
  assign _GEN_31 = 7'h1 == sinAddr ? $signed(16'shc9) : $signed(16'sh0); // @[NCOTable.scala 260:64]
  assign _GEN_32 = 7'h2 == sinAddr ? $signed(16'sh192) : $signed(_GEN_31); // @[NCOTable.scala 260:64]
  assign _GEN_33 = 7'h3 == sinAddr ? $signed(16'sh25b) : $signed(_GEN_32); // @[NCOTable.scala 260:64]
  assign _GEN_34 = 7'h4 == sinAddr ? $signed(16'sh324) : $signed(_GEN_33); // @[NCOTable.scala 260:64]
  assign _GEN_35 = 7'h5 == sinAddr ? $signed(16'sh3ed) : $signed(_GEN_34); // @[NCOTable.scala 260:64]
  assign _GEN_36 = 7'h6 == sinAddr ? $signed(16'sh4b5) : $signed(_GEN_35); // @[NCOTable.scala 260:64]
  assign _GEN_37 = 7'h7 == sinAddr ? $signed(16'sh57e) : $signed(_GEN_36); // @[NCOTable.scala 260:64]
  assign _GEN_38 = 7'h8 == sinAddr ? $signed(16'sh646) : $signed(_GEN_37); // @[NCOTable.scala 260:64]
  assign _GEN_39 = 7'h9 == sinAddr ? $signed(16'sh70e) : $signed(_GEN_38); // @[NCOTable.scala 260:64]
  assign _GEN_40 = 7'ha == sinAddr ? $signed(16'sh7d6) : $signed(_GEN_39); // @[NCOTable.scala 260:64]
  assign _GEN_41 = 7'hb == sinAddr ? $signed(16'sh89d) : $signed(_GEN_40); // @[NCOTable.scala 260:64]
  assign _GEN_42 = 7'hc == sinAddr ? $signed(16'sh964) : $signed(_GEN_41); // @[NCOTable.scala 260:64]
  assign _GEN_43 = 7'hd == sinAddr ? $signed(16'sha2b) : $signed(_GEN_42); // @[NCOTable.scala 260:64]
  assign _GEN_44 = 7'he == sinAddr ? $signed(16'shaf1) : $signed(_GEN_43); // @[NCOTable.scala 260:64]
  assign _GEN_45 = 7'hf == sinAddr ? $signed(16'shbb7) : $signed(_GEN_44); // @[NCOTable.scala 260:64]
  assign _GEN_46 = 7'h10 == sinAddr ? $signed(16'shc7c) : $signed(_GEN_45); // @[NCOTable.scala 260:64]
  assign _GEN_47 = 7'h11 == sinAddr ? $signed(16'shd41) : $signed(_GEN_46); // @[NCOTable.scala 260:64]
  assign _GEN_48 = 7'h12 == sinAddr ? $signed(16'she06) : $signed(_GEN_47); // @[NCOTable.scala 260:64]
  assign _GEN_49 = 7'h13 == sinAddr ? $signed(16'sheca) : $signed(_GEN_48); // @[NCOTable.scala 260:64]
  assign _GEN_50 = 7'h14 == sinAddr ? $signed(16'shf8d) : $signed(_GEN_49); // @[NCOTable.scala 260:64]
  assign _GEN_51 = 7'h15 == sinAddr ? $signed(16'sh1050) : $signed(_GEN_50); // @[NCOTable.scala 260:64]
  assign _GEN_52 = 7'h16 == sinAddr ? $signed(16'sh1112) : $signed(_GEN_51); // @[NCOTable.scala 260:64]
  assign _GEN_53 = 7'h17 == sinAddr ? $signed(16'sh11d3) : $signed(_GEN_52); // @[NCOTable.scala 260:64]
  assign _GEN_54 = 7'h18 == sinAddr ? $signed(16'sh1294) : $signed(_GEN_53); // @[NCOTable.scala 260:64]
  assign _GEN_55 = 7'h19 == sinAddr ? $signed(16'sh1354) : $signed(_GEN_54); // @[NCOTable.scala 260:64]
  assign _GEN_56 = 7'h1a == sinAddr ? $signed(16'sh1413) : $signed(_GEN_55); // @[NCOTable.scala 260:64]
  assign _GEN_57 = 7'h1b == sinAddr ? $signed(16'sh14d2) : $signed(_GEN_56); // @[NCOTable.scala 260:64]
  assign _GEN_58 = 7'h1c == sinAddr ? $signed(16'sh1590) : $signed(_GEN_57); // @[NCOTable.scala 260:64]
  assign _GEN_59 = 7'h1d == sinAddr ? $signed(16'sh164c) : $signed(_GEN_58); // @[NCOTable.scala 260:64]
  assign _GEN_60 = 7'h1e == sinAddr ? $signed(16'sh1709) : $signed(_GEN_59); // @[NCOTable.scala 260:64]
  assign _GEN_61 = 7'h1f == sinAddr ? $signed(16'sh17c4) : $signed(_GEN_60); // @[NCOTable.scala 260:64]
  assign _GEN_62 = 7'h20 == sinAddr ? $signed(16'sh187e) : $signed(_GEN_61); // @[NCOTable.scala 260:64]
  assign _GEN_63 = 7'h21 == sinAddr ? $signed(16'sh1937) : $signed(_GEN_62); // @[NCOTable.scala 260:64]
  assign _GEN_64 = 7'h22 == sinAddr ? $signed(16'sh19ef) : $signed(_GEN_63); // @[NCOTable.scala 260:64]
  assign _GEN_65 = 7'h23 == sinAddr ? $signed(16'sh1aa7) : $signed(_GEN_64); // @[NCOTable.scala 260:64]
  assign _GEN_66 = 7'h24 == sinAddr ? $signed(16'sh1b5d) : $signed(_GEN_65); // @[NCOTable.scala 260:64]
  assign _GEN_67 = 7'h25 == sinAddr ? $signed(16'sh1c12) : $signed(_GEN_66); // @[NCOTable.scala 260:64]
  assign _GEN_68 = 7'h26 == sinAddr ? $signed(16'sh1cc6) : $signed(_GEN_67); // @[NCOTable.scala 260:64]
  assign _GEN_69 = 7'h27 == sinAddr ? $signed(16'sh1d79) : $signed(_GEN_68); // @[NCOTable.scala 260:64]
  assign _GEN_70 = 7'h28 == sinAddr ? $signed(16'sh1e2b) : $signed(_GEN_69); // @[NCOTable.scala 260:64]
  assign _GEN_71 = 7'h29 == sinAddr ? $signed(16'sh1edc) : $signed(_GEN_70); // @[NCOTable.scala 260:64]
  assign _GEN_72 = 7'h2a == sinAddr ? $signed(16'sh1f8c) : $signed(_GEN_71); // @[NCOTable.scala 260:64]
  assign _GEN_73 = 7'h2b == sinAddr ? $signed(16'sh203a) : $signed(_GEN_72); // @[NCOTable.scala 260:64]
  assign _GEN_74 = 7'h2c == sinAddr ? $signed(16'sh20e7) : $signed(_GEN_73); // @[NCOTable.scala 260:64]
  assign _GEN_75 = 7'h2d == sinAddr ? $signed(16'sh2193) : $signed(_GEN_74); // @[NCOTable.scala 260:64]
  assign _GEN_76 = 7'h2e == sinAddr ? $signed(16'sh223d) : $signed(_GEN_75); // @[NCOTable.scala 260:64]
  assign _GEN_77 = 7'h2f == sinAddr ? $signed(16'sh22e7) : $signed(_GEN_76); // @[NCOTable.scala 260:64]
  assign _GEN_78 = 7'h30 == sinAddr ? $signed(16'sh238e) : $signed(_GEN_77); // @[NCOTable.scala 260:64]
  assign _GEN_79 = 7'h31 == sinAddr ? $signed(16'sh2435) : $signed(_GEN_78); // @[NCOTable.scala 260:64]
  assign _GEN_80 = 7'h32 == sinAddr ? $signed(16'sh24da) : $signed(_GEN_79); // @[NCOTable.scala 260:64]
  assign _GEN_81 = 7'h33 == sinAddr ? $signed(16'sh257e) : $signed(_GEN_80); // @[NCOTable.scala 260:64]
  assign _GEN_82 = 7'h34 == sinAddr ? $signed(16'sh2620) : $signed(_GEN_81); // @[NCOTable.scala 260:64]
  assign _GEN_83 = 7'h35 == sinAddr ? $signed(16'sh26c1) : $signed(_GEN_82); // @[NCOTable.scala 260:64]
  assign _GEN_84 = 7'h36 == sinAddr ? $signed(16'sh2760) : $signed(_GEN_83); // @[NCOTable.scala 260:64]
  assign _GEN_85 = 7'h37 == sinAddr ? $signed(16'sh27fe) : $signed(_GEN_84); // @[NCOTable.scala 260:64]
  assign _GEN_86 = 7'h38 == sinAddr ? $signed(16'sh289a) : $signed(_GEN_85); // @[NCOTable.scala 260:64]
  assign _GEN_87 = 7'h39 == sinAddr ? $signed(16'sh2935) : $signed(_GEN_86); // @[NCOTable.scala 260:64]
  assign _GEN_88 = 7'h3a == sinAddr ? $signed(16'sh29ce) : $signed(_GEN_87); // @[NCOTable.scala 260:64]
  assign _GEN_89 = 7'h3b == sinAddr ? $signed(16'sh2a65) : $signed(_GEN_88); // @[NCOTable.scala 260:64]
  assign _GEN_90 = 7'h3c == sinAddr ? $signed(16'sh2afb) : $signed(_GEN_89); // @[NCOTable.scala 260:64]
  assign _GEN_91 = 7'h3d == sinAddr ? $signed(16'sh2b8f) : $signed(_GEN_90); // @[NCOTable.scala 260:64]
  assign _GEN_92 = 7'h3e == sinAddr ? $signed(16'sh2c21) : $signed(_GEN_91); // @[NCOTable.scala 260:64]
  assign _GEN_93 = 7'h3f == sinAddr ? $signed(16'sh2cb2) : $signed(_GEN_92); // @[NCOTable.scala 260:64]
  assign _GEN_94 = 7'h40 == sinAddr ? $signed(16'sh2d41) : $signed(_GEN_93); // @[NCOTable.scala 260:64]
  assign _GEN_95 = 7'h41 == sinAddr ? $signed(16'sh2dcf) : $signed(_GEN_94); // @[NCOTable.scala 260:64]
  assign _GEN_96 = 7'h42 == sinAddr ? $signed(16'sh2e5a) : $signed(_GEN_95); // @[NCOTable.scala 260:64]
  assign _GEN_97 = 7'h43 == sinAddr ? $signed(16'sh2ee4) : $signed(_GEN_96); // @[NCOTable.scala 260:64]
  assign _GEN_98 = 7'h44 == sinAddr ? $signed(16'sh2f6c) : $signed(_GEN_97); // @[NCOTable.scala 260:64]
  assign _GEN_99 = 7'h45 == sinAddr ? $signed(16'sh2ff2) : $signed(_GEN_98); // @[NCOTable.scala 260:64]
  assign _GEN_100 = 7'h46 == sinAddr ? $signed(16'sh3076) : $signed(_GEN_99); // @[NCOTable.scala 260:64]
  assign _GEN_101 = 7'h47 == sinAddr ? $signed(16'sh30f9) : $signed(_GEN_100); // @[NCOTable.scala 260:64]
  assign _GEN_102 = 7'h48 == sinAddr ? $signed(16'sh3179) : $signed(_GEN_101); // @[NCOTable.scala 260:64]
  assign _GEN_103 = 7'h49 == sinAddr ? $signed(16'sh31f8) : $signed(_GEN_102); // @[NCOTable.scala 260:64]
  assign _GEN_104 = 7'h4a == sinAddr ? $signed(16'sh3274) : $signed(_GEN_103); // @[NCOTable.scala 260:64]
  assign _GEN_105 = 7'h4b == sinAddr ? $signed(16'sh32ef) : $signed(_GEN_104); // @[NCOTable.scala 260:64]
  assign _GEN_106 = 7'h4c == sinAddr ? $signed(16'sh3368) : $signed(_GEN_105); // @[NCOTable.scala 260:64]
  assign _GEN_107 = 7'h4d == sinAddr ? $signed(16'sh33df) : $signed(_GEN_106); // @[NCOTable.scala 260:64]
  assign _GEN_108 = 7'h4e == sinAddr ? $signed(16'sh3453) : $signed(_GEN_107); // @[NCOTable.scala 260:64]
  assign _GEN_109 = 7'h4f == sinAddr ? $signed(16'sh34c6) : $signed(_GEN_108); // @[NCOTable.scala 260:64]
  assign _GEN_110 = 7'h50 == sinAddr ? $signed(16'sh3537) : $signed(_GEN_109); // @[NCOTable.scala 260:64]
  assign _GEN_111 = 7'h51 == sinAddr ? $signed(16'sh35a5) : $signed(_GEN_110); // @[NCOTable.scala 260:64]
  assign _GEN_112 = 7'h52 == sinAddr ? $signed(16'sh3612) : $signed(_GEN_111); // @[NCOTable.scala 260:64]
  assign _GEN_113 = 7'h53 == sinAddr ? $signed(16'sh367d) : $signed(_GEN_112); // @[NCOTable.scala 260:64]
  assign _GEN_114 = 7'h54 == sinAddr ? $signed(16'sh36e5) : $signed(_GEN_113); // @[NCOTable.scala 260:64]
  assign _GEN_115 = 7'h55 == sinAddr ? $signed(16'sh374b) : $signed(_GEN_114); // @[NCOTable.scala 260:64]
  assign _GEN_116 = 7'h56 == sinAddr ? $signed(16'sh37b0) : $signed(_GEN_115); // @[NCOTable.scala 260:64]
  assign _GEN_117 = 7'h57 == sinAddr ? $signed(16'sh3812) : $signed(_GEN_116); // @[NCOTable.scala 260:64]
  assign _GEN_118 = 7'h58 == sinAddr ? $signed(16'sh3871) : $signed(_GEN_117); // @[NCOTable.scala 260:64]
  assign _GEN_119 = 7'h59 == sinAddr ? $signed(16'sh38cf) : $signed(_GEN_118); // @[NCOTable.scala 260:64]
  assign _GEN_120 = 7'h5a == sinAddr ? $signed(16'sh392b) : $signed(_GEN_119); // @[NCOTable.scala 260:64]
  assign _GEN_121 = 7'h5b == sinAddr ? $signed(16'sh3984) : $signed(_GEN_120); // @[NCOTable.scala 260:64]
  assign _GEN_122 = 7'h5c == sinAddr ? $signed(16'sh39db) : $signed(_GEN_121); // @[NCOTable.scala 260:64]
  assign _GEN_123 = 7'h5d == sinAddr ? $signed(16'sh3a30) : $signed(_GEN_122); // @[NCOTable.scala 260:64]
  assign _GEN_124 = 7'h5e == sinAddr ? $signed(16'sh3a82) : $signed(_GEN_123); // @[NCOTable.scala 260:64]
  assign _GEN_125 = 7'h5f == sinAddr ? $signed(16'sh3ad3) : $signed(_GEN_124); // @[NCOTable.scala 260:64]
  assign _GEN_126 = 7'h60 == sinAddr ? $signed(16'sh3b21) : $signed(_GEN_125); // @[NCOTable.scala 260:64]
  assign _GEN_127 = 7'h61 == sinAddr ? $signed(16'sh3b6d) : $signed(_GEN_126); // @[NCOTable.scala 260:64]
  assign _GEN_128 = 7'h62 == sinAddr ? $signed(16'sh3bb6) : $signed(_GEN_127); // @[NCOTable.scala 260:64]
  assign _GEN_129 = 7'h63 == sinAddr ? $signed(16'sh3bfd) : $signed(_GEN_128); // @[NCOTable.scala 260:64]
  assign _GEN_130 = 7'h64 == sinAddr ? $signed(16'sh3c42) : $signed(_GEN_129); // @[NCOTable.scala 260:64]
  assign _GEN_131 = 7'h65 == sinAddr ? $signed(16'sh3c85) : $signed(_GEN_130); // @[NCOTable.scala 260:64]
  assign _GEN_132 = 7'h66 == sinAddr ? $signed(16'sh3cc5) : $signed(_GEN_131); // @[NCOTable.scala 260:64]
  assign _GEN_133 = 7'h67 == sinAddr ? $signed(16'sh3d03) : $signed(_GEN_132); // @[NCOTable.scala 260:64]
  assign _GEN_134 = 7'h68 == sinAddr ? $signed(16'sh3d3f) : $signed(_GEN_133); // @[NCOTable.scala 260:64]
  assign _GEN_135 = 7'h69 == sinAddr ? $signed(16'sh3d78) : $signed(_GEN_134); // @[NCOTable.scala 260:64]
  assign _GEN_136 = 7'h6a == sinAddr ? $signed(16'sh3daf) : $signed(_GEN_135); // @[NCOTable.scala 260:64]
  assign _GEN_137 = 7'h6b == sinAddr ? $signed(16'sh3de3) : $signed(_GEN_136); // @[NCOTable.scala 260:64]
  assign _GEN_138 = 7'h6c == sinAddr ? $signed(16'sh3e15) : $signed(_GEN_137); // @[NCOTable.scala 260:64]
  assign _GEN_139 = 7'h6d == sinAddr ? $signed(16'sh3e45) : $signed(_GEN_138); // @[NCOTable.scala 260:64]
  assign _GEN_140 = 7'h6e == sinAddr ? $signed(16'sh3e72) : $signed(_GEN_139); // @[NCOTable.scala 260:64]
  assign _GEN_141 = 7'h6f == sinAddr ? $signed(16'sh3e9d) : $signed(_GEN_140); // @[NCOTable.scala 260:64]
  assign _GEN_142 = 7'h70 == sinAddr ? $signed(16'sh3ec5) : $signed(_GEN_141); // @[NCOTable.scala 260:64]
  assign _GEN_143 = 7'h71 == sinAddr ? $signed(16'sh3eeb) : $signed(_GEN_142); // @[NCOTable.scala 260:64]
  assign _GEN_144 = 7'h72 == sinAddr ? $signed(16'sh3f0f) : $signed(_GEN_143); // @[NCOTable.scala 260:64]
  assign _GEN_145 = 7'h73 == sinAddr ? $signed(16'sh3f30) : $signed(_GEN_144); // @[NCOTable.scala 260:64]
  assign _GEN_146 = 7'h74 == sinAddr ? $signed(16'sh3f4f) : $signed(_GEN_145); // @[NCOTable.scala 260:64]
  assign _GEN_147 = 7'h75 == sinAddr ? $signed(16'sh3f6b) : $signed(_GEN_146); // @[NCOTable.scala 260:64]
  assign _GEN_148 = 7'h76 == sinAddr ? $signed(16'sh3f85) : $signed(_GEN_147); // @[NCOTable.scala 260:64]
  assign _GEN_149 = 7'h77 == sinAddr ? $signed(16'sh3f9c) : $signed(_GEN_148); // @[NCOTable.scala 260:64]
  assign _GEN_150 = 7'h78 == sinAddr ? $signed(16'sh3fb1) : $signed(_GEN_149); // @[NCOTable.scala 260:64]
  assign _GEN_151 = 7'h79 == sinAddr ? $signed(16'sh3fc4) : $signed(_GEN_150); // @[NCOTable.scala 260:64]
  assign _GEN_152 = 7'h7a == sinAddr ? $signed(16'sh3fd4) : $signed(_GEN_151); // @[NCOTable.scala 260:64]
  assign _GEN_153 = 7'h7b == sinAddr ? $signed(16'sh3fe1) : $signed(_GEN_152); // @[NCOTable.scala 260:64]
  assign _GEN_154 = 7'h7c == sinAddr ? $signed(16'sh3fec) : $signed(_GEN_153); // @[NCOTable.scala 260:64]
  assign _GEN_155 = 7'h7d == sinAddr ? $signed(16'sh3ff5) : $signed(_GEN_154); // @[NCOTable.scala 260:64]
  assign _GEN_156 = 7'h7e == sinAddr ? $signed(16'sh3ffb) : $signed(_GEN_155); // @[NCOTable.scala 260:64]
  assign _T_65 = 7'h7f == sinAddr ? $signed(16'sh3fff) : $signed(_GEN_156); // @[NCOTable.scala 260:64]
  assign sinTableOut = _GEN_28 ? $signed(16'sh4000) : $signed(_T_65); // @[NCOTable.scala 260:23]
  assign _GEN_159 = 7'h1 == cosAddr ? $signed(16'shc9) : $signed(16'sh0); // @[NCOTable.scala 261:64]
  assign _GEN_160 = 7'h2 == cosAddr ? $signed(16'sh192) : $signed(_GEN_159); // @[NCOTable.scala 261:64]
  assign _GEN_161 = 7'h3 == cosAddr ? $signed(16'sh25b) : $signed(_GEN_160); // @[NCOTable.scala 261:64]
  assign _GEN_162 = 7'h4 == cosAddr ? $signed(16'sh324) : $signed(_GEN_161); // @[NCOTable.scala 261:64]
  assign _GEN_163 = 7'h5 == cosAddr ? $signed(16'sh3ed) : $signed(_GEN_162); // @[NCOTable.scala 261:64]
  assign _GEN_164 = 7'h6 == cosAddr ? $signed(16'sh4b5) : $signed(_GEN_163); // @[NCOTable.scala 261:64]
  assign _GEN_165 = 7'h7 == cosAddr ? $signed(16'sh57e) : $signed(_GEN_164); // @[NCOTable.scala 261:64]
  assign _GEN_166 = 7'h8 == cosAddr ? $signed(16'sh646) : $signed(_GEN_165); // @[NCOTable.scala 261:64]
  assign _GEN_167 = 7'h9 == cosAddr ? $signed(16'sh70e) : $signed(_GEN_166); // @[NCOTable.scala 261:64]
  assign _GEN_168 = 7'ha == cosAddr ? $signed(16'sh7d6) : $signed(_GEN_167); // @[NCOTable.scala 261:64]
  assign _GEN_169 = 7'hb == cosAddr ? $signed(16'sh89d) : $signed(_GEN_168); // @[NCOTable.scala 261:64]
  assign _GEN_170 = 7'hc == cosAddr ? $signed(16'sh964) : $signed(_GEN_169); // @[NCOTable.scala 261:64]
  assign _GEN_171 = 7'hd == cosAddr ? $signed(16'sha2b) : $signed(_GEN_170); // @[NCOTable.scala 261:64]
  assign _GEN_172 = 7'he == cosAddr ? $signed(16'shaf1) : $signed(_GEN_171); // @[NCOTable.scala 261:64]
  assign _GEN_173 = 7'hf == cosAddr ? $signed(16'shbb7) : $signed(_GEN_172); // @[NCOTable.scala 261:64]
  assign _GEN_174 = 7'h10 == cosAddr ? $signed(16'shc7c) : $signed(_GEN_173); // @[NCOTable.scala 261:64]
  assign _GEN_175 = 7'h11 == cosAddr ? $signed(16'shd41) : $signed(_GEN_174); // @[NCOTable.scala 261:64]
  assign _GEN_176 = 7'h12 == cosAddr ? $signed(16'she06) : $signed(_GEN_175); // @[NCOTable.scala 261:64]
  assign _GEN_177 = 7'h13 == cosAddr ? $signed(16'sheca) : $signed(_GEN_176); // @[NCOTable.scala 261:64]
  assign _GEN_178 = 7'h14 == cosAddr ? $signed(16'shf8d) : $signed(_GEN_177); // @[NCOTable.scala 261:64]
  assign _GEN_179 = 7'h15 == cosAddr ? $signed(16'sh1050) : $signed(_GEN_178); // @[NCOTable.scala 261:64]
  assign _GEN_180 = 7'h16 == cosAddr ? $signed(16'sh1112) : $signed(_GEN_179); // @[NCOTable.scala 261:64]
  assign _GEN_181 = 7'h17 == cosAddr ? $signed(16'sh11d3) : $signed(_GEN_180); // @[NCOTable.scala 261:64]
  assign _GEN_182 = 7'h18 == cosAddr ? $signed(16'sh1294) : $signed(_GEN_181); // @[NCOTable.scala 261:64]
  assign _GEN_183 = 7'h19 == cosAddr ? $signed(16'sh1354) : $signed(_GEN_182); // @[NCOTable.scala 261:64]
  assign _GEN_184 = 7'h1a == cosAddr ? $signed(16'sh1413) : $signed(_GEN_183); // @[NCOTable.scala 261:64]
  assign _GEN_185 = 7'h1b == cosAddr ? $signed(16'sh14d2) : $signed(_GEN_184); // @[NCOTable.scala 261:64]
  assign _GEN_186 = 7'h1c == cosAddr ? $signed(16'sh1590) : $signed(_GEN_185); // @[NCOTable.scala 261:64]
  assign _GEN_187 = 7'h1d == cosAddr ? $signed(16'sh164c) : $signed(_GEN_186); // @[NCOTable.scala 261:64]
  assign _GEN_188 = 7'h1e == cosAddr ? $signed(16'sh1709) : $signed(_GEN_187); // @[NCOTable.scala 261:64]
  assign _GEN_189 = 7'h1f == cosAddr ? $signed(16'sh17c4) : $signed(_GEN_188); // @[NCOTable.scala 261:64]
  assign _GEN_190 = 7'h20 == cosAddr ? $signed(16'sh187e) : $signed(_GEN_189); // @[NCOTable.scala 261:64]
  assign _GEN_191 = 7'h21 == cosAddr ? $signed(16'sh1937) : $signed(_GEN_190); // @[NCOTable.scala 261:64]
  assign _GEN_192 = 7'h22 == cosAddr ? $signed(16'sh19ef) : $signed(_GEN_191); // @[NCOTable.scala 261:64]
  assign _GEN_193 = 7'h23 == cosAddr ? $signed(16'sh1aa7) : $signed(_GEN_192); // @[NCOTable.scala 261:64]
  assign _GEN_194 = 7'h24 == cosAddr ? $signed(16'sh1b5d) : $signed(_GEN_193); // @[NCOTable.scala 261:64]
  assign _GEN_195 = 7'h25 == cosAddr ? $signed(16'sh1c12) : $signed(_GEN_194); // @[NCOTable.scala 261:64]
  assign _GEN_196 = 7'h26 == cosAddr ? $signed(16'sh1cc6) : $signed(_GEN_195); // @[NCOTable.scala 261:64]
  assign _GEN_197 = 7'h27 == cosAddr ? $signed(16'sh1d79) : $signed(_GEN_196); // @[NCOTable.scala 261:64]
  assign _GEN_198 = 7'h28 == cosAddr ? $signed(16'sh1e2b) : $signed(_GEN_197); // @[NCOTable.scala 261:64]
  assign _GEN_199 = 7'h29 == cosAddr ? $signed(16'sh1edc) : $signed(_GEN_198); // @[NCOTable.scala 261:64]
  assign _GEN_200 = 7'h2a == cosAddr ? $signed(16'sh1f8c) : $signed(_GEN_199); // @[NCOTable.scala 261:64]
  assign _GEN_201 = 7'h2b == cosAddr ? $signed(16'sh203a) : $signed(_GEN_200); // @[NCOTable.scala 261:64]
  assign _GEN_202 = 7'h2c == cosAddr ? $signed(16'sh20e7) : $signed(_GEN_201); // @[NCOTable.scala 261:64]
  assign _GEN_203 = 7'h2d == cosAddr ? $signed(16'sh2193) : $signed(_GEN_202); // @[NCOTable.scala 261:64]
  assign _GEN_204 = 7'h2e == cosAddr ? $signed(16'sh223d) : $signed(_GEN_203); // @[NCOTable.scala 261:64]
  assign _GEN_205 = 7'h2f == cosAddr ? $signed(16'sh22e7) : $signed(_GEN_204); // @[NCOTable.scala 261:64]
  assign _GEN_206 = 7'h30 == cosAddr ? $signed(16'sh238e) : $signed(_GEN_205); // @[NCOTable.scala 261:64]
  assign _GEN_207 = 7'h31 == cosAddr ? $signed(16'sh2435) : $signed(_GEN_206); // @[NCOTable.scala 261:64]
  assign _GEN_208 = 7'h32 == cosAddr ? $signed(16'sh24da) : $signed(_GEN_207); // @[NCOTable.scala 261:64]
  assign _GEN_209 = 7'h33 == cosAddr ? $signed(16'sh257e) : $signed(_GEN_208); // @[NCOTable.scala 261:64]
  assign _GEN_210 = 7'h34 == cosAddr ? $signed(16'sh2620) : $signed(_GEN_209); // @[NCOTable.scala 261:64]
  assign _GEN_211 = 7'h35 == cosAddr ? $signed(16'sh26c1) : $signed(_GEN_210); // @[NCOTable.scala 261:64]
  assign _GEN_212 = 7'h36 == cosAddr ? $signed(16'sh2760) : $signed(_GEN_211); // @[NCOTable.scala 261:64]
  assign _GEN_213 = 7'h37 == cosAddr ? $signed(16'sh27fe) : $signed(_GEN_212); // @[NCOTable.scala 261:64]
  assign _GEN_214 = 7'h38 == cosAddr ? $signed(16'sh289a) : $signed(_GEN_213); // @[NCOTable.scala 261:64]
  assign _GEN_215 = 7'h39 == cosAddr ? $signed(16'sh2935) : $signed(_GEN_214); // @[NCOTable.scala 261:64]
  assign _GEN_216 = 7'h3a == cosAddr ? $signed(16'sh29ce) : $signed(_GEN_215); // @[NCOTable.scala 261:64]
  assign _GEN_217 = 7'h3b == cosAddr ? $signed(16'sh2a65) : $signed(_GEN_216); // @[NCOTable.scala 261:64]
  assign _GEN_218 = 7'h3c == cosAddr ? $signed(16'sh2afb) : $signed(_GEN_217); // @[NCOTable.scala 261:64]
  assign _GEN_219 = 7'h3d == cosAddr ? $signed(16'sh2b8f) : $signed(_GEN_218); // @[NCOTable.scala 261:64]
  assign _GEN_220 = 7'h3e == cosAddr ? $signed(16'sh2c21) : $signed(_GEN_219); // @[NCOTable.scala 261:64]
  assign _GEN_221 = 7'h3f == cosAddr ? $signed(16'sh2cb2) : $signed(_GEN_220); // @[NCOTable.scala 261:64]
  assign _GEN_222 = 7'h40 == cosAddr ? $signed(16'sh2d41) : $signed(_GEN_221); // @[NCOTable.scala 261:64]
  assign _GEN_223 = 7'h41 == cosAddr ? $signed(16'sh2dcf) : $signed(_GEN_222); // @[NCOTable.scala 261:64]
  assign _GEN_224 = 7'h42 == cosAddr ? $signed(16'sh2e5a) : $signed(_GEN_223); // @[NCOTable.scala 261:64]
  assign _GEN_225 = 7'h43 == cosAddr ? $signed(16'sh2ee4) : $signed(_GEN_224); // @[NCOTable.scala 261:64]
  assign _GEN_226 = 7'h44 == cosAddr ? $signed(16'sh2f6c) : $signed(_GEN_225); // @[NCOTable.scala 261:64]
  assign _GEN_227 = 7'h45 == cosAddr ? $signed(16'sh2ff2) : $signed(_GEN_226); // @[NCOTable.scala 261:64]
  assign _GEN_228 = 7'h46 == cosAddr ? $signed(16'sh3076) : $signed(_GEN_227); // @[NCOTable.scala 261:64]
  assign _GEN_229 = 7'h47 == cosAddr ? $signed(16'sh30f9) : $signed(_GEN_228); // @[NCOTable.scala 261:64]
  assign _GEN_230 = 7'h48 == cosAddr ? $signed(16'sh3179) : $signed(_GEN_229); // @[NCOTable.scala 261:64]
  assign _GEN_231 = 7'h49 == cosAddr ? $signed(16'sh31f8) : $signed(_GEN_230); // @[NCOTable.scala 261:64]
  assign _GEN_232 = 7'h4a == cosAddr ? $signed(16'sh3274) : $signed(_GEN_231); // @[NCOTable.scala 261:64]
  assign _GEN_233 = 7'h4b == cosAddr ? $signed(16'sh32ef) : $signed(_GEN_232); // @[NCOTable.scala 261:64]
  assign _GEN_234 = 7'h4c == cosAddr ? $signed(16'sh3368) : $signed(_GEN_233); // @[NCOTable.scala 261:64]
  assign _GEN_235 = 7'h4d == cosAddr ? $signed(16'sh33df) : $signed(_GEN_234); // @[NCOTable.scala 261:64]
  assign _GEN_236 = 7'h4e == cosAddr ? $signed(16'sh3453) : $signed(_GEN_235); // @[NCOTable.scala 261:64]
  assign _GEN_237 = 7'h4f == cosAddr ? $signed(16'sh34c6) : $signed(_GEN_236); // @[NCOTable.scala 261:64]
  assign _GEN_238 = 7'h50 == cosAddr ? $signed(16'sh3537) : $signed(_GEN_237); // @[NCOTable.scala 261:64]
  assign _GEN_239 = 7'h51 == cosAddr ? $signed(16'sh35a5) : $signed(_GEN_238); // @[NCOTable.scala 261:64]
  assign _GEN_240 = 7'h52 == cosAddr ? $signed(16'sh3612) : $signed(_GEN_239); // @[NCOTable.scala 261:64]
  assign _GEN_241 = 7'h53 == cosAddr ? $signed(16'sh367d) : $signed(_GEN_240); // @[NCOTable.scala 261:64]
  assign _GEN_242 = 7'h54 == cosAddr ? $signed(16'sh36e5) : $signed(_GEN_241); // @[NCOTable.scala 261:64]
  assign _GEN_243 = 7'h55 == cosAddr ? $signed(16'sh374b) : $signed(_GEN_242); // @[NCOTable.scala 261:64]
  assign _GEN_244 = 7'h56 == cosAddr ? $signed(16'sh37b0) : $signed(_GEN_243); // @[NCOTable.scala 261:64]
  assign _GEN_245 = 7'h57 == cosAddr ? $signed(16'sh3812) : $signed(_GEN_244); // @[NCOTable.scala 261:64]
  assign _GEN_246 = 7'h58 == cosAddr ? $signed(16'sh3871) : $signed(_GEN_245); // @[NCOTable.scala 261:64]
  assign _GEN_247 = 7'h59 == cosAddr ? $signed(16'sh38cf) : $signed(_GEN_246); // @[NCOTable.scala 261:64]
  assign _GEN_248 = 7'h5a == cosAddr ? $signed(16'sh392b) : $signed(_GEN_247); // @[NCOTable.scala 261:64]
  assign _GEN_249 = 7'h5b == cosAddr ? $signed(16'sh3984) : $signed(_GEN_248); // @[NCOTable.scala 261:64]
  assign _GEN_250 = 7'h5c == cosAddr ? $signed(16'sh39db) : $signed(_GEN_249); // @[NCOTable.scala 261:64]
  assign _GEN_251 = 7'h5d == cosAddr ? $signed(16'sh3a30) : $signed(_GEN_250); // @[NCOTable.scala 261:64]
  assign _GEN_252 = 7'h5e == cosAddr ? $signed(16'sh3a82) : $signed(_GEN_251); // @[NCOTable.scala 261:64]
  assign _GEN_253 = 7'h5f == cosAddr ? $signed(16'sh3ad3) : $signed(_GEN_252); // @[NCOTable.scala 261:64]
  assign _GEN_254 = 7'h60 == cosAddr ? $signed(16'sh3b21) : $signed(_GEN_253); // @[NCOTable.scala 261:64]
  assign _GEN_255 = 7'h61 == cosAddr ? $signed(16'sh3b6d) : $signed(_GEN_254); // @[NCOTable.scala 261:64]
  assign _GEN_256 = 7'h62 == cosAddr ? $signed(16'sh3bb6) : $signed(_GEN_255); // @[NCOTable.scala 261:64]
  assign _GEN_257 = 7'h63 == cosAddr ? $signed(16'sh3bfd) : $signed(_GEN_256); // @[NCOTable.scala 261:64]
  assign _GEN_258 = 7'h64 == cosAddr ? $signed(16'sh3c42) : $signed(_GEN_257); // @[NCOTable.scala 261:64]
  assign _GEN_259 = 7'h65 == cosAddr ? $signed(16'sh3c85) : $signed(_GEN_258); // @[NCOTable.scala 261:64]
  assign _GEN_260 = 7'h66 == cosAddr ? $signed(16'sh3cc5) : $signed(_GEN_259); // @[NCOTable.scala 261:64]
  assign _GEN_261 = 7'h67 == cosAddr ? $signed(16'sh3d03) : $signed(_GEN_260); // @[NCOTable.scala 261:64]
  assign _GEN_262 = 7'h68 == cosAddr ? $signed(16'sh3d3f) : $signed(_GEN_261); // @[NCOTable.scala 261:64]
  assign _GEN_263 = 7'h69 == cosAddr ? $signed(16'sh3d78) : $signed(_GEN_262); // @[NCOTable.scala 261:64]
  assign _GEN_264 = 7'h6a == cosAddr ? $signed(16'sh3daf) : $signed(_GEN_263); // @[NCOTable.scala 261:64]
  assign _GEN_265 = 7'h6b == cosAddr ? $signed(16'sh3de3) : $signed(_GEN_264); // @[NCOTable.scala 261:64]
  assign _GEN_266 = 7'h6c == cosAddr ? $signed(16'sh3e15) : $signed(_GEN_265); // @[NCOTable.scala 261:64]
  assign _GEN_267 = 7'h6d == cosAddr ? $signed(16'sh3e45) : $signed(_GEN_266); // @[NCOTable.scala 261:64]
  assign _GEN_268 = 7'h6e == cosAddr ? $signed(16'sh3e72) : $signed(_GEN_267); // @[NCOTable.scala 261:64]
  assign _GEN_269 = 7'h6f == cosAddr ? $signed(16'sh3e9d) : $signed(_GEN_268); // @[NCOTable.scala 261:64]
  assign _GEN_270 = 7'h70 == cosAddr ? $signed(16'sh3ec5) : $signed(_GEN_269); // @[NCOTable.scala 261:64]
  assign _GEN_271 = 7'h71 == cosAddr ? $signed(16'sh3eeb) : $signed(_GEN_270); // @[NCOTable.scala 261:64]
  assign _GEN_272 = 7'h72 == cosAddr ? $signed(16'sh3f0f) : $signed(_GEN_271); // @[NCOTable.scala 261:64]
  assign _GEN_273 = 7'h73 == cosAddr ? $signed(16'sh3f30) : $signed(_GEN_272); // @[NCOTable.scala 261:64]
  assign _GEN_274 = 7'h74 == cosAddr ? $signed(16'sh3f4f) : $signed(_GEN_273); // @[NCOTable.scala 261:64]
  assign _GEN_275 = 7'h75 == cosAddr ? $signed(16'sh3f6b) : $signed(_GEN_274); // @[NCOTable.scala 261:64]
  assign _GEN_276 = 7'h76 == cosAddr ? $signed(16'sh3f85) : $signed(_GEN_275); // @[NCOTable.scala 261:64]
  assign _GEN_277 = 7'h77 == cosAddr ? $signed(16'sh3f9c) : $signed(_GEN_276); // @[NCOTable.scala 261:64]
  assign _GEN_278 = 7'h78 == cosAddr ? $signed(16'sh3fb1) : $signed(_GEN_277); // @[NCOTable.scala 261:64]
  assign _GEN_279 = 7'h79 == cosAddr ? $signed(16'sh3fc4) : $signed(_GEN_278); // @[NCOTable.scala 261:64]
  assign _GEN_280 = 7'h7a == cosAddr ? $signed(16'sh3fd4) : $signed(_GEN_279); // @[NCOTable.scala 261:64]
  assign _GEN_281 = 7'h7b == cosAddr ? $signed(16'sh3fe1) : $signed(_GEN_280); // @[NCOTable.scala 261:64]
  assign _GEN_282 = 7'h7c == cosAddr ? $signed(16'sh3fec) : $signed(_GEN_281); // @[NCOTable.scala 261:64]
  assign _GEN_283 = 7'h7d == cosAddr ? $signed(16'sh3ff5) : $signed(_GEN_282); // @[NCOTable.scala 261:64]
  assign _GEN_284 = 7'h7e == cosAddr ? $signed(16'sh3ffb) : $signed(_GEN_283); // @[NCOTable.scala 261:64]
  assign _T_71 = 7'h7f == cosAddr ? $signed(16'sh3fff) : $signed(_GEN_284); // @[NCOTable.scala 261:64]
  assign cosTableOut = _GEN_26 ? $signed(16'sh4000) : $signed(_T_71); // @[NCOTable.scala 261:23]
  assign _T_75 = 16'sh0 - $signed(sinTableOut); // @[FixedPointTypeClass.scala 39:43]
  assign _T_78 = 16'sh0 - $signed(cosTableOut); // @[FixedPointTypeClass.scala 39:43]
  assign io_sinOut = sinNegative2 ? $signed(_T_75) : $signed(sinTableOut); // @[NCOTable.scala 314:13]
  assign io_cosOut = cosNegative2 ? $signed(_T_78) : $signed(cosTableOut); // @[NCOTable.scala 315:13]
endmodule
module NCOTable(
  input  [8:0]  io_phase,
  output [15:0] io_sinOut,
  output [15:0] io_cosOut
);
  wire [8:0] tableNCO_io_phase; // @[NCOTable.scala 473:13]
  wire [15:0] tableNCO_io_sinOut; // @[NCOTable.scala 473:13]
  wire [15:0] tableNCO_io_cosOut; // @[NCOTable.scala 473:13]
  NCOTableStandardMode tableNCO ( // @[NCOTable.scala 473:13]
    .io_phase(tableNCO_io_phase),
    .io_sinOut(tableNCO_io_sinOut),
    .io_cosOut(tableNCO_io_cosOut)
  );
  assign io_sinOut = tableNCO_io_sinOut; // @[NCOTable.scala 478:13]
  assign io_cosOut = tableNCO_io_cosOut; // @[NCOTable.scala 479:13]
  assign tableNCO_io_phase = io_phase; // @[NCOTable.scala 477:21]
endmodule
module Queue_6(
  input   clock,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input   io_enq_bits,
  input   io_deq_ready,
  output  io_deq_valid,
  output  io_deq_bits
);
  reg  _T [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_0;
  wire  _T__T_18_data; // @[Decoupled.scala 209:24]
  wire  _T__T_18_addr; // @[Decoupled.scala 209:24]
  wire  _T__T_10_data; // @[Decoupled.scala 209:24]
  wire  _T__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T__T_10_en; // @[Decoupled.scala 209:24]
  reg  value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_1;
  reg  value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_2;
  reg  _T_1; // @[Decoupled.scala 212:35]
  reg [31:0] _RAND_3;
  wire  _T_2; // @[Decoupled.scala 214:41]
  wire  _T_3; // @[Decoupled.scala 215:36]
  wire  _T_4; // @[Decoupled.scala 215:33]
  wire  _T_5; // @[Decoupled.scala 216:32]
  wire  _T_6; // @[Decoupled.scala 40:37]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _T_12; // @[Counter.scala 39:22]
  wire  _T_14; // @[Counter.scala 39:22]
  wire  _T_15; // @[Decoupled.scala 227:16]
  wire  _T_17; // @[Decoupled.scala 232:19]
  assign _T__T_18_addr = value_1;
  assign _T__T_18_data = _T[_T__T_18_addr]; // @[Decoupled.scala 209:24]
  assign _T__T_10_data = io_enq_bits;
  assign _T__T_10_addr = value;
  assign _T__T_10_mask = 1'h1;
  assign _T__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_2 = value == value_1; // @[Decoupled.scala 214:41]
  assign _T_3 = ~_T_1; // @[Decoupled.scala 215:36]
  assign _T_4 = _T_2 & _T_3; // @[Decoupled.scala 215:33]
  assign _T_5 = _T_2 & _T_1; // @[Decoupled.scala 216:32]
  assign _T_6 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  assign _T_8 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  assign _T_12 = value + 1'h1; // @[Counter.scala 39:22]
  assign _T_14 = value_1 + 1'h1; // @[Counter.scala 39:22]
  assign _T_15 = _T_6 != _T_8; // @[Decoupled.scala 227:16]
  assign _T_17 = ~_T_5; // @[Decoupled.scala 232:19]
  assign io_enq_ready = io_deq_ready | _T_17; // @[Decoupled.scala 232:16 Decoupled.scala 245:40]
  assign io_deq_valid = ~_T_4; // @[Decoupled.scala 231:16]
  assign io_deq_bits = _T__T_18_data; // @[Decoupled.scala 233:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T[initvar] = _RAND_0[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  value = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  value_1 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_1 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T__T_10_en & _T__T_10_mask) begin
      _T[_T__T_10_addr] <= _T__T_10_data; // @[Decoupled.scala 209:24]
    end
    if (reset) begin
      value <= 1'h0;
    end else if (_T_6) begin
      value <= _T_12;
    end
    if (reset) begin
      value_1 <= 1'h0;
    end else if (_T_8) begin
      value_1 <= _T_14;
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else if (_T_15) begin
      _T_1 <= _T_6;
    end
  end
endmodule
module AXI4NCOLazyModuleBlock(
  input         clock,
  input         reset,
  input         auto_stream_out_ready,
  output        auto_stream_out_valid,
  output [31:0] auto_stream_out_bits_data,
  output        auto_stream_out_bits_last,
  output        auto_freq_in_ready,
  input         auto_freq_in_valid,
  input  [31:0] auto_freq_in_bits_data,
  input         auto_freq_in_bits_last
);
  wire [8:0] phaseConverter_io_phase; // @[NCOLazyModuleBlock.scala 35:32]
  wire [15:0] phaseConverter_io_sinOut; // @[NCOLazyModuleBlock.scala 35:32]
  wire [15:0] phaseConverter_io_cosOut; // @[NCOLazyModuleBlock.scala 35:32]
  wire  Queue_clock; // @[Skid.scala 21:23]
  wire  Queue_reset; // @[Skid.scala 21:23]
  wire  Queue_io_enq_ready; // @[Skid.scala 21:23]
  wire  Queue_io_enq_valid; // @[Skid.scala 21:23]
  wire  Queue_io_enq_bits; // @[Skid.scala 21:23]
  wire  Queue_io_deq_ready; // @[Skid.scala 21:23]
  wire  Queue_io_deq_valid; // @[Skid.scala 21:23]
  wire  Queue_io_deq_bits; // @[Skid.scala 21:23]
  reg [8:0] phaseCounter; // @[NCOLazyModuleBlock.scala 36:33]
  reg [31:0] _RAND_0;
  reg [1:0] _T_35; // @[NCOLazyModuleBlock.scala 213:33]
  reg [31:0] _RAND_1;
  wire  _T_52; // @[NCOLazyModuleBlock.scala 223:48]
  wire  _T_53; // @[NCOLazyModuleBlock.scala 223:78]
  wire  _T_54; // @[NCOLazyModuleBlock.scala 223:92]
  wire  _T_55; // @[NCOLazyModuleBlock.scala 223:61]
  wire  _T_5; // @[Decoupled.scala 40:37]
  wire [31:0] _GEN_15; // @[NCOLazyModuleBlock.scala 190:40]
  wire [31:0] _T_7; // @[NCOLazyModuleBlock.scala 190:40]
  wire [31:0] _GEN_0; // @[NCOLazyModuleBlock.scala 189:40]
  wire [16:0] _T_8; // @[NCOLazyModuleBlock.scala 199:47]
  reg  queueCounter; // @[Skid.scala 22:31]
  reg [31:0] _RAND_2;
  wire  _T_26; // @[Skid.scala 29:31]
  wire  _T_28; // @[Skid.scala 29:75]
  wire  _T_29; // @[Skid.scala 29:44]
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire [1:0] _T_15; // @[Skid.scala 23:34]
  wire  _T_11_valid; // @[NCOLazyModuleBlock.scala 202:29 Skid.scala 31:15]
  wire  _T_16; // @[Decoupled.scala 40:37]
  wire [1:0] _GEN_16; // @[Skid.scala 23:47]
  wire [2:0] _T_17; // @[Skid.scala 23:47]
  reg  _T_20; // @[Reg.scala 27:20]
  reg [31:0] _RAND_3;
  wire  _T_21; // @[Skid.scala 26:12]
  wire  _T_22; // @[Skid.scala 26:32]
  wire  _T_24; // @[Skid.scala 26:11]
  wire  _T_25; // @[Skid.scala 26:11]
  reg  ioout_bits_last; // @[NCOLazyModuleBlock.scala 207:28]
  reg [31:0] _RAND_4;
  reg  _T_31; // @[NCOLazyModuleBlock.scala 208:30]
  reg [31:0] _RAND_5;
  wire  _T_11_bits; // @[NCOLazyModuleBlock.scala 202:29 Skid.scala 32:14]
  wire  _GEN_2; // @[NCOLazyModuleBlock.scala 209:30]
  wire  _T_32; // @[NCOLazyModuleBlock.scala 210:32]
  wire  _T_33; // @[NCOLazyModuleBlock.scala 210:29]
  wire  _T_57; // @[NCOLazyModuleBlock.scala 224:65]
  reg [1:0] _T_46; // @[NCOLazyModuleBlock.scala 218:64]
  reg [31:0] _RAND_6;
  wire  _T_47; // @[NCOLazyModuleBlock.scala 218:53]
  reg [1:0] _T_48; // @[NCOLazyModuleBlock.scala 218:87]
  reg [31:0] _RAND_7;
  reg [1:0] _T_41; // @[NCOLazyModuleBlock.scala 215:42]
  reg [31:0] _RAND_8;
  wire [1:0] _T_49; // @[NCOLazyModuleBlock.scala 218:39]
  wire  _T_58; // @[NCOLazyModuleBlock.scala 224:104]
  wire  _T_59; // @[NCOLazyModuleBlock.scala 224:74]
  wire  _T_60; // @[NCOLazyModuleBlock.scala 224:47]
  wire  ioout_valid; // @[NCOLazyModuleBlock.scala 224:115]
  wire [1:0] _GEN_17; // @[NCOLazyModuleBlock.scala 214:36]
  wire [2:0] _T_37; // @[NCOLazyModuleBlock.scala 214:36]
  wire  _T_38; // @[Decoupled.scala 40:37]
  wire [2:0] _GEN_18; // @[NCOLazyModuleBlock.scala 214:64]
  wire [3:0] _T_39; // @[NCOLazyModuleBlock.scala 214:64]
  reg [1:0] _T_42; // @[NCOLazyModuleBlock.scala 216:37]
  reg [31:0] _RAND_9;
  wire  _T_43; // @[NCOLazyModuleBlock.scala 216:26]
  reg [1:0] _T_44; // @[NCOLazyModuleBlock.scala 216:86]
  reg [31:0] _RAND_10;
  reg  _T_50; // @[NCOLazyModuleBlock.scala 220:27]
  reg [31:0] _RAND_11;
  reg [15:0] _T_64; // @[NCOLazyModuleBlock.scala 226:36]
  reg [31:0] _RAND_12;
  reg [15:0] _T_67; // @[NCOLazyModuleBlock.scala 227:36]
  reg [31:0] _RAND_13;
  reg [15:0] _T_70; // @[NCOLazyModuleBlock.scala 229:37]
  reg [31:0] _RAND_14;
  reg [15:0] _T_73; // @[NCOLazyModuleBlock.scala 230:37]
  reg [31:0] _RAND_15;
  wire  _T_76; // @[NCOLazyModuleBlock.scala 258:39]
  wire [31:0] _T_79; // @[Cat.scala 29:58]
  wire  _T_81; // @[NCOLazyModuleBlock.scala 260:48]
  wire  _T_82; // @[NCOLazyModuleBlock.scala 260:45]
  wire [31:0] _T_85; // @[Cat.scala 29:58]
  wire  _T_87; // @[NCOLazyModuleBlock.scala 262:20]
  wire  _T_88; // @[NCOLazyModuleBlock.scala 262:46]
  wire [31:0] _GEN_11; // @[NCOLazyModuleBlock.scala 262:56]
  wire [31:0] _GEN_12; // @[NCOLazyModuleBlock.scala 260:56]
  wire [31:0] _GEN_13; // @[NCOLazyModuleBlock.scala 258:49]
  NCOTable phaseConverter ( // @[NCOLazyModuleBlock.scala 35:32]
    .io_phase(phaseConverter_io_phase),
    .io_sinOut(phaseConverter_io_sinOut),
    .io_cosOut(phaseConverter_io_cosOut)
  );
  Queue_6 Queue ( // @[Skid.scala 21:23]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits(Queue_io_enq_bits),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits(Queue_io_deq_bits)
  );
  assign _T_52 = _T_35 < 2'h2; // @[NCOLazyModuleBlock.scala 223:48]
  assign _T_53 = _T_35 == 2'h2; // @[NCOLazyModuleBlock.scala 223:78]
  assign _T_54 = _T_53 & auto_stream_out_ready; // @[NCOLazyModuleBlock.scala 223:92]
  assign _T_55 = _T_52 | _T_54; // @[NCOLazyModuleBlock.scala 223:61]
  assign _T_5 = _T_55 & auto_freq_in_valid; // @[Decoupled.scala 40:37]
  assign _GEN_15 = {{23'd0}, phaseCounter}; // @[NCOLazyModuleBlock.scala 190:40]
  assign _T_7 = _GEN_15 + auto_freq_in_bits_data; // @[NCOLazyModuleBlock.scala 190:40]
  assign _GEN_0 = _T_5 ? _T_7 : {{23'd0}, phaseCounter}; // @[NCOLazyModuleBlock.scala 189:40]
  assign _T_8 = {{8'd0}, phaseCounter}; // @[NCOLazyModuleBlock.scala 199:47]
  assign _T_26 = queueCounter < 1'h1; // @[Skid.scala 29:31]
  assign _T_28 = queueCounter & auto_stream_out_ready; // @[Skid.scala 29:75]
  assign _T_29 = _T_26 | _T_28; // @[Skid.scala 29:44]
  assign _T_14 = _T_29 & auto_freq_in_valid; // @[Decoupled.scala 40:37]
  assign _T_15 = queueCounter + _T_14; // @[Skid.scala 23:34]
  assign _T_11_valid = Queue_io_deq_valid; // @[NCOLazyModuleBlock.scala 202:29 Skid.scala 31:15]
  assign _T_16 = auto_stream_out_ready & _T_11_valid; // @[Decoupled.scala 40:37]
  assign _GEN_16 = {{1'd0}, _T_16}; // @[Skid.scala 23:47]
  assign _T_17 = _T_15 - _GEN_16; // @[Skid.scala 23:47]
  assign _T_21 = ~Queue_io_enq_valid; // @[Skid.scala 26:12]
  assign _T_22 = _T_21 | Queue_io_enq_ready; // @[Skid.scala 26:32]
  assign _T_24 = _T_22 | reset; // @[Skid.scala 26:11]
  assign _T_25 = ~_T_24; // @[Skid.scala 26:11]
  assign _T_11_bits = Queue_io_deq_bits; // @[NCOLazyModuleBlock.scala 202:29 Skid.scala 32:14]
  assign _GEN_2 = _T_11_bits | _T_31; // @[NCOLazyModuleBlock.scala 209:30]
  assign _T_32 = ~_T_31; // @[NCOLazyModuleBlock.scala 210:32]
  assign _T_33 = _T_11_bits & _T_32; // @[NCOLazyModuleBlock.scala 210:29]
  assign _T_57 = _T_35 == 2'h1; // @[NCOLazyModuleBlock.scala 224:65]
  assign _T_47 = _T_35 != _T_46; // @[NCOLazyModuleBlock.scala 218:53]
  assign _T_49 = _T_47 ? _T_48 : _T_41; // @[NCOLazyModuleBlock.scala 218:39]
  assign _T_58 = _T_49 == 2'h2; // @[NCOLazyModuleBlock.scala 224:104]
  assign _T_59 = _T_57 & _T_58; // @[NCOLazyModuleBlock.scala 224:74]
  assign _T_60 = _T_53 | _T_59; // @[NCOLazyModuleBlock.scala 224:47]
  assign ioout_valid = _T_60 & auto_stream_out_ready; // @[NCOLazyModuleBlock.scala 224:115]
  assign _GEN_17 = {{1'd0}, _T_5}; // @[NCOLazyModuleBlock.scala 214:36]
  assign _T_37 = _T_35 + _GEN_17; // @[NCOLazyModuleBlock.scala 214:36]
  assign _T_38 = auto_stream_out_ready & ioout_valid; // @[Decoupled.scala 40:37]
  assign _GEN_18 = {{2'd0}, _T_38}; // @[NCOLazyModuleBlock.scala 214:64]
  assign _T_39 = _T_37 - _GEN_18; // @[NCOLazyModuleBlock.scala 214:64]
  assign _T_43 = _T_35 != _T_42; // @[NCOLazyModuleBlock.scala 216:26]
  assign _T_76 = _T_5 & _T_50; // @[NCOLazyModuleBlock.scala 258:39]
  assign _T_79 = {_T_67,_T_64}; // @[Cat.scala 29:58]
  assign _T_81 = ~_T_50; // @[NCOLazyModuleBlock.scala 260:48]
  assign _T_82 = _T_5 & _T_81; // @[NCOLazyModuleBlock.scala 260:45]
  assign _T_85 = {_T_73,_T_70}; // @[Cat.scala 29:58]
  assign _T_87 = ~_T_5; // @[NCOLazyModuleBlock.scala 262:20]
  assign _T_88 = _T_87 & _T_50; // @[NCOLazyModuleBlock.scala 262:46]
  assign _GEN_11 = _T_88 ? _T_79 : _T_85; // @[NCOLazyModuleBlock.scala 262:56]
  assign _GEN_12 = _T_82 ? _T_85 : _GEN_11; // @[NCOLazyModuleBlock.scala 260:56]
  assign _GEN_13 = _T_76 ? _T_79 : _GEN_12; // @[NCOLazyModuleBlock.scala 258:49]
  assign auto_stream_out_valid = _T_60 & auto_stream_out_ready; // @[LazyModule.scala 173:49]
  assign auto_stream_out_bits_data = _T_53 ? _GEN_13 : _T_79; // @[LazyModule.scala 173:49]
  assign auto_stream_out_bits_last = ioout_bits_last; // @[LazyModule.scala 173:49]
  assign auto_freq_in_ready = _T_52 | _T_54; // @[LazyModule.scala 173:31]
  assign phaseConverter_io_phase = _T_8[8:0]; // @[NCOLazyModuleBlock.scala 199:31]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = _T_20; // @[Skid.scala 25:24]
  assign Queue_io_enq_bits = auto_freq_in_bits_last & _T_5; // @[NCOLazyModuleBlock.scala 206:41]
  assign Queue_io_deq_ready = auto_stream_out_ready; // @[Skid.scala 30:24]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  phaseCounter = _RAND_0[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_35 = _RAND_1[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  queueCounter = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_20 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  ioout_bits_last = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_31 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_46 = _RAND_6[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_48 = _RAND_7[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_41 = _RAND_8[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_42 = _RAND_9[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_44 = _RAND_10[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_50 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_64 = _RAND_12[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_67 = _RAND_13[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_70 = _RAND_14[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_73 = _RAND_15[15:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      phaseCounter <= 9'h0;
    end else begin
      phaseCounter <= _GEN_0[8:0];
    end
    if (reset) begin
      _T_35 <= 2'h0;
    end else begin
      _T_35 <= _T_39[1:0];
    end
    if (reset) begin
      queueCounter <= 1'h0;
    end else begin
      queueCounter <= _T_17[0];
    end
    if (reset) begin
      _T_20 <= 1'h0;
    end else begin
      _T_20 <= _T_14;
    end
    if (reset) begin
      ioout_bits_last <= 1'h0;
    end else begin
      ioout_bits_last <= _T_33;
    end
    if (reset) begin
      _T_31 <= 1'h0;
    end else begin
      _T_31 <= _GEN_2;
    end
    _T_46 <= _T_35;
    _T_48 <= _T_35;
    if (reset) begin
      _T_41 <= 2'h0;
    end else if (_T_43) begin
      _T_41 <= _T_44;
    end
    _T_42 <= _T_35;
    _T_44 <= _T_35;
    if (reset) begin
      _T_50 <= 1'h0;
    end else begin
      _T_50 <= _T_5;
    end
    if (reset) begin
      _T_64 <= 16'sh0;
    end else if (_T_50) begin
      _T_64 <= phaseConverter_io_sinOut;
    end
    if (reset) begin
      _T_67 <= 16'sh0;
    end else if (_T_50) begin
      _T_67 <= phaseConverter_io_cosOut;
    end
    if (reset) begin
      _T_70 <= 16'sh0;
    end else if (_T_50) begin
      _T_70 <= _T_64;
    end
    if (reset) begin
      _T_73 <= 16'sh0;
    end else if (_T_50) begin
      _T_73 <= _T_67;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_25) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Skid.scala:26 assert(!queue.io.enq.valid || queue.io.enq.ready) // we control in.ready such that the queue can't fill up!\n"); // @[Skid.scala 26:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_25) begin
          $fatal; // @[Skid.scala 26:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module AXI4Splitter_2(
  input         clock,
  input         reset,
  output        auto_mem_in_aw_ready,
  input         auto_mem_in_aw_valid,
  input         auto_mem_in_aw_bits_id,
  input  [29:0] auto_mem_in_aw_bits_addr,
  output        auto_mem_in_w_ready,
  input         auto_mem_in_w_valid,
  input  [31:0] auto_mem_in_w_bits_data,
  input  [3:0]  auto_mem_in_w_bits_strb,
  input         auto_mem_in_b_ready,
  output        auto_mem_in_b_valid,
  output        auto_mem_in_b_bits_id,
  output        auto_mem_in_ar_ready,
  input         auto_mem_in_ar_valid,
  input         auto_mem_in_ar_bits_id,
  input  [29:0] auto_mem_in_ar_bits_addr,
  input  [2:0]  auto_mem_in_ar_bits_size,
  input         auto_mem_in_r_ready,
  output        auto_mem_in_r_valid,
  output        auto_mem_in_r_bits_id,
  output [31:0] auto_mem_in_r_bits_data,
  output        auto_stream_in_ready,
  input         auto_stream_in_valid,
  input  [31:0] auto_stream_in_bits_data,
  input         auto_stream_in_bits_last,
  input         auto_stream_out_1_ready,
  output        auto_stream_out_1_valid,
  output [31:0] auto_stream_out_1_bits_data,
  output        auto_stream_out_1_bits_last,
  input         auto_stream_out_0_ready,
  output        auto_stream_out_0_valid,
  output [31:0] auto_stream_out_0_bits_data,
  output        auto_stream_out_0_bits_last
);
  wire  Queue_clock; // @[Decoupled.scala 287:21]
  wire  Queue_reset; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_read; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_enq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_extra; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_read; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_deq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_extra; // @[Decoupled.scala 287:21]
  reg [31:0] ctrlReg; // @[Splitter.scala 27:26]
  reg [31:0] _RAND_0;
  reg [31:0] maskReg; // @[Splitter.scala 28:26]
  reg [31:0] _RAND_1;
  wire  _T_4; // @[RegisterRouter.scala 40:39]
  wire  _T_5; // @[RegisterRouter.scala 40:26]
  wire  _T_6; // @[RegisterRouter.scala 42:29]
  wire  _T_49_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 290:17]
  wire [29:0] _T_13; // @[RegisterRouter.scala 48:19]
  wire [1:0] _T_53; // @[RegisterRouter.scala 59:16]
  wire  _T_55; // @[RegisterRouter.scala 59:16]
  wire  _T_7; // @[RegisterRouter.scala 42:26]
  wire [1:0] _T_16; // @[OneHot.scala 65:12]
  wire [1:0] _T_18; // @[Misc.scala 200:81]
  wire  _T_19; // @[Misc.scala 204:21]
  wire  _T_22; // @[Misc.scala 209:20]
  wire  _T_24; // @[Misc.scala 213:38]
  wire  _T_25; // @[Misc.scala 213:29]
  wire  _T_27; // @[Misc.scala 213:38]
  wire  _T_28; // @[Misc.scala 213:29]
  wire  _T_31; // @[Misc.scala 209:20]
  wire  _T_32; // @[Misc.scala 212:27]
  wire  _T_33; // @[Misc.scala 213:38]
  wire  _T_34; // @[Misc.scala 213:29]
  wire  _T_35; // @[Misc.scala 212:27]
  wire  _T_36; // @[Misc.scala 213:38]
  wire  _T_37; // @[Misc.scala 213:29]
  wire  _T_38; // @[Misc.scala 212:27]
  wire  _T_39; // @[Misc.scala 213:38]
  wire  _T_40; // @[Misc.scala 213:29]
  wire  _T_41; // @[Misc.scala 212:27]
  wire  _T_42; // @[Misc.scala 213:38]
  wire  _T_43; // @[Misc.scala 213:29]
  wire [3:0] _T_46; // @[Cat.scala 29:58]
  wire [3:0] _T_48; // @[RegisterRouter.scala 54:25]
  wire [7:0] _T_67; // @[Bitwise.scala 72:12]
  wire [7:0] _T_69; // @[Bitwise.scala 72:12]
  wire [7:0] _T_71; // @[Bitwise.scala 72:12]
  wire [7:0] _T_73; // @[Bitwise.scala 72:12]
  wire [31:0] _T_76; // @[Cat.scala 29:58]
  wire  _T_95; // @[RegisterRouter.scala 59:16]
  wire  _T_148; // @[RegisterRouter.scala 59:16]
  wire [1:0] _T_142; // @[OneHot.scala 58:35]
  wire  _T_165; // @[RegisterRouter.scala 59:16]
  wire  _T_172; // @[RegisterRouter.scala 59:16]
  wire  _T_173; // @[RegisterRouter.scala 59:16]
  wire  _T_102; // @[RegisterRouter.scala 59:16]
  wire  _T_167; // @[RegisterRouter.scala 59:16]
  wire  _T_168; // @[RegisterRouter.scala 59:16]
  wire  _T_125; // @[RegisterRouter.scala 59:16]
  wire  _GEN_11; // @[MuxLiteral.scala 48:10]
  wire [31:0] _GEN_13; // @[MuxLiteral.scala 48:10]
  wire  _T_223_bits_read; // @[Decoupled.scala 308:19 Decoupled.scala 309:14]
  wire  _T_223_valid; // @[Decoupled.scala 308:19 Decoupled.scala 310:15]
  wire  _T_226; // @[RegisterRouter.scala 65:29]
  wire  readyOR; // @[Splitter.scala 45:34]
  wire  readyAND; // @[Splitter.scala 46:34]
  wire  _T_229; // @[Splitter.scala 49:19]
  wire  _T_230; // @[Splitter.scala 52:24]
  wire  _GEN_14; // @[Splitter.scala 52:33]
  wire  _T_233; // @[Splitter.scala 62:34]
  wire  _T_237; // @[Splitter.scala 62:34]
  Queue Queue ( // @[Decoupled.scala 287:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_read(Queue_io_enq_bits_read),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_extra(Queue_io_enq_bits_extra),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_read(Queue_io_deq_bits_read),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_extra(Queue_io_deq_bits_extra)
  );
  assign _T_4 = auto_mem_in_aw_valid & auto_mem_in_w_valid; // @[RegisterRouter.scala 40:39]
  assign _T_5 = auto_mem_in_ar_valid | _T_4; // @[RegisterRouter.scala 40:26]
  assign _T_6 = ~auto_mem_in_ar_valid; // @[RegisterRouter.scala 42:29]
  assign _T_49_ready = Queue_io_enq_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 290:17]
  assign _T_13 = auto_mem_in_ar_valid ? auto_mem_in_ar_bits_addr : auto_mem_in_aw_bits_addr; // @[RegisterRouter.scala 48:19]
  assign _T_53 = _T_13[3:2] & 2'h2; // @[RegisterRouter.scala 59:16]
  assign _T_55 = _T_53 == 2'h0; // @[RegisterRouter.scala 59:16]
  assign _T_7 = _T_49_ready & _T_6; // @[RegisterRouter.scala 42:26]
  assign _T_16 = 2'h1 << auto_mem_in_ar_bits_size[0]; // @[OneHot.scala 65:12]
  assign _T_18 = _T_16 | 2'h1; // @[Misc.scala 200:81]
  assign _T_19 = auto_mem_in_ar_bits_size >= 3'h2; // @[Misc.scala 204:21]
  assign _T_22 = ~auto_mem_in_ar_bits_addr[1]; // @[Misc.scala 209:20]
  assign _T_24 = _T_18[1] & _T_22; // @[Misc.scala 213:38]
  assign _T_25 = _T_19 | _T_24; // @[Misc.scala 213:29]
  assign _T_27 = _T_18[1] & auto_mem_in_ar_bits_addr[1]; // @[Misc.scala 213:38]
  assign _T_28 = _T_19 | _T_27; // @[Misc.scala 213:29]
  assign _T_31 = ~auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 209:20]
  assign _T_32 = _T_22 & _T_31; // @[Misc.scala 212:27]
  assign _T_33 = _T_18[0] & _T_32; // @[Misc.scala 213:38]
  assign _T_34 = _T_25 | _T_33; // @[Misc.scala 213:29]
  assign _T_35 = _T_22 & auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  assign _T_36 = _T_18[0] & _T_35; // @[Misc.scala 213:38]
  assign _T_37 = _T_25 | _T_36; // @[Misc.scala 213:29]
  assign _T_38 = auto_mem_in_ar_bits_addr[1] & _T_31; // @[Misc.scala 212:27]
  assign _T_39 = _T_18[0] & _T_38; // @[Misc.scala 213:38]
  assign _T_40 = _T_28 | _T_39; // @[Misc.scala 213:29]
  assign _T_41 = auto_mem_in_ar_bits_addr[1] & auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  assign _T_42 = _T_18[0] & _T_41; // @[Misc.scala 213:38]
  assign _T_43 = _T_28 | _T_42; // @[Misc.scala 213:29]
  assign _T_46 = {_T_43,_T_40,_T_37,_T_34}; // @[Cat.scala 29:58]
  assign _T_48 = auto_mem_in_ar_valid ? _T_46 : auto_mem_in_w_bits_strb; // @[RegisterRouter.scala 54:25]
  assign _T_67 = _T_48[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_69 = _T_48[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_71 = _T_48[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_73 = _T_48[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_76 = {_T_73,_T_71,_T_69,_T_67}; // @[Cat.scala 29:58]
  assign _T_95 = _T_76 == 32'hffffffff; // @[RegisterRouter.scala 59:16]
  assign _T_148 = _T_5 & _T_49_ready; // @[RegisterRouter.scala 59:16]
  assign _T_142 = 2'h1 << _T_13[2]; // @[OneHot.scala 58:35]
  assign _T_165 = _T_148 & _T_6; // @[RegisterRouter.scala 59:16]
  assign _T_172 = _T_165 & _T_142[1]; // @[RegisterRouter.scala 59:16]
  assign _T_173 = _T_172 & _T_55; // @[RegisterRouter.scala 59:16]
  assign _T_102 = _T_173 & _T_95; // @[RegisterRouter.scala 59:16]
  assign _T_167 = _T_165 & _T_142[0]; // @[RegisterRouter.scala 59:16]
  assign _T_168 = _T_167 & _T_55; // @[RegisterRouter.scala 59:16]
  assign _T_125 = _T_168 & _T_95; // @[RegisterRouter.scala 59:16]
  assign _GEN_11 = _T_13[2] ? _T_55 : _T_55; // @[MuxLiteral.scala 48:10]
  assign _GEN_13 = _T_13[2] ? maskReg : ctrlReg; // @[MuxLiteral.scala 48:10]
  assign _T_223_bits_read = Queue_io_deq_bits_read; // @[Decoupled.scala 308:19 Decoupled.scala 309:14]
  assign _T_223_valid = Queue_io_deq_valid; // @[Decoupled.scala 308:19 Decoupled.scala 310:15]
  assign _T_226 = ~_T_223_bits_read; // @[RegisterRouter.scala 65:29]
  assign readyOR = auto_stream_out_0_ready | auto_stream_out_1_ready; // @[Splitter.scala 45:34]
  assign readyAND = auto_stream_out_0_ready & auto_stream_out_1_ready; // @[Splitter.scala 46:34]
  assign _T_229 = ctrlReg == 32'h0; // @[Splitter.scala 49:19]
  assign _T_230 = ctrlReg == 32'h1; // @[Splitter.scala 52:24]
  assign _GEN_14 = _T_230 & readyOR; // @[Splitter.scala 52:33]
  assign _T_233 = ~maskReg[0]; // @[Splitter.scala 62:34]
  assign _T_237 = ~maskReg[1]; // @[Splitter.scala 62:34]
  assign auto_mem_in_aw_ready = _T_7 & auto_mem_in_w_valid; // @[LazyModule.scala 173:31]
  assign auto_mem_in_w_ready = _T_7 & auto_mem_in_aw_valid; // @[LazyModule.scala 173:31]
  assign auto_mem_in_b_valid = _T_223_valid & _T_226; // @[LazyModule.scala 173:31]
  assign auto_mem_in_b_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_mem_in_ar_ready = Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_valid = _T_223_valid & _T_223_bits_read; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 173:31]
  assign auto_stream_in_ready = _T_229 ? readyAND : _GEN_14; // @[LazyModule.scala 173:31]
  assign auto_stream_out_1_valid = auto_stream_in_valid & _T_237; // @[LazyModule.scala 173:49]
  assign auto_stream_out_1_bits_data = auto_stream_in_bits_data; // @[LazyModule.scala 173:49]
  assign auto_stream_out_1_bits_last = auto_stream_in_bits_last; // @[LazyModule.scala 173:49]
  assign auto_stream_out_0_valid = auto_stream_in_valid & _T_233; // @[LazyModule.scala 173:49]
  assign auto_stream_out_0_bits_data = auto_stream_in_bits_data; // @[LazyModule.scala 173:49]
  assign auto_stream_out_0_bits_last = auto_stream_in_bits_last; // @[LazyModule.scala 173:49]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_mem_in_ar_valid | _T_4; // @[Decoupled.scala 288:22]
  assign Queue_io_enq_bits_read = auto_mem_in_ar_valid; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_data = _GEN_11 ? _GEN_13 : 32'h0; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_extra = auto_mem_in_ar_valid ? auto_mem_in_ar_bits_id : auto_mem_in_aw_bits_id; // @[Decoupled.scala 289:21]
  assign Queue_io_deq_ready = _T_223_bits_read ? auto_mem_in_r_ready : auto_mem_in_b_ready; // @[Decoupled.scala 311:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ctrlReg = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  maskReg = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      ctrlReg <= 32'h0;
    end else if (_T_125) begin
      ctrlReg <= auto_mem_in_w_bits_data;
    end
    if (reset) begin
      maskReg <= 32'h0;
    end else if (_T_102) begin
      maskReg <= auto_mem_in_w_bits_data;
    end
  end
endmodule
module AXI4StreamMux_2(
  input         clock,
  input         reset,
  output        auto_register_in_aw_ready,
  input         auto_register_in_aw_valid,
  input         auto_register_in_aw_bits_id,
  input  [29:0] auto_register_in_aw_bits_addr,
  output        auto_register_in_w_ready,
  input         auto_register_in_w_valid,
  input  [31:0] auto_register_in_w_bits_data,
  input  [3:0]  auto_register_in_w_bits_strb,
  input         auto_register_in_b_ready,
  output        auto_register_in_b_valid,
  output        auto_register_in_b_bits_id,
  output        auto_register_in_ar_ready,
  input         auto_register_in_ar_valid,
  input         auto_register_in_ar_bits_id,
  input  [29:0] auto_register_in_ar_bits_addr,
  input  [2:0]  auto_register_in_ar_bits_size,
  input         auto_register_in_r_ready,
  output        auto_register_in_r_valid,
  output        auto_register_in_r_bits_id,
  output [31:0] auto_register_in_r_bits_data,
  output        auto_stream_in_2_ready,
  input         auto_stream_in_2_valid,
  input  [31:0] auto_stream_in_2_bits_data,
  input         auto_stream_in_2_bits_last,
  output        auto_stream_in_1_ready,
  input         auto_stream_in_1_valid,
  input  [31:0] auto_stream_in_1_bits_data,
  input         auto_stream_in_1_bits_last,
  output        auto_stream_in_0_ready,
  input         auto_stream_in_0_valid,
  input  [31:0] auto_stream_in_0_bits_data,
  input         auto_stream_in_0_bits_last,
  input         auto_stream_out_0_ready,
  output        auto_stream_out_0_valid,
  output [31:0] auto_stream_out_0_bits_data,
  output        auto_stream_out_0_bits_last
);
  wire  Queue_clock; // @[Decoupled.scala 287:21]
  wire  Queue_reset; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_read; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_enq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_extra; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_read; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_deq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_extra; // @[Decoupled.scala 287:21]
  reg [2:0] sels_0; // @[Mux.scala 32:23]
  reg [31:0] _RAND_0;
  reg [2:0] sels_1; // @[Mux.scala 32:23]
  reg [31:0] _RAND_1;
  wire  _T_3; // @[Mux.scala 45:28]
  wire  _GEN_7; // @[Mux.scala 45:41]
  wire  _GEN_8; // @[Mux.scala 45:41]
  wire  _T_4; // @[Mux.scala 45:28]
  wire  _GEN_12; // @[Mux.scala 45:41]
  wire [31:0] _GEN_15; // @[Mux.scala 45:41]
  wire  _GEN_16; // @[Mux.scala 45:41]
  wire  _GEN_17; // @[Mux.scala 45:41]
  wire  _T_5; // @[Mux.scala 45:28]
  wire  _GEN_21; // @[Mux.scala 45:41]
  wire [31:0] _GEN_24; // @[Mux.scala 45:41]
  wire  _GEN_25; // @[Mux.scala 45:41]
  wire  _GEN_26; // @[Mux.scala 45:41]
  wire  _T_6; // @[Mux.scala 45:28]
  wire  _GEN_30; // @[Mux.scala 45:41]
  wire [31:0] _GEN_33; // @[Mux.scala 45:41]
  wire  _GEN_34; // @[Mux.scala 45:41]
  wire  _T_7; // @[Mux.scala 45:28]
  wire  _T_8; // @[Mux.scala 40:46]
  wire [2:0] _T_10; // @[Mux.scala 41:29]
  wire  _T_11; // @[Mux.scala 45:28]
  wire  _T_12; // @[Mux.scala 45:28]
  wire  _T_13; // @[Mux.scala 45:28]
  wire  _T_17; // @[RegisterRouter.scala 40:39]
  wire  _T_18; // @[RegisterRouter.scala 40:26]
  wire  _T_19; // @[RegisterRouter.scala 42:29]
  wire  _T_62_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 290:17]
  wire [29:0] _T_26; // @[RegisterRouter.scala 48:19]
  wire [1:0] _T_66; // @[RegisterRouter.scala 59:16]
  wire  _T_68; // @[RegisterRouter.scala 59:16]
  wire  _T_20; // @[RegisterRouter.scala 42:26]
  wire [1:0] _T_29; // @[OneHot.scala 65:12]
  wire [1:0] _T_31; // @[Misc.scala 200:81]
  wire  _T_32; // @[Misc.scala 204:21]
  wire  _T_35; // @[Misc.scala 209:20]
  wire  _T_37; // @[Misc.scala 213:38]
  wire  _T_38; // @[Misc.scala 213:29]
  wire  _T_40; // @[Misc.scala 213:38]
  wire  _T_41; // @[Misc.scala 213:29]
  wire  _T_44; // @[Misc.scala 209:20]
  wire  _T_45; // @[Misc.scala 212:27]
  wire  _T_46; // @[Misc.scala 213:38]
  wire  _T_47; // @[Misc.scala 213:29]
  wire  _T_48; // @[Misc.scala 212:27]
  wire  _T_49; // @[Misc.scala 213:38]
  wire  _T_50; // @[Misc.scala 213:29]
  wire  _T_51; // @[Misc.scala 212:27]
  wire  _T_52; // @[Misc.scala 213:38]
  wire  _T_53; // @[Misc.scala 213:29]
  wire  _T_54; // @[Misc.scala 212:27]
  wire  _T_55; // @[Misc.scala 213:38]
  wire  _T_56; // @[Misc.scala 213:29]
  wire [3:0] _T_59; // @[Cat.scala 29:58]
  wire [3:0] _T_61; // @[RegisterRouter.scala 54:25]
  wire [7:0] _T_80; // @[Bitwise.scala 72:12]
  wire [7:0] _T_82; // @[Bitwise.scala 72:12]
  wire [7:0] _T_84; // @[Bitwise.scala 72:12]
  wire [7:0] _T_86; // @[Bitwise.scala 72:12]
  wire [31:0] _T_89; // @[Cat.scala 29:58]
  wire  _T_108; // @[RegisterRouter.scala 59:16]
  wire  _T_161; // @[RegisterRouter.scala 59:16]
  wire [1:0] _T_155; // @[OneHot.scala 58:35]
  wire  _T_178; // @[RegisterRouter.scala 59:16]
  wire  _T_185; // @[RegisterRouter.scala 59:16]
  wire  _T_186; // @[RegisterRouter.scala 59:16]
  wire  _T_115; // @[RegisterRouter.scala 59:16]
  wire  _T_180; // @[RegisterRouter.scala 59:16]
  wire  _T_181; // @[RegisterRouter.scala 59:16]
  wire  _T_138; // @[RegisterRouter.scala 59:16]
  wire  _GEN_101; // @[MuxLiteral.scala 48:10]
  wire [2:0] _GEN_103; // @[MuxLiteral.scala 48:10]
  wire [2:0] _T_235; // @[RegisterRouter.scala 59:16]
  wire  _T_236_bits_read; // @[Decoupled.scala 308:19 Decoupled.scala 309:14]
  wire  _T_236_valid; // @[Decoupled.scala 308:19 Decoupled.scala 310:15]
  wire  _T_239; // @[RegisterRouter.scala 65:29]
  Queue Queue ( // @[Decoupled.scala 287:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_read(Queue_io_enq_bits_read),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_extra(Queue_io_enq_bits_extra),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_read(Queue_io_deq_bits_read),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_extra(Queue_io_deq_bits_extra)
  );
  assign _T_3 = sels_0 == 3'h0; // @[Mux.scala 45:28]
  assign _GEN_7 = _T_3 & auto_stream_in_0_valid; // @[Mux.scala 45:41]
  assign _GEN_8 = _T_3 & auto_stream_out_0_ready; // @[Mux.scala 45:41]
  assign _T_4 = sels_0 == 3'h1; // @[Mux.scala 45:28]
  assign _GEN_12 = _T_4 ? auto_stream_in_1_bits_last : auto_stream_in_0_bits_last; // @[Mux.scala 45:41]
  assign _GEN_15 = _T_4 ? auto_stream_in_1_bits_data : auto_stream_in_0_bits_data; // @[Mux.scala 45:41]
  assign _GEN_16 = _T_4 ? auto_stream_in_1_valid : _GEN_7; // @[Mux.scala 45:41]
  assign _GEN_17 = _T_4 & auto_stream_out_0_ready; // @[Mux.scala 45:41]
  assign _T_5 = sels_0 == 3'h2; // @[Mux.scala 45:28]
  assign _GEN_21 = _T_5 ? auto_stream_in_2_bits_last : _GEN_12; // @[Mux.scala 45:41]
  assign _GEN_24 = _T_5 ? auto_stream_in_2_bits_data : _GEN_15; // @[Mux.scala 45:41]
  assign _GEN_25 = _T_5 ? auto_stream_in_2_valid : _GEN_16; // @[Mux.scala 45:41]
  assign _GEN_26 = _T_5 & auto_stream_out_0_ready; // @[Mux.scala 45:41]
  assign _T_6 = sels_0 == 3'h3; // @[Mux.scala 45:28]
  assign _GEN_30 = _T_6 ? 1'h0 : _GEN_21; // @[Mux.scala 45:41]
  assign _GEN_33 = _T_6 ? 32'hffffffff : _GEN_24; // @[Mux.scala 45:41]
  assign _GEN_34 = _T_6 | _GEN_25; // @[Mux.scala 45:41]
  assign _T_7 = sels_0 == 3'h4; // @[Mux.scala 45:28]
  assign _T_8 = sels_0 == sels_1; // @[Mux.scala 40:46]
  assign _T_10 = _T_8 ? 3'h5 : sels_1; // @[Mux.scala 41:29]
  assign _T_11 = _T_10 == 3'h0; // @[Mux.scala 45:28]
  assign _T_12 = _T_10 == 3'h1; // @[Mux.scala 45:28]
  assign _T_13 = _T_10 == 3'h2; // @[Mux.scala 45:28]
  assign _T_17 = auto_register_in_aw_valid & auto_register_in_w_valid; // @[RegisterRouter.scala 40:39]
  assign _T_18 = auto_register_in_ar_valid | _T_17; // @[RegisterRouter.scala 40:26]
  assign _T_19 = ~auto_register_in_ar_valid; // @[RegisterRouter.scala 42:29]
  assign _T_62_ready = Queue_io_enq_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 290:17]
  assign _T_26 = auto_register_in_ar_valid ? auto_register_in_ar_bits_addr : auto_register_in_aw_bits_addr; // @[RegisterRouter.scala 48:19]
  assign _T_66 = _T_26[3:2] & 2'h2; // @[RegisterRouter.scala 59:16]
  assign _T_68 = _T_66 == 2'h0; // @[RegisterRouter.scala 59:16]
  assign _T_20 = _T_62_ready & _T_19; // @[RegisterRouter.scala 42:26]
  assign _T_29 = 2'h1 << auto_register_in_ar_bits_size[0]; // @[OneHot.scala 65:12]
  assign _T_31 = _T_29 | 2'h1; // @[Misc.scala 200:81]
  assign _T_32 = auto_register_in_ar_bits_size >= 3'h2; // @[Misc.scala 204:21]
  assign _T_35 = ~auto_register_in_ar_bits_addr[1]; // @[Misc.scala 209:20]
  assign _T_37 = _T_31[1] & _T_35; // @[Misc.scala 213:38]
  assign _T_38 = _T_32 | _T_37; // @[Misc.scala 213:29]
  assign _T_40 = _T_31[1] & auto_register_in_ar_bits_addr[1]; // @[Misc.scala 213:38]
  assign _T_41 = _T_32 | _T_40; // @[Misc.scala 213:29]
  assign _T_44 = ~auto_register_in_ar_bits_addr[0]; // @[Misc.scala 209:20]
  assign _T_45 = _T_35 & _T_44; // @[Misc.scala 212:27]
  assign _T_46 = _T_31[0] & _T_45; // @[Misc.scala 213:38]
  assign _T_47 = _T_38 | _T_46; // @[Misc.scala 213:29]
  assign _T_48 = _T_35 & auto_register_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  assign _T_49 = _T_31[0] & _T_48; // @[Misc.scala 213:38]
  assign _T_50 = _T_38 | _T_49; // @[Misc.scala 213:29]
  assign _T_51 = auto_register_in_ar_bits_addr[1] & _T_44; // @[Misc.scala 212:27]
  assign _T_52 = _T_31[0] & _T_51; // @[Misc.scala 213:38]
  assign _T_53 = _T_41 | _T_52; // @[Misc.scala 213:29]
  assign _T_54 = auto_register_in_ar_bits_addr[1] & auto_register_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  assign _T_55 = _T_31[0] & _T_54; // @[Misc.scala 213:38]
  assign _T_56 = _T_41 | _T_55; // @[Misc.scala 213:29]
  assign _T_59 = {_T_56,_T_53,_T_50,_T_47}; // @[Cat.scala 29:58]
  assign _T_61 = auto_register_in_ar_valid ? _T_59 : auto_register_in_w_bits_strb; // @[RegisterRouter.scala 54:25]
  assign _T_80 = _T_61[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_82 = _T_61[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_84 = _T_61[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_86 = _T_61[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_89 = {_T_86,_T_84,_T_82,_T_80}; // @[Cat.scala 29:58]
  assign _T_108 = _T_89[2:0] == 3'h7; // @[RegisterRouter.scala 59:16]
  assign _T_161 = _T_18 & _T_62_ready; // @[RegisterRouter.scala 59:16]
  assign _T_155 = 2'h1 << _T_26[2]; // @[OneHot.scala 58:35]
  assign _T_178 = _T_161 & _T_19; // @[RegisterRouter.scala 59:16]
  assign _T_185 = _T_178 & _T_155[1]; // @[RegisterRouter.scala 59:16]
  assign _T_186 = _T_185 & _T_68; // @[RegisterRouter.scala 59:16]
  assign _T_115 = _T_186 & _T_108; // @[RegisterRouter.scala 59:16]
  assign _T_180 = _T_178 & _T_155[0]; // @[RegisterRouter.scala 59:16]
  assign _T_181 = _T_180 & _T_68; // @[RegisterRouter.scala 59:16]
  assign _T_138 = _T_181 & _T_108; // @[RegisterRouter.scala 59:16]
  assign _GEN_101 = _T_26[2] ? _T_68 : _T_68; // @[MuxLiteral.scala 48:10]
  assign _GEN_103 = _T_26[2] ? sels_1 : sels_0; // @[MuxLiteral.scala 48:10]
  assign _T_235 = _GEN_101 ? _GEN_103 : 3'h0; // @[RegisterRouter.scala 59:16]
  assign _T_236_bits_read = Queue_io_deq_bits_read; // @[Decoupled.scala 308:19 Decoupled.scala 309:14]
  assign _T_236_valid = Queue_io_deq_valid; // @[Decoupled.scala 308:19 Decoupled.scala 310:15]
  assign _T_239 = ~_T_236_bits_read; // @[RegisterRouter.scala 65:29]
  assign auto_register_in_aw_ready = _T_20 & auto_register_in_w_valid; // @[LazyModule.scala 173:31]
  assign auto_register_in_w_ready = _T_20 & auto_register_in_aw_valid; // @[LazyModule.scala 173:31]
  assign auto_register_in_b_valid = _T_236_valid & _T_239; // @[LazyModule.scala 173:31]
  assign auto_register_in_b_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_register_in_ar_ready = Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_register_in_r_valid = _T_236_valid & _T_236_bits_read; // @[LazyModule.scala 173:31]
  assign auto_register_in_r_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_register_in_r_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 173:31]
  assign auto_stream_in_2_ready = _T_13 | _GEN_26; // @[LazyModule.scala 173:31]
  assign auto_stream_in_1_ready = _T_12 | _GEN_17; // @[LazyModule.scala 173:31]
  assign auto_stream_in_0_ready = _T_11 | _GEN_8; // @[LazyModule.scala 173:31]
  assign auto_stream_out_0_valid = _T_7 | _GEN_34; // @[LazyModule.scala 173:49]
  assign auto_stream_out_0_bits_data = _T_7 ? 32'h0 : _GEN_33; // @[LazyModule.scala 173:49]
  assign auto_stream_out_0_bits_last = _T_7 ? 1'h0 : _GEN_30; // @[LazyModule.scala 173:49]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_register_in_ar_valid | _T_17; // @[Decoupled.scala 288:22]
  assign Queue_io_enq_bits_read = auto_register_in_ar_valid; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_data = {{29'd0}, _T_235}; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_extra = auto_register_in_ar_valid ? auto_register_in_ar_bits_id : auto_register_in_aw_bits_id; // @[Decoupled.scala 289:21]
  assign Queue_io_deq_ready = _T_236_bits_read ? auto_register_in_r_ready : auto_register_in_b_ready; // @[Decoupled.scala 311:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  sels_0 = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  sels_1 = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      sels_0 <= 3'h5;
    end else if (_T_138) begin
      sels_0 <= auto_register_in_w_bits_data[2:0];
    end
    if (reset) begin
      sels_1 <= 3'h5;
    end else if (_T_115) begin
      sels_1 <= auto_register_in_w_bits_data[2:0];
    end
  end
endmodule
module SDFStageRadix22(
  input         clock,
  input         reset,
  input  [15:0] io_in_real,
  input  [15:0] io_in_imag,
  output [15:0] io_out_real,
  output [15:0] io_out_imag,
  input  [5:0]  io_cntr,
  input         io_en
);
  wire  load_input; // @[SDFChainRadix22.scala 426:66]
  reg [15:0] shift_out_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_0;
  wire [16:0] butt_outputs_1_real; // @[FixedPointTypeClass.scala 33:22]
  wire [17:0] _T_140; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_142; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_145; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] butterfly_outputs_1_real; // @[FixedPointTypeClass.scala 176:41]
  reg [15:0] shift_out_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1;
  wire [16:0] butt_outputs_1_imag; // @[FixedPointTypeClass.scala 33:22]
  wire [17:0] _T_147; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_149; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_152; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] butterfly_outputs_1_imag; // @[FixedPointTypeClass.scala 176:41]
  reg [15:0] _T_21_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2;
  reg [15:0] _T_21_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3;
  reg [15:0] _T_24_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4;
  reg [15:0] _T_24_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5;
  reg [15:0] _T_27_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6;
  reg [15:0] _T_27_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7;
  reg [15:0] _T_30_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8;
  reg [15:0] _T_30_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9;
  reg [15:0] _T_33_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10;
  reg [15:0] _T_33_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11;
  reg [15:0] _T_36_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12;
  reg [15:0] _T_36_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_13;
  reg [15:0] _T_39_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_14;
  reg [15:0] _T_39_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_15;
  reg [15:0] _T_42_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_16;
  reg [15:0] _T_42_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_17;
  reg [15:0] _T_45_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_18;
  reg [15:0] _T_45_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_19;
  reg [15:0] _T_48_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_20;
  reg [15:0] _T_48_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_21;
  reg [15:0] _T_51_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_22;
  reg [15:0] _T_51_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_23;
  reg [15:0] _T_54_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_24;
  reg [15:0] _T_54_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_25;
  reg [15:0] _T_57_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_26;
  reg [15:0] _T_57_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_27;
  reg [15:0] _T_60_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_28;
  reg [15:0] _T_60_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_29;
  reg [15:0] _T_63_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_30;
  reg [15:0] _T_63_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_31;
  reg [15:0] _T_66_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_32;
  reg [15:0] _T_66_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_33;
  reg [15:0] _T_69_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_34;
  reg [15:0] _T_69_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_35;
  reg [15:0] _T_72_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_36;
  reg [15:0] _T_72_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_37;
  reg [15:0] _T_75_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_38;
  reg [15:0] _T_75_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_39;
  reg [15:0] _T_78_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_40;
  reg [15:0] _T_78_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_41;
  reg [15:0] _T_81_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_42;
  reg [15:0] _T_81_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_43;
  reg [15:0] _T_84_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_44;
  reg [15:0] _T_84_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_45;
  reg [15:0] _T_87_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_46;
  reg [15:0] _T_87_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_47;
  reg [15:0] _T_90_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_48;
  reg [15:0] _T_90_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_49;
  reg [15:0] _T_93_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_50;
  reg [15:0] _T_93_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_51;
  reg [15:0] _T_96_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_52;
  reg [15:0] _T_96_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_53;
  reg [15:0] _T_99_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_54;
  reg [15:0] _T_99_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_55;
  reg [15:0] _T_102_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_56;
  reg [15:0] _T_102_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_57;
  reg [15:0] _T_105_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_58;
  reg [15:0] _T_105_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_59;
  reg [15:0] _T_108_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_60;
  reg [15:0] _T_108_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_61;
  reg [15:0] _T_111_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_62;
  reg [15:0] _T_111_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_63;
  wire [16:0] butt_outputs_0_real; // @[FixedPointTypeClass.scala 24:22]
  wire [16:0] butt_outputs_0_imag; // @[FixedPointTypeClass.scala 24:22]
  wire [17:0] _T_123; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_125; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_128; // @[FixedPointTypeClass.scala 20:58]
  wire [17:0] _T_130; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_132; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_135; // @[FixedPointTypeClass.scala 20:58]
  reg [15:0] feedback_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_64;
  reg [15:0] feedback_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_65;
  reg [15:0] butt_out_0_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_66;
  reg [15:0] butt_out_0_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_67;
  reg  load_output; // @[Reg.scala 27:20]
  reg [31:0] _RAND_68;
  assign load_input = io_cntr < 6'h20; // @[SDFChainRadix22.scala 426:66]
  assign butt_outputs_1_real = $signed(shift_out_real) - $signed(io_in_real); // @[FixedPointTypeClass.scala 33:22]
  assign _T_140 = {$signed(butt_outputs_1_real), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign _T_142 = _T_140[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign _T_145 = $signed(_T_142) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign butterfly_outputs_1_real = _T_145[16:1]; // @[FixedPointTypeClass.scala 176:41]
  assign butt_outputs_1_imag = $signed(shift_out_imag) - $signed(io_in_imag); // @[FixedPointTypeClass.scala 33:22]
  assign _T_147 = {$signed(butt_outputs_1_imag), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign _T_149 = _T_147[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign _T_152 = $signed(_T_149) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign butterfly_outputs_1_imag = _T_152[16:1]; // @[FixedPointTypeClass.scala 176:41]
  assign butt_outputs_0_real = $signed(shift_out_real) + $signed(io_in_real); // @[FixedPointTypeClass.scala 24:22]
  assign butt_outputs_0_imag = $signed(shift_out_imag) + $signed(io_in_imag); // @[FixedPointTypeClass.scala 24:22]
  assign _T_123 = {$signed(butt_outputs_0_real), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign _T_125 = _T_123[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign _T_128 = $signed(_T_125) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign _T_130 = {$signed(butt_outputs_0_imag), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign _T_132 = _T_130[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign _T_135 = $signed(_T_132) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign io_out_real = load_output ? $signed(feedback_real) : $signed(butt_out_0_real); // @[SDFChainRadix22.scala 422:10]
  assign io_out_imag = load_output ? $signed(feedback_imag) : $signed(butt_out_0_imag); // @[SDFChainRadix22.scala 422:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  shift_out_real = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  shift_out_imag = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_21_real = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_21_imag = _RAND_3[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_24_real = _RAND_4[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_24_imag = _RAND_5[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_27_real = _RAND_6[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_27_imag = _RAND_7[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_30_real = _RAND_8[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_30_imag = _RAND_9[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_33_real = _RAND_10[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_33_imag = _RAND_11[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_36_real = _RAND_12[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_36_imag = _RAND_13[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_39_real = _RAND_14[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_39_imag = _RAND_15[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_42_real = _RAND_16[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_42_imag = _RAND_17[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_45_real = _RAND_18[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_45_imag = _RAND_19[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_48_real = _RAND_20[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_48_imag = _RAND_21[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_51_real = _RAND_22[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_51_imag = _RAND_23[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_54_real = _RAND_24[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_54_imag = _RAND_25[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_57_real = _RAND_26[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T_57_imag = _RAND_27[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_60_real = _RAND_28[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_60_imag = _RAND_29[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_63_real = _RAND_30[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T_63_imag = _RAND_31[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _T_66_real = _RAND_32[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _T_66_imag = _RAND_33[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _T_69_real = _RAND_34[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _T_69_imag = _RAND_35[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _T_72_real = _RAND_36[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _T_72_imag = _RAND_37[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _T_75_real = _RAND_38[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _T_75_imag = _RAND_39[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _T_78_real = _RAND_40[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  _T_78_imag = _RAND_41[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  _T_81_real = _RAND_42[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  _T_81_imag = _RAND_43[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  _T_84_real = _RAND_44[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  _T_84_imag = _RAND_45[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  _T_87_real = _RAND_46[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  _T_87_imag = _RAND_47[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  _T_90_real = _RAND_48[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  _T_90_imag = _RAND_49[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  _T_93_real = _RAND_50[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  _T_93_imag = _RAND_51[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  _T_96_real = _RAND_52[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  _T_96_imag = _RAND_53[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  _T_99_real = _RAND_54[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  _T_99_imag = _RAND_55[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  _T_102_real = _RAND_56[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  _T_102_imag = _RAND_57[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  _T_105_real = _RAND_58[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  _T_105_imag = _RAND_59[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  _T_108_real = _RAND_60[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  _T_108_imag = _RAND_61[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  _T_111_real = _RAND_62[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  _T_111_imag = _RAND_63[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  feedback_real = _RAND_64[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  feedback_imag = _RAND_65[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  butt_out_0_real = _RAND_66[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  butt_out_0_imag = _RAND_67[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  load_output = _RAND_68[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (io_en) begin
      shift_out_real <= _T_111_real;
    end
    if (io_en) begin
      shift_out_imag <= _T_111_imag;
    end
    if (io_en) begin
      if (load_input) begin
        _T_21_real <= io_in_real;
      end else begin
        _T_21_real <= butterfly_outputs_1_real;
      end
    end
    if (io_en) begin
      if (load_input) begin
        _T_21_imag <= io_in_imag;
      end else begin
        _T_21_imag <= butterfly_outputs_1_imag;
      end
    end
    if (io_en) begin
      _T_24_real <= _T_21_real;
    end
    if (io_en) begin
      _T_24_imag <= _T_21_imag;
    end
    if (io_en) begin
      _T_27_real <= _T_24_real;
    end
    if (io_en) begin
      _T_27_imag <= _T_24_imag;
    end
    if (io_en) begin
      _T_30_real <= _T_27_real;
    end
    if (io_en) begin
      _T_30_imag <= _T_27_imag;
    end
    if (io_en) begin
      _T_33_real <= _T_30_real;
    end
    if (io_en) begin
      _T_33_imag <= _T_30_imag;
    end
    if (io_en) begin
      _T_36_real <= _T_33_real;
    end
    if (io_en) begin
      _T_36_imag <= _T_33_imag;
    end
    if (io_en) begin
      _T_39_real <= _T_36_real;
    end
    if (io_en) begin
      _T_39_imag <= _T_36_imag;
    end
    if (io_en) begin
      _T_42_real <= _T_39_real;
    end
    if (io_en) begin
      _T_42_imag <= _T_39_imag;
    end
    if (io_en) begin
      _T_45_real <= _T_42_real;
    end
    if (io_en) begin
      _T_45_imag <= _T_42_imag;
    end
    if (io_en) begin
      _T_48_real <= _T_45_real;
    end
    if (io_en) begin
      _T_48_imag <= _T_45_imag;
    end
    if (io_en) begin
      _T_51_real <= _T_48_real;
    end
    if (io_en) begin
      _T_51_imag <= _T_48_imag;
    end
    if (io_en) begin
      _T_54_real <= _T_51_real;
    end
    if (io_en) begin
      _T_54_imag <= _T_51_imag;
    end
    if (io_en) begin
      _T_57_real <= _T_54_real;
    end
    if (io_en) begin
      _T_57_imag <= _T_54_imag;
    end
    if (io_en) begin
      _T_60_real <= _T_57_real;
    end
    if (io_en) begin
      _T_60_imag <= _T_57_imag;
    end
    if (io_en) begin
      _T_63_real <= _T_60_real;
    end
    if (io_en) begin
      _T_63_imag <= _T_60_imag;
    end
    if (io_en) begin
      _T_66_real <= _T_63_real;
    end
    if (io_en) begin
      _T_66_imag <= _T_63_imag;
    end
    if (io_en) begin
      _T_69_real <= _T_66_real;
    end
    if (io_en) begin
      _T_69_imag <= _T_66_imag;
    end
    if (io_en) begin
      _T_72_real <= _T_69_real;
    end
    if (io_en) begin
      _T_72_imag <= _T_69_imag;
    end
    if (io_en) begin
      _T_75_real <= _T_72_real;
    end
    if (io_en) begin
      _T_75_imag <= _T_72_imag;
    end
    if (io_en) begin
      _T_78_real <= _T_75_real;
    end
    if (io_en) begin
      _T_78_imag <= _T_75_imag;
    end
    if (io_en) begin
      _T_81_real <= _T_78_real;
    end
    if (io_en) begin
      _T_81_imag <= _T_78_imag;
    end
    if (io_en) begin
      _T_84_real <= _T_81_real;
    end
    if (io_en) begin
      _T_84_imag <= _T_81_imag;
    end
    if (io_en) begin
      _T_87_real <= _T_84_real;
    end
    if (io_en) begin
      _T_87_imag <= _T_84_imag;
    end
    if (io_en) begin
      _T_90_real <= _T_87_real;
    end
    if (io_en) begin
      _T_90_imag <= _T_87_imag;
    end
    if (io_en) begin
      _T_93_real <= _T_90_real;
    end
    if (io_en) begin
      _T_93_imag <= _T_90_imag;
    end
    if (io_en) begin
      _T_96_real <= _T_93_real;
    end
    if (io_en) begin
      _T_96_imag <= _T_93_imag;
    end
    if (io_en) begin
      _T_99_real <= _T_96_real;
    end
    if (io_en) begin
      _T_99_imag <= _T_96_imag;
    end
    if (io_en) begin
      _T_102_real <= _T_99_real;
    end
    if (io_en) begin
      _T_102_imag <= _T_99_imag;
    end
    if (io_en) begin
      _T_105_real <= _T_102_real;
    end
    if (io_en) begin
      _T_105_imag <= _T_102_imag;
    end
    if (io_en) begin
      _T_108_real <= _T_105_real;
    end
    if (io_en) begin
      _T_108_imag <= _T_105_imag;
    end
    if (io_en) begin
      _T_111_real <= _T_108_real;
    end
    if (io_en) begin
      _T_111_imag <= _T_108_imag;
    end
    feedback_real <= shift_out_real;
    feedback_imag <= shift_out_imag;
    butt_out_0_real <= _T_128[16:1];
    butt_out_0_imag <= _T_135[16:1];
    if (reset) begin
      load_output <= 1'h0;
    end else begin
      load_output <= load_input;
    end
  end
endmodule
module SDFStageRadix22_1(
  input         clock,
  input         reset,
  input  [15:0] io_in_real,
  input  [15:0] io_in_imag,
  output [15:0] io_out_real,
  output [15:0] io_out_imag,
  input  [5:0]  io_cntr,
  input         io_en
);
  wire  load_input; // @[SDFChainRadix22.scala 426:66]
  reg [15:0] shift_out_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_0;
  wire [16:0] butt_outputs_1_real; // @[FixedPointTypeClass.scala 33:22]
  wire [17:0] _T_92; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_94; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_97; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] butterfly_outputs_1_real; // @[FixedPointTypeClass.scala 176:41]
  reg [15:0] shift_out_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1;
  wire [16:0] butt_outputs_1_imag; // @[FixedPointTypeClass.scala 33:22]
  wire [17:0] _T_99; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_101; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_104; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] butterfly_outputs_1_imag; // @[FixedPointTypeClass.scala 176:41]
  reg [15:0] _T_21_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2;
  reg [15:0] _T_21_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3;
  reg [15:0] _T_24_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4;
  reg [15:0] _T_24_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5;
  reg [15:0] _T_27_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6;
  reg [15:0] _T_27_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7;
  reg [15:0] _T_30_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8;
  reg [15:0] _T_30_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9;
  reg [15:0] _T_33_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10;
  reg [15:0] _T_33_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11;
  reg [15:0] _T_36_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12;
  reg [15:0] _T_36_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_13;
  reg [15:0] _T_39_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_14;
  reg [15:0] _T_39_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_15;
  reg [15:0] _T_42_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_16;
  reg [15:0] _T_42_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_17;
  reg [15:0] _T_45_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_18;
  reg [15:0] _T_45_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_19;
  reg [15:0] _T_48_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_20;
  reg [15:0] _T_48_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_21;
  reg [15:0] _T_51_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_22;
  reg [15:0] _T_51_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_23;
  reg [15:0] _T_54_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_24;
  reg [15:0] _T_54_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_25;
  reg [15:0] _T_57_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_26;
  reg [15:0] _T_57_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_27;
  reg [15:0] _T_60_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_28;
  reg [15:0] _T_60_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_29;
  reg [15:0] _T_63_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_30;
  reg [15:0] _T_63_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_31;
  wire [16:0] butt_outputs_0_real; // @[FixedPointTypeClass.scala 24:22]
  wire [16:0] butt_outputs_0_imag; // @[FixedPointTypeClass.scala 24:22]
  wire [17:0] _T_75; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_77; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_80; // @[FixedPointTypeClass.scala 20:58]
  wire [17:0] _T_82; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_84; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_87; // @[FixedPointTypeClass.scala 20:58]
  reg [15:0] feedback_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_32;
  reg [15:0] feedback_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_33;
  reg [15:0] butt_out_0_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_34;
  reg [15:0] butt_out_0_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_35;
  reg  load_output; // @[Reg.scala 27:20]
  reg [31:0] _RAND_36;
  assign load_input = io_cntr < 6'h10; // @[SDFChainRadix22.scala 426:66]
  assign butt_outputs_1_real = $signed(shift_out_real) - $signed(io_in_real); // @[FixedPointTypeClass.scala 33:22]
  assign _T_92 = {$signed(butt_outputs_1_real), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign _T_94 = _T_92[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign _T_97 = $signed(_T_94) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign butterfly_outputs_1_real = _T_97[16:1]; // @[FixedPointTypeClass.scala 176:41]
  assign butt_outputs_1_imag = $signed(shift_out_imag) - $signed(io_in_imag); // @[FixedPointTypeClass.scala 33:22]
  assign _T_99 = {$signed(butt_outputs_1_imag), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign _T_101 = _T_99[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign _T_104 = $signed(_T_101) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign butterfly_outputs_1_imag = _T_104[16:1]; // @[FixedPointTypeClass.scala 176:41]
  assign butt_outputs_0_real = $signed(shift_out_real) + $signed(io_in_real); // @[FixedPointTypeClass.scala 24:22]
  assign butt_outputs_0_imag = $signed(shift_out_imag) + $signed(io_in_imag); // @[FixedPointTypeClass.scala 24:22]
  assign _T_75 = {$signed(butt_outputs_0_real), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign _T_77 = _T_75[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign _T_80 = $signed(_T_77) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign _T_82 = {$signed(butt_outputs_0_imag), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign _T_84 = _T_82[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign _T_87 = $signed(_T_84) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign io_out_real = load_output ? $signed(feedback_real) : $signed(butt_out_0_real); // @[SDFChainRadix22.scala 422:10]
  assign io_out_imag = load_output ? $signed(feedback_imag) : $signed(butt_out_0_imag); // @[SDFChainRadix22.scala 422:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  shift_out_real = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  shift_out_imag = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_21_real = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_21_imag = _RAND_3[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_24_real = _RAND_4[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_24_imag = _RAND_5[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_27_real = _RAND_6[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_27_imag = _RAND_7[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_30_real = _RAND_8[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_30_imag = _RAND_9[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_33_real = _RAND_10[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_33_imag = _RAND_11[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_36_real = _RAND_12[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_36_imag = _RAND_13[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_39_real = _RAND_14[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_39_imag = _RAND_15[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_42_real = _RAND_16[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_42_imag = _RAND_17[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_45_real = _RAND_18[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_45_imag = _RAND_19[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_48_real = _RAND_20[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_48_imag = _RAND_21[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_51_real = _RAND_22[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_51_imag = _RAND_23[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_54_real = _RAND_24[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_54_imag = _RAND_25[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_57_real = _RAND_26[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T_57_imag = _RAND_27[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_60_real = _RAND_28[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_60_imag = _RAND_29[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_63_real = _RAND_30[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T_63_imag = _RAND_31[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  feedback_real = _RAND_32[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  feedback_imag = _RAND_33[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  butt_out_0_real = _RAND_34[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  butt_out_0_imag = _RAND_35[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  load_output = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (io_en) begin
      shift_out_real <= _T_63_real;
    end
    if (io_en) begin
      shift_out_imag <= _T_63_imag;
    end
    if (io_en) begin
      if (load_input) begin
        _T_21_real <= io_in_real;
      end else begin
        _T_21_real <= butterfly_outputs_1_real;
      end
    end
    if (io_en) begin
      if (load_input) begin
        _T_21_imag <= io_in_imag;
      end else begin
        _T_21_imag <= butterfly_outputs_1_imag;
      end
    end
    if (io_en) begin
      _T_24_real <= _T_21_real;
    end
    if (io_en) begin
      _T_24_imag <= _T_21_imag;
    end
    if (io_en) begin
      _T_27_real <= _T_24_real;
    end
    if (io_en) begin
      _T_27_imag <= _T_24_imag;
    end
    if (io_en) begin
      _T_30_real <= _T_27_real;
    end
    if (io_en) begin
      _T_30_imag <= _T_27_imag;
    end
    if (io_en) begin
      _T_33_real <= _T_30_real;
    end
    if (io_en) begin
      _T_33_imag <= _T_30_imag;
    end
    if (io_en) begin
      _T_36_real <= _T_33_real;
    end
    if (io_en) begin
      _T_36_imag <= _T_33_imag;
    end
    if (io_en) begin
      _T_39_real <= _T_36_real;
    end
    if (io_en) begin
      _T_39_imag <= _T_36_imag;
    end
    if (io_en) begin
      _T_42_real <= _T_39_real;
    end
    if (io_en) begin
      _T_42_imag <= _T_39_imag;
    end
    if (io_en) begin
      _T_45_real <= _T_42_real;
    end
    if (io_en) begin
      _T_45_imag <= _T_42_imag;
    end
    if (io_en) begin
      _T_48_real <= _T_45_real;
    end
    if (io_en) begin
      _T_48_imag <= _T_45_imag;
    end
    if (io_en) begin
      _T_51_real <= _T_48_real;
    end
    if (io_en) begin
      _T_51_imag <= _T_48_imag;
    end
    if (io_en) begin
      _T_54_real <= _T_51_real;
    end
    if (io_en) begin
      _T_54_imag <= _T_51_imag;
    end
    if (io_en) begin
      _T_57_real <= _T_54_real;
    end
    if (io_en) begin
      _T_57_imag <= _T_54_imag;
    end
    if (io_en) begin
      _T_60_real <= _T_57_real;
    end
    if (io_en) begin
      _T_60_imag <= _T_57_imag;
    end
    if (io_en) begin
      _T_63_real <= _T_60_real;
    end
    if (io_en) begin
      _T_63_imag <= _T_60_imag;
    end
    feedback_real <= shift_out_real;
    feedback_imag <= shift_out_imag;
    butt_out_0_real <= _T_80[16:1];
    butt_out_0_imag <= _T_87[16:1];
    if (reset) begin
      load_output <= 1'h0;
    end else begin
      load_output <= load_input;
    end
  end
endmodule
module SDFStageRadix22_2(
  input         clock,
  input         reset,
  input  [15:0] io_in_real,
  input  [15:0] io_in_imag,
  output [15:0] io_out_real,
  output [15:0] io_out_imag,
  input  [5:0]  io_cntr,
  input         io_en
);
  wire  load_input; // @[SDFChainRadix22.scala 426:66]
  reg [15:0] shift_out_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_0;
  wire [16:0] butt_outputs_1_real; // @[FixedPointTypeClass.scala 33:22]
  wire [17:0] _T_68; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_70; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_73; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] butterfly_outputs_1_real; // @[FixedPointTypeClass.scala 176:41]
  reg [15:0] shift_out_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1;
  wire [16:0] butt_outputs_1_imag; // @[FixedPointTypeClass.scala 33:22]
  wire [17:0] _T_75; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_77; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_80; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] butterfly_outputs_1_imag; // @[FixedPointTypeClass.scala 176:41]
  reg [15:0] _T_21_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2;
  reg [15:0] _T_21_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3;
  reg [15:0] _T_24_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4;
  reg [15:0] _T_24_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5;
  reg [15:0] _T_27_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6;
  reg [15:0] _T_27_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7;
  reg [15:0] _T_30_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8;
  reg [15:0] _T_30_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9;
  reg [15:0] _T_33_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10;
  reg [15:0] _T_33_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11;
  reg [15:0] _T_36_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12;
  reg [15:0] _T_36_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_13;
  reg [15:0] _T_39_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_14;
  reg [15:0] _T_39_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_15;
  wire [16:0] butt_outputs_0_real; // @[FixedPointTypeClass.scala 24:22]
  wire [16:0] butt_outputs_0_imag; // @[FixedPointTypeClass.scala 24:22]
  wire [17:0] _T_51; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_53; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_56; // @[FixedPointTypeClass.scala 20:58]
  wire [17:0] _T_58; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_60; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_63; // @[FixedPointTypeClass.scala 20:58]
  reg [15:0] feedback_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_16;
  reg [15:0] feedback_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_17;
  reg [15:0] butt_out_0_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_18;
  reg [15:0] butt_out_0_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_19;
  reg  load_output; // @[Reg.scala 27:20]
  reg [31:0] _RAND_20;
  assign load_input = io_cntr < 6'h8; // @[SDFChainRadix22.scala 426:66]
  assign butt_outputs_1_real = $signed(shift_out_real) - $signed(io_in_real); // @[FixedPointTypeClass.scala 33:22]
  assign _T_68 = {$signed(butt_outputs_1_real), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign _T_70 = _T_68[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign _T_73 = $signed(_T_70) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign butterfly_outputs_1_real = _T_73[16:1]; // @[FixedPointTypeClass.scala 176:41]
  assign butt_outputs_1_imag = $signed(shift_out_imag) - $signed(io_in_imag); // @[FixedPointTypeClass.scala 33:22]
  assign _T_75 = {$signed(butt_outputs_1_imag), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign _T_77 = _T_75[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign _T_80 = $signed(_T_77) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign butterfly_outputs_1_imag = _T_80[16:1]; // @[FixedPointTypeClass.scala 176:41]
  assign butt_outputs_0_real = $signed(shift_out_real) + $signed(io_in_real); // @[FixedPointTypeClass.scala 24:22]
  assign butt_outputs_0_imag = $signed(shift_out_imag) + $signed(io_in_imag); // @[FixedPointTypeClass.scala 24:22]
  assign _T_51 = {$signed(butt_outputs_0_real), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign _T_53 = _T_51[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign _T_56 = $signed(_T_53) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign _T_58 = {$signed(butt_outputs_0_imag), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign _T_60 = _T_58[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign _T_63 = $signed(_T_60) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign io_out_real = load_output ? $signed(feedback_real) : $signed(butt_out_0_real); // @[SDFChainRadix22.scala 422:10]
  assign io_out_imag = load_output ? $signed(feedback_imag) : $signed(butt_out_0_imag); // @[SDFChainRadix22.scala 422:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  shift_out_real = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  shift_out_imag = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_21_real = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_21_imag = _RAND_3[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_24_real = _RAND_4[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_24_imag = _RAND_5[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_27_real = _RAND_6[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_27_imag = _RAND_7[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_30_real = _RAND_8[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_30_imag = _RAND_9[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_33_real = _RAND_10[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_33_imag = _RAND_11[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_36_real = _RAND_12[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_36_imag = _RAND_13[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_39_real = _RAND_14[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_39_imag = _RAND_15[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  feedback_real = _RAND_16[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  feedback_imag = _RAND_17[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  butt_out_0_real = _RAND_18[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  butt_out_0_imag = _RAND_19[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  load_output = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (io_en) begin
      shift_out_real <= _T_39_real;
    end
    if (io_en) begin
      shift_out_imag <= _T_39_imag;
    end
    if (io_en) begin
      if (load_input) begin
        _T_21_real <= io_in_real;
      end else begin
        _T_21_real <= butterfly_outputs_1_real;
      end
    end
    if (io_en) begin
      if (load_input) begin
        _T_21_imag <= io_in_imag;
      end else begin
        _T_21_imag <= butterfly_outputs_1_imag;
      end
    end
    if (io_en) begin
      _T_24_real <= _T_21_real;
    end
    if (io_en) begin
      _T_24_imag <= _T_21_imag;
    end
    if (io_en) begin
      _T_27_real <= _T_24_real;
    end
    if (io_en) begin
      _T_27_imag <= _T_24_imag;
    end
    if (io_en) begin
      _T_30_real <= _T_27_real;
    end
    if (io_en) begin
      _T_30_imag <= _T_27_imag;
    end
    if (io_en) begin
      _T_33_real <= _T_30_real;
    end
    if (io_en) begin
      _T_33_imag <= _T_30_imag;
    end
    if (io_en) begin
      _T_36_real <= _T_33_real;
    end
    if (io_en) begin
      _T_36_imag <= _T_33_imag;
    end
    if (io_en) begin
      _T_39_real <= _T_36_real;
    end
    if (io_en) begin
      _T_39_imag <= _T_36_imag;
    end
    feedback_real <= shift_out_real;
    feedback_imag <= shift_out_imag;
    butt_out_0_real <= _T_56[16:1];
    butt_out_0_imag <= _T_63[16:1];
    if (reset) begin
      load_output <= 1'h0;
    end else begin
      load_output <= load_input;
    end
  end
endmodule
module SDFStageRadix22_3(
  input         clock,
  input         reset,
  input  [15:0] io_in_real,
  input  [15:0] io_in_imag,
  output [15:0] io_out_real,
  output [15:0] io_out_imag,
  input  [5:0]  io_cntr,
  input         io_en
);
  wire  load_input; // @[SDFChainRadix22.scala 426:66]
  reg [15:0] shift_out_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_0;
  wire [16:0] butt_outputs_1_real; // @[FixedPointTypeClass.scala 33:22]
  wire [17:0] _T_56; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_58; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_61; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] butterfly_outputs_1_real; // @[FixedPointTypeClass.scala 176:41]
  reg [15:0] shift_out_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1;
  wire [16:0] butt_outputs_1_imag; // @[FixedPointTypeClass.scala 33:22]
  wire [17:0] _T_63; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_65; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_68; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] butterfly_outputs_1_imag; // @[FixedPointTypeClass.scala 176:41]
  reg [15:0] _T_21_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2;
  reg [15:0] _T_21_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3;
  reg [15:0] _T_24_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4;
  reg [15:0] _T_24_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5;
  reg [15:0] _T_27_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6;
  reg [15:0] _T_27_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7;
  wire [16:0] butt_outputs_0_real; // @[FixedPointTypeClass.scala 24:22]
  wire [16:0] butt_outputs_0_imag; // @[FixedPointTypeClass.scala 24:22]
  wire [17:0] _T_39; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_41; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_44; // @[FixedPointTypeClass.scala 20:58]
  wire [17:0] _T_46; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_48; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_51; // @[FixedPointTypeClass.scala 20:58]
  reg [15:0] feedback_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8;
  reg [15:0] feedback_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9;
  reg [15:0] butt_out_0_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10;
  reg [15:0] butt_out_0_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11;
  reg  load_output; // @[Reg.scala 27:20]
  reg [31:0] _RAND_12;
  assign load_input = io_cntr < 6'h4; // @[SDFChainRadix22.scala 426:66]
  assign butt_outputs_1_real = $signed(shift_out_real) - $signed(io_in_real); // @[FixedPointTypeClass.scala 33:22]
  assign _T_56 = {$signed(butt_outputs_1_real), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign _T_58 = _T_56[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign _T_61 = $signed(_T_58) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign butterfly_outputs_1_real = _T_61[16:1]; // @[FixedPointTypeClass.scala 176:41]
  assign butt_outputs_1_imag = $signed(shift_out_imag) - $signed(io_in_imag); // @[FixedPointTypeClass.scala 33:22]
  assign _T_63 = {$signed(butt_outputs_1_imag), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign _T_65 = _T_63[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign _T_68 = $signed(_T_65) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign butterfly_outputs_1_imag = _T_68[16:1]; // @[FixedPointTypeClass.scala 176:41]
  assign butt_outputs_0_real = $signed(shift_out_real) + $signed(io_in_real); // @[FixedPointTypeClass.scala 24:22]
  assign butt_outputs_0_imag = $signed(shift_out_imag) + $signed(io_in_imag); // @[FixedPointTypeClass.scala 24:22]
  assign _T_39 = {$signed(butt_outputs_0_real), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign _T_41 = _T_39[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign _T_44 = $signed(_T_41) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign _T_46 = {$signed(butt_outputs_0_imag), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign _T_48 = _T_46[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign _T_51 = $signed(_T_48) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign io_out_real = load_output ? $signed(feedback_real) : $signed(butt_out_0_real); // @[SDFChainRadix22.scala 422:10]
  assign io_out_imag = load_output ? $signed(feedback_imag) : $signed(butt_out_0_imag); // @[SDFChainRadix22.scala 422:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  shift_out_real = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  shift_out_imag = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_21_real = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_21_imag = _RAND_3[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_24_real = _RAND_4[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_24_imag = _RAND_5[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_27_real = _RAND_6[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_27_imag = _RAND_7[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  feedback_real = _RAND_8[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  feedback_imag = _RAND_9[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  butt_out_0_real = _RAND_10[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  butt_out_0_imag = _RAND_11[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  load_output = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (io_en) begin
      shift_out_real <= _T_27_real;
    end
    if (io_en) begin
      shift_out_imag <= _T_27_imag;
    end
    if (io_en) begin
      if (load_input) begin
        _T_21_real <= io_in_real;
      end else begin
        _T_21_real <= butterfly_outputs_1_real;
      end
    end
    if (io_en) begin
      if (load_input) begin
        _T_21_imag <= io_in_imag;
      end else begin
        _T_21_imag <= butterfly_outputs_1_imag;
      end
    end
    if (io_en) begin
      _T_24_real <= _T_21_real;
    end
    if (io_en) begin
      _T_24_imag <= _T_21_imag;
    end
    if (io_en) begin
      _T_27_real <= _T_24_real;
    end
    if (io_en) begin
      _T_27_imag <= _T_24_imag;
    end
    feedback_real <= shift_out_real;
    feedback_imag <= shift_out_imag;
    butt_out_0_real <= _T_44[16:1];
    butt_out_0_imag <= _T_51[16:1];
    if (reset) begin
      load_output <= 1'h0;
    end else begin
      load_output <= load_input;
    end
  end
endmodule
module SDFStageRadix22_4(
  input         clock,
  input         reset,
  input  [15:0] io_in_real,
  input  [15:0] io_in_imag,
  output [15:0] io_out_real,
  output [15:0] io_out_imag,
  input  [5:0]  io_cntr,
  input         io_en
);
  wire  load_input; // @[SDFChainRadix22.scala 426:66]
  reg [15:0] shift_out_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_0;
  wire [16:0] butt_outputs_1_real; // @[FixedPointTypeClass.scala 33:22]
  wire [17:0] _T_50; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_52; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_55; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] butterfly_outputs_1_real; // @[FixedPointTypeClass.scala 176:41]
  reg [15:0] shift_out_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1;
  wire [16:0] butt_outputs_1_imag; // @[FixedPointTypeClass.scala 33:22]
  wire [17:0] _T_57; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_59; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_62; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] butterfly_outputs_1_imag; // @[FixedPointTypeClass.scala 176:41]
  reg [15:0] _T_21_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2;
  reg [15:0] _T_21_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3;
  wire [16:0] butt_outputs_0_real; // @[FixedPointTypeClass.scala 24:22]
  wire [16:0] butt_outputs_0_imag; // @[FixedPointTypeClass.scala 24:22]
  wire [17:0] _T_33; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_35; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_38; // @[FixedPointTypeClass.scala 20:58]
  wire [17:0] _T_40; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_42; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_45; // @[FixedPointTypeClass.scala 20:58]
  reg [15:0] feedback_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4;
  reg [15:0] feedback_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5;
  reg [15:0] butt_out_0_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6;
  reg [15:0] butt_out_0_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7;
  reg  load_output; // @[Reg.scala 27:20]
  reg [31:0] _RAND_8;
  assign load_input = io_cntr < 6'h2; // @[SDFChainRadix22.scala 426:66]
  assign butt_outputs_1_real = $signed(shift_out_real) - $signed(io_in_real); // @[FixedPointTypeClass.scala 33:22]
  assign _T_50 = {$signed(butt_outputs_1_real), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign _T_52 = _T_50[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign _T_55 = $signed(_T_52) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign butterfly_outputs_1_real = _T_55[16:1]; // @[FixedPointTypeClass.scala 176:41]
  assign butt_outputs_1_imag = $signed(shift_out_imag) - $signed(io_in_imag); // @[FixedPointTypeClass.scala 33:22]
  assign _T_57 = {$signed(butt_outputs_1_imag), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign _T_59 = _T_57[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign _T_62 = $signed(_T_59) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign butterfly_outputs_1_imag = _T_62[16:1]; // @[FixedPointTypeClass.scala 176:41]
  assign butt_outputs_0_real = $signed(shift_out_real) + $signed(io_in_real); // @[FixedPointTypeClass.scala 24:22]
  assign butt_outputs_0_imag = $signed(shift_out_imag) + $signed(io_in_imag); // @[FixedPointTypeClass.scala 24:22]
  assign _T_33 = {$signed(butt_outputs_0_real), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign _T_35 = _T_33[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign _T_38 = $signed(_T_35) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign _T_40 = {$signed(butt_outputs_0_imag), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign _T_42 = _T_40[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign _T_45 = $signed(_T_42) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign io_out_real = load_output ? $signed(feedback_real) : $signed(butt_out_0_real); // @[SDFChainRadix22.scala 422:10]
  assign io_out_imag = load_output ? $signed(feedback_imag) : $signed(butt_out_0_imag); // @[SDFChainRadix22.scala 422:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  shift_out_real = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  shift_out_imag = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_21_real = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_21_imag = _RAND_3[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  feedback_real = _RAND_4[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  feedback_imag = _RAND_5[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  butt_out_0_real = _RAND_6[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  butt_out_0_imag = _RAND_7[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  load_output = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (io_en) begin
      shift_out_real <= _T_21_real;
    end
    if (io_en) begin
      shift_out_imag <= _T_21_imag;
    end
    if (io_en) begin
      if (load_input) begin
        _T_21_real <= io_in_real;
      end else begin
        _T_21_real <= butterfly_outputs_1_real;
      end
    end
    if (io_en) begin
      if (load_input) begin
        _T_21_imag <= io_in_imag;
      end else begin
        _T_21_imag <= butterfly_outputs_1_imag;
      end
    end
    feedback_real <= shift_out_real;
    feedback_imag <= shift_out_imag;
    butt_out_0_real <= _T_38[16:1];
    butt_out_0_imag <= _T_45[16:1];
    if (reset) begin
      load_output <= 1'h0;
    end else begin
      load_output <= load_input;
    end
  end
endmodule
module SDFStageRadix22_5(
  input         clock,
  input         reset,
  input  [15:0] io_in_real,
  input  [15:0] io_in_imag,
  output [15:0] io_out_real,
  output [15:0] io_out_imag,
  input  [5:0]  io_cntr,
  input         io_en
);
  wire  load_input; // @[SDFChainRadix22.scala 426:66]
  reg [15:0] shift_out_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_0;
  wire [16:0] butt_outputs_1_real; // @[FixedPointTypeClass.scala 33:22]
  wire [17:0] _T_47; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_49; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_52; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] butterfly_outputs_1_real; // @[FixedPointTypeClass.scala 176:41]
  reg [15:0] shift_out_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1;
  wire [16:0] butt_outputs_1_imag; // @[FixedPointTypeClass.scala 33:22]
  wire [17:0] _T_54; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_56; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_59; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] butterfly_outputs_1_imag; // @[FixedPointTypeClass.scala 176:41]
  wire [16:0] butt_outputs_0_real; // @[FixedPointTypeClass.scala 24:22]
  wire [16:0] butt_outputs_0_imag; // @[FixedPointTypeClass.scala 24:22]
  wire [17:0] _T_30; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_32; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_35; // @[FixedPointTypeClass.scala 20:58]
  wire [17:0] _T_37; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_39; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_42; // @[FixedPointTypeClass.scala 20:58]
  reg [15:0] feedback_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2;
  reg [15:0] feedback_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3;
  reg [15:0] butt_out_0_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4;
  reg [15:0] butt_out_0_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5;
  reg  load_output; // @[Reg.scala 27:20]
  reg [31:0] _RAND_6;
  assign load_input = io_cntr < 6'h1; // @[SDFChainRadix22.scala 426:66]
  assign butt_outputs_1_real = $signed(shift_out_real) - $signed(io_in_real); // @[FixedPointTypeClass.scala 33:22]
  assign _T_47 = {$signed(butt_outputs_1_real), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign _T_49 = _T_47[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign _T_52 = $signed(_T_49) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign butterfly_outputs_1_real = _T_52[16:1]; // @[FixedPointTypeClass.scala 176:41]
  assign butt_outputs_1_imag = $signed(shift_out_imag) - $signed(io_in_imag); // @[FixedPointTypeClass.scala 33:22]
  assign _T_54 = {$signed(butt_outputs_1_imag), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign _T_56 = _T_54[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign _T_59 = $signed(_T_56) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign butterfly_outputs_1_imag = _T_59[16:1]; // @[FixedPointTypeClass.scala 176:41]
  assign butt_outputs_0_real = $signed(shift_out_real) + $signed(io_in_real); // @[FixedPointTypeClass.scala 24:22]
  assign butt_outputs_0_imag = $signed(shift_out_imag) + $signed(io_in_imag); // @[FixedPointTypeClass.scala 24:22]
  assign _T_30 = {$signed(butt_outputs_0_real), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign _T_32 = _T_30[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign _T_35 = $signed(_T_32) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign _T_37 = {$signed(butt_outputs_0_imag), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  assign _T_39 = _T_37[17:1]; // @[FixedPointTypeClass.scala 133:23]
  assign _T_42 = $signed(_T_39) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign io_out_real = load_output ? $signed(feedback_real) : $signed(butt_out_0_real); // @[SDFChainRadix22.scala 422:10]
  assign io_out_imag = load_output ? $signed(feedback_imag) : $signed(butt_out_0_imag); // @[SDFChainRadix22.scala 422:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  shift_out_real = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  shift_out_imag = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  feedback_real = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  feedback_imag = _RAND_3[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  butt_out_0_real = _RAND_4[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  butt_out_0_imag = _RAND_5[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  load_output = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (io_en) begin
      if (load_input) begin
        shift_out_real <= io_in_real;
      end else begin
        shift_out_real <= butterfly_outputs_1_real;
      end
    end
    if (io_en) begin
      if (load_input) begin
        shift_out_imag <= io_in_imag;
      end else begin
        shift_out_imag <= butterfly_outputs_1_imag;
      end
    end
    feedback_real <= shift_out_real;
    feedback_imag <= shift_out_imag;
    butt_out_0_real <= _T_35[16:1];
    butt_out_0_imag <= _T_42[16:1];
    if (reset) begin
      load_output <= 1'h0;
    end else begin
      load_output <= load_input;
    end
  end
endmodule
module Queue_10(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [15:0] io_enq_bits_real,
  input  [15:0] io_enq_bits_imag,
  input         io_deq_ready,
  output        io_deq_valid,
  output [15:0] io_deq_bits_real,
  output [15:0] io_deq_bits_imag
);
  reg [15:0] _T_4_real [0:24]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_0;
  wire [15:0] _T_4_real__T_26_data; // @[Decoupled.scala 209:24]
  wire [4:0] _T_4_real__T_26_addr; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_1;
  wire [15:0] _T_4_real__T_16_data; // @[Decoupled.scala 209:24]
  wire [4:0] _T_4_real__T_16_addr; // @[Decoupled.scala 209:24]
  wire  _T_4_real__T_16_mask; // @[Decoupled.scala 209:24]
  wire  _T_4_real__T_16_en; // @[Decoupled.scala 209:24]
  reg [15:0] _T_4_imag [0:24]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_2;
  wire [15:0] _T_4_imag__T_26_data; // @[Decoupled.scala 209:24]
  wire [4:0] _T_4_imag__T_26_addr; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_3;
  wire [15:0] _T_4_imag__T_16_data; // @[Decoupled.scala 209:24]
  wire [4:0] _T_4_imag__T_16_addr; // @[Decoupled.scala 209:24]
  wire  _T_4_imag__T_16_mask; // @[Decoupled.scala 209:24]
  wire  _T_4_imag__T_16_en; // @[Decoupled.scala 209:24]
  reg [4:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_4;
  reg [4:0] value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  reg  _T_5; // @[Decoupled.scala 212:35]
  reg [31:0] _RAND_6;
  wire  _T_6; // @[Decoupled.scala 214:41]
  wire  _T_7; // @[Decoupled.scala 215:36]
  wire  _T_8; // @[Decoupled.scala 215:33]
  wire  _T_9; // @[Decoupled.scala 216:32]
  wire  _T_10; // @[Decoupled.scala 40:37]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  wrap; // @[Counter.scala 38:24]
  wire [4:0] _T_18; // @[Counter.scala 39:22]
  wire  _GEN_12; // @[Decoupled.scala 240:27]
  wire  _GEN_16; // @[Decoupled.scala 237:18]
  wire  wrap_1; // @[Counter.scala 38:24]
  wire [4:0] _T_20; // @[Counter.scala 39:22]
  wire  _GEN_15; // @[Decoupled.scala 237:18]
  wire  _T_21; // @[Decoupled.scala 227:16]
  wire  _T_22; // @[Decoupled.scala 231:19]
  wire  _T_23; // @[Decoupled.scala 232:19]
  assign _T_4_real__T_26_addr = value_1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_4_real__T_26_data = _T_4_real[_T_4_real__T_26_addr]; // @[Decoupled.scala 209:24]
  `else
  assign _T_4_real__T_26_data = _T_4_real__T_26_addr >= 5'h19 ? _RAND_1[15:0] : _T_4_real[_T_4_real__T_26_addr]; // @[Decoupled.scala 209:24]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_4_real__T_16_data = io_enq_bits_real;
  assign _T_4_real__T_16_addr = value;
  assign _T_4_real__T_16_mask = 1'h1;
  assign _T_4_real__T_16_en = _T_8 ? _GEN_12 : _T_10;
  assign _T_4_imag__T_26_addr = value_1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_4_imag__T_26_data = _T_4_imag[_T_4_imag__T_26_addr]; // @[Decoupled.scala 209:24]
  `else
  assign _T_4_imag__T_26_data = _T_4_imag__T_26_addr >= 5'h19 ? _RAND_3[15:0] : _T_4_imag[_T_4_imag__T_26_addr]; // @[Decoupled.scala 209:24]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_4_imag__T_16_data = io_enq_bits_imag;
  assign _T_4_imag__T_16_addr = value;
  assign _T_4_imag__T_16_mask = 1'h1;
  assign _T_4_imag__T_16_en = _T_8 ? _GEN_12 : _T_10;
  assign _T_6 = value == value_1; // @[Decoupled.scala 214:41]
  assign _T_7 = ~_T_5; // @[Decoupled.scala 215:36]
  assign _T_8 = _T_6 & _T_7; // @[Decoupled.scala 215:33]
  assign _T_9 = _T_6 & _T_5; // @[Decoupled.scala 216:32]
  assign _T_10 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  assign _T_12 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  assign wrap = value == 5'h18; // @[Counter.scala 38:24]
  assign _T_18 = value + 5'h1; // @[Counter.scala 39:22]
  assign _GEN_12 = io_deq_ready ? 1'h0 : _T_10; // @[Decoupled.scala 240:27]
  assign _GEN_16 = _T_8 ? _GEN_12 : _T_10; // @[Decoupled.scala 237:18]
  assign wrap_1 = value_1 == 5'h18; // @[Counter.scala 38:24]
  assign _T_20 = value_1 + 5'h1; // @[Counter.scala 39:22]
  assign _GEN_15 = _T_8 ? 1'h0 : _T_12; // @[Decoupled.scala 237:18]
  assign _T_21 = _GEN_16 != _GEN_15; // @[Decoupled.scala 227:16]
  assign _T_22 = ~_T_8; // @[Decoupled.scala 231:19]
  assign _T_23 = ~_T_9; // @[Decoupled.scala 232:19]
  assign io_enq_ready = io_deq_ready | _T_23; // @[Decoupled.scala 232:16 Decoupled.scala 245:40]
  assign io_deq_valid = io_enq_valid | _T_22; // @[Decoupled.scala 231:16 Decoupled.scala 236:40]
  assign io_deq_bits_real = _T_8 ? $signed(io_enq_bits_real) : $signed(_T_4_real__T_26_data); // @[Decoupled.scala 233:15 Decoupled.scala 238:19]
  assign io_deq_bits_imag = _T_8 ? $signed(io_enq_bits_imag) : $signed(_T_4_imag__T_26_data); // @[Decoupled.scala 233:15 Decoupled.scala 238:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 25; initvar = initvar+1)
    _T_4_real[initvar] = _RAND_0[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  _RAND_2 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 25; initvar = initvar+1)
    _T_4_imag[initvar] = _RAND_2[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  value = _RAND_4[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value_1 = _RAND_5[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_5 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T_4_real__T_16_en & _T_4_real__T_16_mask) begin
      _T_4_real[_T_4_real__T_16_addr] <= _T_4_real__T_16_data; // @[Decoupled.scala 209:24]
    end
    if(_T_4_imag__T_16_en & _T_4_imag__T_16_mask) begin
      _T_4_imag[_T_4_imag__T_16_addr] <= _T_4_imag__T_16_data; // @[Decoupled.scala 209:24]
    end
    if (reset) begin
      value <= 5'h0;
    end else if (_GEN_16) begin
      if (wrap) begin
        value <= 5'h0;
      end else begin
        value <= _T_18;
      end
    end
    if (reset) begin
      value_1 <= 5'h0;
    end else if (_GEN_15) begin
      if (wrap_1) begin
        value_1 <= 5'h0;
      end else begin
        value_1 <= _T_20;
      end
    end
    if (reset) begin
      _T_5 <= 1'h0;
    end else if (_T_21) begin
      if (_T_8) begin
        if (io_deq_ready) begin
          _T_5 <= 1'h0;
        end else begin
          _T_5 <= _T_10;
        end
      end else begin
        _T_5 <= _T_10;
      end
    end
  end
endmodule
module SDFChainRadix22(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [15:0] io_in_bits_real,
  input  [15:0] io_in_bits_imag,
  input         io_out_ready,
  output        io_out_valid,
  output [15:0] io_out_bits_real,
  output [15:0] io_out_bits_imag,
  output        io_lastOut,
  input         io_lastIn,
  input  [5:0]  io_fftSize,
  output        io_busy
);
  wire  sdf_stages_0_clock; // @[SDFChainRadix22.scala 155:25]
  wire  sdf_stages_0_reset; // @[SDFChainRadix22.scala 155:25]
  wire [15:0] sdf_stages_0_io_in_real; // @[SDFChainRadix22.scala 155:25]
  wire [15:0] sdf_stages_0_io_in_imag; // @[SDFChainRadix22.scala 155:25]
  wire [15:0] sdf_stages_0_io_out_real; // @[SDFChainRadix22.scala 155:25]
  wire [15:0] sdf_stages_0_io_out_imag; // @[SDFChainRadix22.scala 155:25]
  wire [5:0] sdf_stages_0_io_cntr; // @[SDFChainRadix22.scala 155:25]
  wire  sdf_stages_0_io_en; // @[SDFChainRadix22.scala 155:25]
  wire  sdf_stages_1_clock; // @[SDFChainRadix22.scala 155:25]
  wire  sdf_stages_1_reset; // @[SDFChainRadix22.scala 155:25]
  wire [15:0] sdf_stages_1_io_in_real; // @[SDFChainRadix22.scala 155:25]
  wire [15:0] sdf_stages_1_io_in_imag; // @[SDFChainRadix22.scala 155:25]
  wire [15:0] sdf_stages_1_io_out_real; // @[SDFChainRadix22.scala 155:25]
  wire [15:0] sdf_stages_1_io_out_imag; // @[SDFChainRadix22.scala 155:25]
  wire [5:0] sdf_stages_1_io_cntr; // @[SDFChainRadix22.scala 155:25]
  wire  sdf_stages_1_io_en; // @[SDFChainRadix22.scala 155:25]
  wire  sdf_stages_2_clock; // @[SDFChainRadix22.scala 155:25]
  wire  sdf_stages_2_reset; // @[SDFChainRadix22.scala 155:25]
  wire [15:0] sdf_stages_2_io_in_real; // @[SDFChainRadix22.scala 155:25]
  wire [15:0] sdf_stages_2_io_in_imag; // @[SDFChainRadix22.scala 155:25]
  wire [15:0] sdf_stages_2_io_out_real; // @[SDFChainRadix22.scala 155:25]
  wire [15:0] sdf_stages_2_io_out_imag; // @[SDFChainRadix22.scala 155:25]
  wire [5:0] sdf_stages_2_io_cntr; // @[SDFChainRadix22.scala 155:25]
  wire  sdf_stages_2_io_en; // @[SDFChainRadix22.scala 155:25]
  wire  sdf_stages_3_clock; // @[SDFChainRadix22.scala 155:25]
  wire  sdf_stages_3_reset; // @[SDFChainRadix22.scala 155:25]
  wire [15:0] sdf_stages_3_io_in_real; // @[SDFChainRadix22.scala 155:25]
  wire [15:0] sdf_stages_3_io_in_imag; // @[SDFChainRadix22.scala 155:25]
  wire [15:0] sdf_stages_3_io_out_real; // @[SDFChainRadix22.scala 155:25]
  wire [15:0] sdf_stages_3_io_out_imag; // @[SDFChainRadix22.scala 155:25]
  wire [5:0] sdf_stages_3_io_cntr; // @[SDFChainRadix22.scala 155:25]
  wire  sdf_stages_3_io_en; // @[SDFChainRadix22.scala 155:25]
  wire  sdf_stages_4_clock; // @[SDFChainRadix22.scala 155:25]
  wire  sdf_stages_4_reset; // @[SDFChainRadix22.scala 155:25]
  wire [15:0] sdf_stages_4_io_in_real; // @[SDFChainRadix22.scala 155:25]
  wire [15:0] sdf_stages_4_io_in_imag; // @[SDFChainRadix22.scala 155:25]
  wire [15:0] sdf_stages_4_io_out_real; // @[SDFChainRadix22.scala 155:25]
  wire [15:0] sdf_stages_4_io_out_imag; // @[SDFChainRadix22.scala 155:25]
  wire [5:0] sdf_stages_4_io_cntr; // @[SDFChainRadix22.scala 155:25]
  wire  sdf_stages_4_io_en; // @[SDFChainRadix22.scala 155:25]
  wire  sdf_stages_5_clock; // @[SDFChainRadix22.scala 155:25]
  wire  sdf_stages_5_reset; // @[SDFChainRadix22.scala 155:25]
  wire [15:0] sdf_stages_5_io_in_real; // @[SDFChainRadix22.scala 155:25]
  wire [15:0] sdf_stages_5_io_in_imag; // @[SDFChainRadix22.scala 155:25]
  wire [15:0] sdf_stages_5_io_out_real; // @[SDFChainRadix22.scala 155:25]
  wire [15:0] sdf_stages_5_io_out_imag; // @[SDFChainRadix22.scala 155:25]
  wire [5:0] sdf_stages_5_io_cntr; // @[SDFChainRadix22.scala 155:25]
  wire  sdf_stages_5_io_en; // @[SDFChainRadix22.scala 155:25]
  wire  outQueue_clock; // @[SDFChainRadix22.scala 356:25]
  wire  outQueue_reset; // @[SDFChainRadix22.scala 356:25]
  wire  outQueue_io_enq_ready; // @[SDFChainRadix22.scala 356:25]
  wire  outQueue_io_enq_valid; // @[SDFChainRadix22.scala 356:25]
  wire [15:0] outQueue_io_enq_bits_real; // @[SDFChainRadix22.scala 356:25]
  wire [15:0] outQueue_io_enq_bits_imag; // @[SDFChainRadix22.scala 356:25]
  wire  outQueue_io_deq_ready; // @[SDFChainRadix22.scala 356:25]
  wire  outQueue_io_deq_valid; // @[SDFChainRadix22.scala 356:25]
  wire [15:0] outQueue_io_deq_bits_real; // @[SDFChainRadix22.scala 356:25]
  wire [15:0] outQueue_io_deq_bits_imag; // @[SDFChainRadix22.scala 356:25]
  reg [5:0] regNumStages; // @[SDFChainRadix22.scala 41:29]
  reg [31:0] _RAND_0;
  reg [1:0] state; // @[SDFChainRadix22.scala 52:22]
  reg [31:0] _RAND_1;
  reg  initialOutDone; // @[SDFChainRadix22.scala 55:31]
  reg [31:0] _RAND_2;
  reg [6:0] cnt; // @[SDFChainRadix22.scala 56:20]
  reg [31:0] _RAND_3;
  wire [5:0] _T_35; // @[SDFChainRadix22.scala 69:39]
  wire [64:0] _T_36; // @[SDFChainRadix22.scala 69:23]
  wire  _T_37; // @[Decoupled.scala 40:37]
  wire  fireLast; // @[SDFChainRadix22.scala 75:28]
  wire  _T_38; // @[Conditional.scala 37:30]
  wire [1:0] _GEN_0; // @[SDFChainRadix22.scala 82:27]
  wire  _T_41; // @[Conditional.scala 37:30]
  wire [1:0] _GEN_1; // @[SDFChainRadix22.scala 85:23]
  wire  _T_42; // @[Conditional.scala 37:30]
  wire [1:0] _GEN_2; // @[SDFChainRadix22.scala 90:25]
  wire [1:0] _GEN_3; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_4; // @[Conditional.scala 39:67]
  wire [1:0] state_next; // @[Conditional.scala 40:58]
  reg [5:0] cntValidOut; // @[SDFChainRadix22.scala 99:28]
  reg [31:0] _RAND_4;
  reg  lastWait; // @[SDFChainRadix22.scala 100:25]
  reg [31:0] _RAND_5;
  reg  lastIndeed; // @[SDFChainRadix22.scala 101:27]
  reg [31:0] _RAND_6;
  reg  initialInDone; // @[SDFChainRadix22.scala 102:30]
  reg [31:0] _RAND_7;
  reg  initialInDonePrev; // @[SDFChainRadix22.scala 103:34]
  reg [31:0] _RAND_8;
  wire [6:0] numPoints; // @[SDFChainRadix22.scala 46:23 SDFChainRadix22.scala 69:15]
  wire [6:0] _T_44; // @[SDFChainRadix22.scala 104:44]
  wire [6:0] _GEN_576; // @[SDFChainRadix22.scala 104:29]
  wire  _T_45; // @[SDFChainRadix22.scala 104:29]
  wire  _T_46; // @[Decoupled.scala 40:37]
  wire  pktEnd; // @[SDFChainRadix22.scala 104:52]
  wire  _T_47; // @[SDFChainRadix22.scala 106:20]
  wire  _T_50; // @[SDFChainRadix22.scala 109:18]
  wire  _T_52; // @[SDFChainRadix22.scala 109:40]
  wire  _GEN_14; // @[SDFChainRadix22.scala 109:57]
  wire  _T_54; // @[SDFChainRadix22.scala 117:41]
  wire  _T_55; // @[SDFChainRadix22.scala 117:23]
  wire  _GEN_16; // @[SDFChainRadix22.scala 117:64]
  wire  _T_57; // @[SDFChainRadix22.scala 121:30]
  wire [5:0] _T_60; // @[SDFChainRadix22.scala 125:32]
  wire  _T_62; // @[SDFChainRadix22.scala 131:23]
  wire  _GEN_20; // @[SDFChainRadix22.scala 131:34]
  wire  _T_63; // @[SDFChainRadix22.scala 135:132]
  wire  _T_64; // @[SDFChainRadix22.scala 135:159]
  wire  _T_65; // @[SDFChainRadix22.scala 135:150]
  wire [5:0] _T_67; // @[SDFChainRadix22.scala 138:62]
  wire [5:0] _GEN_23; // @[SDFChainRadix22.scala 138:25]
  wire [5:0] _GEN_24; // @[SDFChainRadix22.scala 138:25]
  wire [5:0] _GEN_25; // @[SDFChainRadix22.scala 138:25]
  wire [5:0] _GEN_26; // @[SDFChainRadix22.scala 138:25]
  wire [5:0] _GEN_27; // @[SDFChainRadix22.scala 138:25]
  wire [5:0] cumulativeDelayWire; // @[SDFChainRadix22.scala 138:25]
  wire  activeStages_0; // @[SDFChainRadix22.scala 146:48]
  wire  activeStages_1; // @[SDFChainRadix22.scala 146:48]
  wire  activeStages_2; // @[SDFChainRadix22.scala 146:48]
  wire  activeStages_3; // @[SDFChainRadix22.scala 146:48]
  wire  activeStages_4; // @[SDFChainRadix22.scala 146:48]
  wire  activeStages_5; // @[SDFChainRadix22.scala 146:48]
  wire  _T_95; // @[SDFChainRadix22.scala 164:54]
  wire  enableInit; // @[SDFChainRadix22.scala 164:33]
  wire [6:0] _T_98; // @[SDFChainRadix22.scala 170:16]
  reg  _T_100; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_9;
  reg  _T_101; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_10;
  reg  _T_102; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_11;
  reg  enableVector_1; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_12;
  reg [6:0] _T_105; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_13;
  reg [6:0] _T_106; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_14;
  reg [6:0] _T_107; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_15;
  reg [6:0] _T_108; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_16;
  reg  _T_110; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_17;
  reg  _T_111; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_18;
  reg  _T_112; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_19;
  reg  enableVector_2; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_20;
  reg [6:0] _T_115; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_21;
  reg [6:0] _T_116; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_22;
  reg [6:0] _T_117; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_23;
  reg [6:0] _T_118; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_24;
  reg  _T_120; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_25;
  reg  _T_121; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_26;
  reg  _T_122; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_27;
  reg  enableVector_3; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_28;
  reg [6:0] _T_125; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_29;
  reg [6:0] _T_126; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_30;
  reg [6:0] _T_127; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_31;
  reg [6:0] _T_128; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_32;
  reg  _T_130; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_33;
  reg  _T_131; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_34;
  reg  _T_132; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_35;
  reg  enableVector_4; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_36;
  reg [6:0] _T_135; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_37;
  reg [6:0] _T_136; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_38;
  reg [6:0] _T_137; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_39;
  reg [6:0] _T_138; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_40;
  reg  _T_140; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_41;
  reg  _T_141; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_42;
  reg  _T_142; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_43;
  reg  enableVector_5; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_44;
  reg [6:0] _T_145; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_45;
  reg [6:0] _T_146; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_46;
  reg [6:0] _T_147; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_47;
  reg [6:0] _T_148; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_48;
  wire [6:0] _T_166; // @[SDFChainRadix22.scala 186:37]
  wire [5:0] cntr_wires_0; // @[SDFChainRadix22.scala 48:24 SDFChainRadix22.scala 176:29]
  wire [5:0] cntr_wires_1; // @[SDFChainRadix22.scala 48:24 SDFChainRadix22.scala 176:29]
  wire [5:0] _GEN_128; // @[SDFChainRadix22.scala 186:22]
  wire [5:0] cntr_wires_2; // @[SDFChainRadix22.scala 48:24 SDFChainRadix22.scala 176:29]
  wire [5:0] _GEN_129; // @[SDFChainRadix22.scala 186:22]
  wire [5:0] cntr_wires_3; // @[SDFChainRadix22.scala 48:24 SDFChainRadix22.scala 176:29]
  wire [5:0] _GEN_130; // @[SDFChainRadix22.scala 186:22]
  wire [5:0] cntr_wires_4; // @[SDFChainRadix22.scala 48:24 SDFChainRadix22.scala 176:29]
  wire [5:0] _GEN_131; // @[SDFChainRadix22.scala 186:22]
  wire [5:0] cntr_wires_5; // @[SDFChainRadix22.scala 48:24 SDFChainRadix22.scala 176:29]
  wire [5:0] _GEN_132; // @[SDFChainRadix22.scala 186:22]
  wire [6:0] _GEN_577; // @[SDFChainRadix22.scala 186:22]
  wire  _T_167; // @[SDFChainRadix22.scala 186:22]
  wire  _GEN_134; // @[SDFChainRadix22.scala 186:44]
  wire  _GEN_135; // @[SDFChainRadix22.scala 186:44]
  wire  _GEN_136; // @[SDFChainRadix22.scala 186:44]
  wire  _GEN_137; // @[SDFChainRadix22.scala 186:44]
  wire  _GEN_138; // @[SDFChainRadix22.scala 186:44]
  wire  _T_168; // @[SDFChainRadix22.scala 186:44]
  wire  _GEN_139; // @[SDFChainRadix22.scala 189:36]
  wire  _GEN_140; // @[SDFChainRadix22.scala 186:60]
  wire  _T_170; // @[SDFChainRadix22.scala 193:43]
  reg  _T_171; // @[SDFChainRadix22.scala 193:59]
  reg [31:0] _RAND_49;
  wire  _T_173; // @[SDFChainRadix22.scala 193:72]
  wire  _T_174; // @[SDFChainRadix22.scala 193:101]
  wire [15:0] input_data_real; // @[SDFChainRadix22.scala 211:23]
  wire [15:0] input_data_imag; // @[SDFChainRadix22.scala 211:23]
  wire  _T_184; // @[SDFChainRadix22.scala 214:67]
  wire [5:0] _T_188; // @[SDFChainRadix22.scala 215:63]
  wire  _GEN_144; // @[SDFChainRadix22.scala 216:20]
  wire  _GEN_145; // @[SDFChainRadix22.scala 216:20]
  wire  _GEN_146; // @[SDFChainRadix22.scala 216:20]
  wire  _GEN_147; // @[SDFChainRadix22.scala 216:20]
  wire  _GEN_148; // @[SDFChainRadix22.scala 216:20]
  wire [5:0] _T_193; // @[SDFChainRadix22.scala 217:68]
  wire [5:0] _GEN_150; // @[SDFChainRadix22.scala 217:38]
  wire [5:0] _GEN_151; // @[SDFChainRadix22.scala 217:38]
  wire [5:0] _GEN_152; // @[SDFChainRadix22.scala 217:38]
  wire [5:0] _GEN_153; // @[SDFChainRadix22.scala 217:38]
  wire [5:0] _GEN_154; // @[SDFChainRadix22.scala 217:38]
  wire  _T_199; // @[SDFChainRadix22.scala 214:67]
  wire [5:0] _T_203; // @[SDFChainRadix22.scala 215:63]
  wire  _GEN_156; // @[SDFChainRadix22.scala 216:20]
  wire  _GEN_157; // @[SDFChainRadix22.scala 216:20]
  wire  _GEN_158; // @[SDFChainRadix22.scala 216:20]
  wire  _GEN_159; // @[SDFChainRadix22.scala 216:20]
  wire  _GEN_160; // @[SDFChainRadix22.scala 216:20]
  wire [5:0] _T_208; // @[SDFChainRadix22.scala 217:68]
  wire [5:0] _GEN_162; // @[SDFChainRadix22.scala 217:38]
  wire [5:0] _GEN_163; // @[SDFChainRadix22.scala 217:38]
  wire [5:0] _GEN_164; // @[SDFChainRadix22.scala 217:38]
  wire [5:0] _GEN_165; // @[SDFChainRadix22.scala 217:38]
  wire [5:0] _GEN_166; // @[SDFChainRadix22.scala 217:38]
  wire [5:0] _T_210; // @[SDFChainRadix22.scala 217:38]
  wire  _T_214; // @[SDFChainRadix22.scala 214:67]
  wire [5:0] _T_218; // @[SDFChainRadix22.scala 215:63]
  wire  _GEN_168; // @[SDFChainRadix22.scala 216:20]
  wire  _GEN_169; // @[SDFChainRadix22.scala 216:20]
  wire  _GEN_170; // @[SDFChainRadix22.scala 216:20]
  wire  _GEN_171; // @[SDFChainRadix22.scala 216:20]
  wire  _GEN_172; // @[SDFChainRadix22.scala 216:20]
  wire [5:0] _T_223; // @[SDFChainRadix22.scala 217:68]
  wire [5:0] _GEN_174; // @[SDFChainRadix22.scala 217:38]
  wire [5:0] _GEN_175; // @[SDFChainRadix22.scala 217:38]
  wire [5:0] _GEN_176; // @[SDFChainRadix22.scala 217:38]
  wire [5:0] _GEN_177; // @[SDFChainRadix22.scala 217:38]
  wire [5:0] _GEN_178; // @[SDFChainRadix22.scala 217:38]
  wire [5:0] _T_225; // @[SDFChainRadix22.scala 217:38]
  wire  _T_229; // @[SDFChainRadix22.scala 214:67]
  wire [5:0] _T_233; // @[SDFChainRadix22.scala 215:63]
  wire  _GEN_180; // @[SDFChainRadix22.scala 216:20]
  wire  _GEN_181; // @[SDFChainRadix22.scala 216:20]
  wire  _GEN_182; // @[SDFChainRadix22.scala 216:20]
  wire  _GEN_183; // @[SDFChainRadix22.scala 216:20]
  wire  _GEN_184; // @[SDFChainRadix22.scala 216:20]
  wire [5:0] _T_238; // @[SDFChainRadix22.scala 217:68]
  wire [5:0] _GEN_186; // @[SDFChainRadix22.scala 217:38]
  wire [5:0] _GEN_187; // @[SDFChainRadix22.scala 217:38]
  wire [5:0] _GEN_188; // @[SDFChainRadix22.scala 217:38]
  wire [5:0] _GEN_189; // @[SDFChainRadix22.scala 217:38]
  wire [5:0] _GEN_190; // @[SDFChainRadix22.scala 217:38]
  wire [5:0] _T_240; // @[SDFChainRadix22.scala 217:38]
  wire  _T_244; // @[SDFChainRadix22.scala 214:67]
  wire [5:0] _T_248; // @[SDFChainRadix22.scala 215:63]
  wire  _GEN_192; // @[SDFChainRadix22.scala 216:20]
  wire  _GEN_193; // @[SDFChainRadix22.scala 216:20]
  wire  _GEN_194; // @[SDFChainRadix22.scala 216:20]
  wire  _GEN_195; // @[SDFChainRadix22.scala 216:20]
  wire  _GEN_196; // @[SDFChainRadix22.scala 216:20]
  wire [5:0] _T_253; // @[SDFChainRadix22.scala 217:68]
  wire [5:0] _GEN_198; // @[SDFChainRadix22.scala 217:38]
  wire [5:0] _GEN_199; // @[SDFChainRadix22.scala 217:38]
  wire [5:0] _GEN_200; // @[SDFChainRadix22.scala 217:38]
  wire [5:0] _GEN_201; // @[SDFChainRadix22.scala 217:38]
  wire [5:0] _GEN_202; // @[SDFChainRadix22.scala 217:38]
  wire [5:0] _T_255; // @[SDFChainRadix22.scala 217:38]
  wire  _T_259; // @[SDFChainRadix22.scala 214:67]
  wire [5:0] _T_263; // @[SDFChainRadix22.scala 215:63]
  wire  _GEN_204; // @[SDFChainRadix22.scala 216:20]
  wire  _GEN_205; // @[SDFChainRadix22.scala 216:20]
  wire  _GEN_206; // @[SDFChainRadix22.scala 216:20]
  wire  _GEN_207; // @[SDFChainRadix22.scala 216:20]
  wire  _GEN_208; // @[SDFChainRadix22.scala 216:20]
  wire [5:0] _T_268; // @[SDFChainRadix22.scala 217:68]
  wire [5:0] _GEN_210; // @[SDFChainRadix22.scala 217:38]
  wire [5:0] _GEN_211; // @[SDFChainRadix22.scala 217:38]
  wire [5:0] _GEN_212; // @[SDFChainRadix22.scala 217:38]
  wire [5:0] _GEN_213; // @[SDFChainRadix22.scala 217:38]
  wire [5:0] _GEN_214; // @[SDFChainRadix22.scala 217:38]
  wire [5:0] _T_270; // @[SDFChainRadix22.scala 217:38]
  wire  _T_277; // @[SDFChainRadix22.scala 234:23]
  wire [15:0] _GEN_215; // @[SDFChainRadix22.scala 234:55]
  wire [15:0] _GEN_216; // @[SDFChainRadix22.scala 234:55]
  wire  _T_278; // @[SDFChainRadix22.scala 320:98]
  wire  _T_280; // @[SDFChainRadix22.scala 320:135]
  wire  _T_281; // @[SDFChainRadix22.scala 320:122]
  reg  _T_283; // @[Reg.scala 15:16]
  reg [31:0] _RAND_50;
  wire [15:0] _T_289; // @[FixedPointTypeClass.scala 39:43]
  wire [15:0] _T_286_real; // @[SDFChainRadix22.scala 322:32 SDFChainRadix22.scala 325:29]
  reg [15:0] _T_295_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_51;
  reg [15:0] _T_295_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_52;
  reg [15:0] _T_298_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_53;
  reg [15:0] _T_298_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_54;
  reg [15:0] outputWires_0_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_55;
  reg [15:0] outputWires_0_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_56;
  wire  _T_307; // @[SDFChainRadix22.scala 234:23]
  wire [15:0] _GEN_226; // @[SDFChainRadix22.scala 234:55]
  wire [15:0] _GEN_227; // @[SDFChainRadix22.scala 234:55]
  wire [5:0] _T_475; // @[SDFChainRadix22.scala 276:83]
  wire [5:0] _T_479; // @[SDFChainRadix22.scala 276:89]
  reg [5:0] _T_481; // @[Reg.scala 15:16]
  reg [31:0] _RAND_57;
  reg [15:0] twiddles_1_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_58;
  reg [15:0] twiddles_1_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_59;
  wire [4:0] _GEN_266; // @[Reg.scala 16:23]
  wire [4:0] _GEN_267; // @[Reg.scala 16:23]
  wire [4:0] _GEN_268; // @[Reg.scala 16:23]
  wire [4:0] _GEN_269; // @[Reg.scala 16:23]
  wire [4:0] _GEN_270; // @[Reg.scala 16:23]
  wire [4:0] _GEN_271; // @[Reg.scala 16:23]
  wire [4:0] _GEN_272; // @[Reg.scala 16:23]
  wire [4:0] _GEN_273; // @[Reg.scala 16:23]
  wire [4:0] _GEN_274; // @[Reg.scala 16:23]
  wire [4:0] _GEN_275; // @[Reg.scala 16:23]
  wire [4:0] _GEN_276; // @[Reg.scala 16:23]
  wire [4:0] _GEN_277; // @[Reg.scala 16:23]
  wire [4:0] _GEN_278; // @[Reg.scala 16:23]
  wire [4:0] _GEN_279; // @[Reg.scala 16:23]
  wire [4:0] _GEN_280; // @[Reg.scala 16:23]
  wire [4:0] _GEN_281; // @[Reg.scala 16:23]
  wire [4:0] _GEN_282; // @[Reg.scala 16:23]
  wire [4:0] _GEN_283; // @[Reg.scala 16:23]
  wire [4:0] _GEN_284; // @[Reg.scala 16:23]
  wire [4:0] _GEN_285; // @[Reg.scala 16:23]
  wire [4:0] _GEN_286; // @[Reg.scala 16:23]
  wire [4:0] _GEN_287; // @[Reg.scala 16:23]
  wire [4:0] _GEN_288; // @[Reg.scala 16:23]
  wire [4:0] _GEN_289; // @[Reg.scala 16:23]
  wire [4:0] _GEN_290; // @[Reg.scala 16:23]
  wire [4:0] _GEN_291; // @[Reg.scala 16:23]
  wire [4:0] _GEN_292; // @[Reg.scala 16:23]
  wire [4:0] _GEN_293; // @[Reg.scala 16:23]
  wire [4:0] _GEN_294; // @[Reg.scala 16:23]
  wire [4:0] _GEN_295; // @[Reg.scala 16:23]
  wire [4:0] _GEN_296; // @[Reg.scala 16:23]
  wire [4:0] _GEN_297; // @[Reg.scala 16:23]
  wire [4:0] _GEN_298; // @[Reg.scala 16:23]
  wire [4:0] _GEN_299; // @[Reg.scala 16:23]
  wire [4:0] _GEN_300; // @[Reg.scala 16:23]
  wire [4:0] _GEN_301; // @[Reg.scala 16:23]
  wire [4:0] _GEN_302; // @[Reg.scala 16:23]
  wire [4:0] _GEN_303; // @[Reg.scala 16:23]
  wire [4:0] _GEN_304; // @[Reg.scala 16:23]
  wire [4:0] _GEN_305; // @[Reg.scala 16:23]
  wire [4:0] _GEN_306; // @[Reg.scala 16:23]
  wire [4:0] _GEN_307; // @[Reg.scala 16:23]
  wire [4:0] _GEN_308; // @[Reg.scala 16:23]
  wire [4:0] _GEN_309; // @[Reg.scala 16:23]
  wire [4:0] _GEN_310; // @[Reg.scala 16:23]
  wire [4:0] _GEN_311; // @[Reg.scala 16:23]
  wire [4:0] _GEN_312; // @[Reg.scala 16:23]
  reg [15:0] _T_490; // @[Reg.scala 15:16]
  reg [31:0] _RAND_60;
  reg [15:0] _T_491; // @[Reg.scala 15:16]
  reg [31:0] _RAND_61;
  reg [15:0] _T_492; // @[Reg.scala 15:16]
  reg [31:0] _RAND_62;
  reg [16:0] _T_494; // @[Reg.scala 15:16]
  reg [31:0] _RAND_63;
  reg [16:0] _T_496; // @[Reg.scala 15:16]
  reg [31:0] _RAND_64;
  reg [16:0] _T_498; // @[Reg.scala 15:16]
  reg [31:0] _RAND_65;
  wire [16:0] _GEN_578; // @[FixedPointTypeClass.scala 211:35]
  reg [32:0] _T_500; // @[Reg.scala 15:16]
  reg [63:0] _RAND_66;
  wire [34:0] _GEN_579; // @[FixedPointTypeClass.scala 20:58]
  wire [34:0] _T_503; // @[FixedPointTypeClass.scala 20:58]
  wire [33:0] _T_504; // @[FixedPointTypeClass.scala 176:41]
  wire [16:0] _GEN_580; // @[FixedPointTypeClass.scala 211:35]
  reg [32:0] _T_506; // @[Reg.scala 15:16]
  reg [63:0] _RAND_67;
  wire [34:0] _GEN_581; // @[FixedPointTypeClass.scala 20:58]
  wire [34:0] _T_509; // @[FixedPointTypeClass.scala 20:58]
  wire [33:0] _T_510; // @[FixedPointTypeClass.scala 176:41]
  wire [16:0] _GEN_582; // @[FixedPointTypeClass.scala 211:35]
  reg [32:0] _T_512; // @[Reg.scala 15:16]
  reg [63:0] _RAND_68;
  wire [34:0] _GEN_583; // @[FixedPointTypeClass.scala 20:58]
  wire [34:0] _T_515; // @[FixedPointTypeClass.scala 20:58]
  wire [33:0] _T_516; // @[FixedPointTypeClass.scala 176:41]
  reg [34:0] _T_518; // @[Reg.scala 15:16]
  reg [63:0] _RAND_69;
  reg [34:0] _T_520; // @[Reg.scala 15:16]
  reg [63:0] _RAND_70;
  wire [34:0] _T_526; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] _T_527; // @[FixedPointTypeClass.scala 176:41]
  wire [34:0] _T_530; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] _T_531; // @[FixedPointTypeClass.scala 176:41]
  wire  _T_540; // @[SDFChainRadix22.scala 234:23]
  wire [15:0] outputWires_1_imag; // @[SDFChainRadix22.scala 286:27 SDFChainRadix22.scala 306:19]
  wire [15:0] _GEN_450; // @[SDFChainRadix22.scala 234:55]
  wire [15:0] outputWires_1_real; // @[SDFChainRadix22.scala 286:27 SDFChainRadix22.scala 306:19]
  wire [15:0] _GEN_451; // @[SDFChainRadix22.scala 234:55]
  wire  _T_541; // @[SDFChainRadix22.scala 320:98]
  wire  _T_543; // @[SDFChainRadix22.scala 320:135]
  wire  _T_544; // @[SDFChainRadix22.scala 320:122]
  reg  _T_546; // @[Reg.scala 15:16]
  reg [31:0] _RAND_71;
  wire [15:0] _T_552; // @[FixedPointTypeClass.scala 39:43]
  wire [15:0] _T_549_real; // @[SDFChainRadix22.scala 322:32 SDFChainRadix22.scala 325:29]
  reg [15:0] _T_558_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_72;
  reg [15:0] _T_558_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_73;
  reg [15:0] _T_561_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_74;
  reg [15:0] _T_561_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_75;
  reg [15:0] outputWires_2_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_76;
  reg [15:0] outputWires_2_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_77;
  wire  _T_570; // @[SDFChainRadix22.scala 234:23]
  wire [15:0] _GEN_461; // @[SDFChainRadix22.scala 234:55]
  wire [15:0] _GEN_462; // @[SDFChainRadix22.scala 234:55]
  wire [5:0] _T_618; // @[SDFChainRadix22.scala 276:83]
  wire [5:0] _T_622; // @[SDFChainRadix22.scala 276:89]
  reg [5:0] _T_624; // @[Reg.scala 15:16]
  reg [31:0] _RAND_78;
  reg [15:0] twiddles_3_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_79;
  reg [15:0] twiddles_3_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_80;
  wire [2:0] _GEN_489; // @[Reg.scala 16:23]
  wire [2:0] _GEN_490; // @[Reg.scala 16:23]
  wire [2:0] _GEN_491; // @[Reg.scala 16:23]
  wire [2:0] _GEN_492; // @[Reg.scala 16:23]
  wire [2:0] _GEN_493; // @[Reg.scala 16:23]
  wire [2:0] _GEN_494; // @[Reg.scala 16:23]
  wire [2:0] _GEN_495; // @[Reg.scala 16:23]
  wire [2:0] _GEN_496; // @[Reg.scala 16:23]
  wire [2:0] _GEN_497; // @[Reg.scala 16:23]
  wire [2:0] _GEN_498; // @[Reg.scala 16:23]
  wire [2:0] _GEN_499; // @[Reg.scala 16:23]
  reg [15:0] _T_634; // @[Reg.scala 15:16]
  reg [31:0] _RAND_81;
  reg [15:0] _T_635; // @[Reg.scala 15:16]
  reg [31:0] _RAND_82;
  reg [15:0] _T_636; // @[Reg.scala 15:16]
  reg [31:0] _RAND_83;
  reg [16:0] _T_638; // @[Reg.scala 15:16]
  reg [31:0] _RAND_84;
  reg [16:0] _T_640; // @[Reg.scala 15:16]
  reg [31:0] _RAND_85;
  reg [16:0] _T_642; // @[Reg.scala 15:16]
  reg [31:0] _RAND_86;
  wire [16:0] _GEN_586; // @[FixedPointTypeClass.scala 211:35]
  reg [32:0] _T_644; // @[Reg.scala 15:16]
  reg [63:0] _RAND_87;
  wire [34:0] _GEN_587; // @[FixedPointTypeClass.scala 20:58]
  wire [34:0] _T_647; // @[FixedPointTypeClass.scala 20:58]
  wire [33:0] _T_648; // @[FixedPointTypeClass.scala 176:41]
  wire [16:0] _GEN_588; // @[FixedPointTypeClass.scala 211:35]
  reg [32:0] _T_650; // @[Reg.scala 15:16]
  reg [63:0] _RAND_88;
  wire [34:0] _GEN_589; // @[FixedPointTypeClass.scala 20:58]
  wire [34:0] _T_653; // @[FixedPointTypeClass.scala 20:58]
  wire [33:0] _T_654; // @[FixedPointTypeClass.scala 176:41]
  wire [16:0] _GEN_590; // @[FixedPointTypeClass.scala 211:35]
  reg [32:0] _T_656; // @[Reg.scala 15:16]
  reg [63:0] _RAND_89;
  wire [34:0] _GEN_591; // @[FixedPointTypeClass.scala 20:58]
  wire [34:0] _T_659; // @[FixedPointTypeClass.scala 20:58]
  wire [33:0] _T_660; // @[FixedPointTypeClass.scala 176:41]
  reg [34:0] _T_662; // @[Reg.scala 15:16]
  reg [63:0] _RAND_90;
  reg [34:0] _T_664; // @[Reg.scala 15:16]
  reg [63:0] _RAND_91;
  wire [34:0] _T_670; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] _T_671; // @[FixedPointTypeClass.scala 176:41]
  wire [34:0] _T_674; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] _T_675; // @[FixedPointTypeClass.scala 176:41]
  wire  _T_684; // @[SDFChainRadix22.scala 234:23]
  wire [15:0] outputWires_3_imag; // @[SDFChainRadix22.scala 286:27 SDFChainRadix22.scala 306:19]
  wire [15:0] _GEN_541; // @[SDFChainRadix22.scala 234:55]
  wire [15:0] outputWires_3_real; // @[SDFChainRadix22.scala 286:27 SDFChainRadix22.scala 306:19]
  wire [15:0] _GEN_542; // @[SDFChainRadix22.scala 234:55]
  wire  _T_685; // @[SDFChainRadix22.scala 320:98]
  wire  _T_687; // @[SDFChainRadix22.scala 320:135]
  wire  _T_688; // @[SDFChainRadix22.scala 320:122]
  reg  _T_690; // @[Reg.scala 15:16]
  reg [31:0] _RAND_92;
  wire [15:0] _T_696; // @[FixedPointTypeClass.scala 39:43]
  wire [15:0] _T_693_real; // @[SDFChainRadix22.scala 322:32 SDFChainRadix22.scala 325:29]
  reg [15:0] _T_702_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_93;
  reg [15:0] _T_702_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_94;
  reg [15:0] _T_705_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_95;
  reg [15:0] _T_705_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_96;
  reg [15:0] outputWires_4_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_97;
  reg [15:0] outputWires_4_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_98;
  wire  _T_714; // @[SDFChainRadix22.scala 234:23]
  wire [15:0] _GEN_552; // @[SDFChainRadix22.scala 234:55]
  wire [15:0] _GEN_553; // @[SDFChainRadix22.scala 234:55]
  reg [15:0] _T_717_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_99;
  reg [15:0] _T_717_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_100;
  reg [15:0] _T_720_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_101;
  reg [15:0] _T_720_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_102;
  reg [15:0] outputWires_5_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_103;
  reg [15:0] outputWires_5_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_104;
  reg  _T_725; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_105;
  reg  _T_726; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_106;
  reg  _T_727; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_107;
  reg  outValid; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_108;
  wire  _T_728; // @[SDFChainRadix22.scala 361:33]
  reg  _T_729; // @[Reg.scala 27:20]
  reg [31:0] _RAND_109;
  reg  _T_730; // @[Reg.scala 27:20]
  reg [31:0] _RAND_110;
  reg  _T_731; // @[Reg.scala 27:20]
  reg [31:0] _RAND_111;
  reg  _T_732; // @[Reg.scala 27:20]
  reg [31:0] _RAND_112;
  wire  _T_733; // @[SDFChainRadix22.scala 361:127]
  wire  _T_734; // @[SDFChainRadix22.scala 361:117]
  wire [29:0] _GEN_594; // @[SDFChainRadix22.scala 375:33]
  wire [31:0] _GEN_574; // @[SDFChainRadix22.scala 375:33]
  wire [29:0] _GEN_595; // @[SDFChainRadix22.scala 375:33]
  wire [31:0] _GEN_575; // @[SDFChainRadix22.scala 375:33]
  wire [17:0] _GEN_596; // @[SDFChainRadix22.scala 59:26 SDFChainRadix22.scala 376:20 SDFChainRadix22.scala 379:25]
  wire [17:0] _GEN_598; // @[SDFChainRadix22.scala 59:26 SDFChainRadix22.scala 376:20 SDFChainRadix22.scala 380:25]
  SDFStageRadix22 sdf_stages_0 ( // @[SDFChainRadix22.scala 155:25]
    .clock(sdf_stages_0_clock),
    .reset(sdf_stages_0_reset),
    .io_in_real(sdf_stages_0_io_in_real),
    .io_in_imag(sdf_stages_0_io_in_imag),
    .io_out_real(sdf_stages_0_io_out_real),
    .io_out_imag(sdf_stages_0_io_out_imag),
    .io_cntr(sdf_stages_0_io_cntr),
    .io_en(sdf_stages_0_io_en)
  );
  SDFStageRadix22_1 sdf_stages_1 ( // @[SDFChainRadix22.scala 155:25]
    .clock(sdf_stages_1_clock),
    .reset(sdf_stages_1_reset),
    .io_in_real(sdf_stages_1_io_in_real),
    .io_in_imag(sdf_stages_1_io_in_imag),
    .io_out_real(sdf_stages_1_io_out_real),
    .io_out_imag(sdf_stages_1_io_out_imag),
    .io_cntr(sdf_stages_1_io_cntr),
    .io_en(sdf_stages_1_io_en)
  );
  SDFStageRadix22_2 sdf_stages_2 ( // @[SDFChainRadix22.scala 155:25]
    .clock(sdf_stages_2_clock),
    .reset(sdf_stages_2_reset),
    .io_in_real(sdf_stages_2_io_in_real),
    .io_in_imag(sdf_stages_2_io_in_imag),
    .io_out_real(sdf_stages_2_io_out_real),
    .io_out_imag(sdf_stages_2_io_out_imag),
    .io_cntr(sdf_stages_2_io_cntr),
    .io_en(sdf_stages_2_io_en)
  );
  SDFStageRadix22_3 sdf_stages_3 ( // @[SDFChainRadix22.scala 155:25]
    .clock(sdf_stages_3_clock),
    .reset(sdf_stages_3_reset),
    .io_in_real(sdf_stages_3_io_in_real),
    .io_in_imag(sdf_stages_3_io_in_imag),
    .io_out_real(sdf_stages_3_io_out_real),
    .io_out_imag(sdf_stages_3_io_out_imag),
    .io_cntr(sdf_stages_3_io_cntr),
    .io_en(sdf_stages_3_io_en)
  );
  SDFStageRadix22_4 sdf_stages_4 ( // @[SDFChainRadix22.scala 155:25]
    .clock(sdf_stages_4_clock),
    .reset(sdf_stages_4_reset),
    .io_in_real(sdf_stages_4_io_in_real),
    .io_in_imag(sdf_stages_4_io_in_imag),
    .io_out_real(sdf_stages_4_io_out_real),
    .io_out_imag(sdf_stages_4_io_out_imag),
    .io_cntr(sdf_stages_4_io_cntr),
    .io_en(sdf_stages_4_io_en)
  );
  SDFStageRadix22_5 sdf_stages_5 ( // @[SDFChainRadix22.scala 155:25]
    .clock(sdf_stages_5_clock),
    .reset(sdf_stages_5_reset),
    .io_in_real(sdf_stages_5_io_in_real),
    .io_in_imag(sdf_stages_5_io_in_imag),
    .io_out_real(sdf_stages_5_io_out_real),
    .io_out_imag(sdf_stages_5_io_out_imag),
    .io_cntr(sdf_stages_5_io_cntr),
    .io_en(sdf_stages_5_io_en)
  );
  Queue_10 outQueue ( // @[SDFChainRadix22.scala 356:25]
    .clock(outQueue_clock),
    .reset(outQueue_reset),
    .io_enq_ready(outQueue_io_enq_ready),
    .io_enq_valid(outQueue_io_enq_valid),
    .io_enq_bits_real(outQueue_io_enq_bits_real),
    .io_enq_bits_imag(outQueue_io_enq_bits_imag),
    .io_deq_ready(outQueue_io_deq_ready),
    .io_deq_valid(outQueue_io_deq_valid),
    .io_deq_bits_real(outQueue_io_deq_bits_real),
    .io_deq_bits_imag(outQueue_io_deq_bits_imag)
  );
  assign _T_35 = regNumStages - 6'h1; // @[SDFChainRadix22.scala 69:39]
  assign _T_36 = 65'h2 << _T_35; // @[SDFChainRadix22.scala 69:23]
  assign _T_37 = io_in_ready & io_in_valid; // @[Decoupled.scala 40:37]
  assign fireLast = io_lastIn & _T_37; // @[SDFChainRadix22.scala 75:28]
  assign _T_38 = 2'h0 == state; // @[Conditional.scala 37:30]
  assign _GEN_0 = _T_37 ? 2'h1 : state; // @[SDFChainRadix22.scala 82:27]
  assign _T_41 = 2'h1 == state; // @[Conditional.scala 37:30]
  assign _GEN_1 = fireLast ? 2'h2 : state; // @[SDFChainRadix22.scala 85:23]
  assign _T_42 = 2'h2 == state; // @[Conditional.scala 37:30]
  assign _GEN_2 = io_lastOut ? 2'h0 : state; // @[SDFChainRadix22.scala 90:25]
  assign _GEN_3 = _T_42 ? _GEN_2 : state; // @[Conditional.scala 39:67]
  assign _GEN_4 = _T_41 ? _GEN_1 : _GEN_3; // @[Conditional.scala 39:67]
  assign state_next = _T_38 ? _GEN_0 : _GEN_4; // @[Conditional.scala 40:58]
  assign numPoints = _T_36[6:0]; // @[SDFChainRadix22.scala 46:23 SDFChainRadix22.scala 69:15]
  assign _T_44 = numPoints - 7'h1; // @[SDFChainRadix22.scala 104:44]
  assign _GEN_576 = {{1'd0}, cntValidOut}; // @[SDFChainRadix22.scala 104:29]
  assign _T_45 = _GEN_576 == _T_44; // @[SDFChainRadix22.scala 104:29]
  assign _T_46 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  assign pktEnd = _T_45 & _T_46; // @[SDFChainRadix22.scala 104:52]
  assign _T_47 = state_next == 2'h0; // @[SDFChainRadix22.scala 106:20]
  assign _T_50 = cnt == _T_44; // @[SDFChainRadix22.scala 109:18]
  assign _T_52 = _T_50 & _T_37; // @[SDFChainRadix22.scala 109:40]
  assign _GEN_14 = _T_52 | initialInDone; // @[SDFChainRadix22.scala 109:57]
  assign _T_54 = initialInDone & initialInDonePrev; // @[SDFChainRadix22.scala 117:41]
  assign _T_55 = fireLast & _T_54; // @[SDFChainRadix22.scala 117:23]
  assign _GEN_16 = _T_55 | lastWait; // @[SDFChainRadix22.scala 117:64]
  assign _T_57 = _T_47 & pktEnd; // @[SDFChainRadix22.scala 121:30]
  assign _T_60 = cntValidOut + 6'h1; // @[SDFChainRadix22.scala 125:32]
  assign _T_62 = lastWait & pktEnd; // @[SDFChainRadix22.scala 131:23]
  assign _GEN_20 = _T_62 | lastIndeed; // @[SDFChainRadix22.scala 131:34]
  assign _T_63 = lastIndeed & pktEnd; // @[SDFChainRadix22.scala 135:132]
  assign _T_64 = state == 2'h2; // @[SDFChainRadix22.scala 135:159]
  assign _T_65 = pktEnd & _T_64; // @[SDFChainRadix22.scala 135:150]
  assign _T_67 = 6'h6 - regNumStages; // @[SDFChainRadix22.scala 138:62]
  assign _GEN_23 = 3'h1 == _T_67[2:0] ? 6'h20 : 6'h0; // @[SDFChainRadix22.scala 138:25]
  assign _GEN_24 = 3'h2 == _T_67[2:0] ? 6'h30 : _GEN_23; // @[SDFChainRadix22.scala 138:25]
  assign _GEN_25 = 3'h3 == _T_67[2:0] ? 6'h38 : _GEN_24; // @[SDFChainRadix22.scala 138:25]
  assign _GEN_26 = 3'h4 == _T_67[2:0] ? 6'h3c : _GEN_25; // @[SDFChainRadix22.scala 138:25]
  assign _GEN_27 = 3'h5 == _T_67[2:0] ? 6'h3e : _GEN_26; // @[SDFChainRadix22.scala 138:25]
  assign cumulativeDelayWire = 3'h6 == _T_67[2:0] ? 6'h3f : _GEN_27; // @[SDFChainRadix22.scala 138:25]
  assign activeStages_0 = _T_67 <= 6'h0; // @[SDFChainRadix22.scala 146:48]
  assign activeStages_1 = _T_67 <= 6'h1; // @[SDFChainRadix22.scala 146:48]
  assign activeStages_2 = _T_67 <= 6'h2; // @[SDFChainRadix22.scala 146:48]
  assign activeStages_3 = _T_67 <= 6'h3; // @[SDFChainRadix22.scala 146:48]
  assign activeStages_4 = _T_67 <= 6'h4; // @[SDFChainRadix22.scala 146:48]
  assign activeStages_5 = _T_67 <= 6'h5; // @[SDFChainRadix22.scala 146:48]
  assign _T_95 = _T_64 & io_out_ready; // @[SDFChainRadix22.scala 164:54]
  assign enableInit = _T_37 | _T_95; // @[SDFChainRadix22.scala 164:33]
  assign _T_98 = cnt + 7'h1; // @[SDFChainRadix22.scala 170:16]
  assign _T_166 = numPoints - 7'h2; // @[SDFChainRadix22.scala 186:37]
  assign cntr_wires_0 = cnt[5:0]; // @[SDFChainRadix22.scala 48:24 SDFChainRadix22.scala 176:29]
  assign cntr_wires_1 = _T_108[5:0]; // @[SDFChainRadix22.scala 48:24 SDFChainRadix22.scala 176:29]
  assign _GEN_128 = 3'h1 == _T_35[2:0] ? cntr_wires_1 : cntr_wires_0; // @[SDFChainRadix22.scala 186:22]
  assign cntr_wires_2 = _T_118[5:0]; // @[SDFChainRadix22.scala 48:24 SDFChainRadix22.scala 176:29]
  assign _GEN_129 = 3'h2 == _T_35[2:0] ? cntr_wires_2 : _GEN_128; // @[SDFChainRadix22.scala 186:22]
  assign cntr_wires_3 = _T_128[5:0]; // @[SDFChainRadix22.scala 48:24 SDFChainRadix22.scala 176:29]
  assign _GEN_130 = 3'h3 == _T_35[2:0] ? cntr_wires_3 : _GEN_129; // @[SDFChainRadix22.scala 186:22]
  assign cntr_wires_4 = _T_138[5:0]; // @[SDFChainRadix22.scala 48:24 SDFChainRadix22.scala 176:29]
  assign _GEN_131 = 3'h4 == _T_35[2:0] ? cntr_wires_4 : _GEN_130; // @[SDFChainRadix22.scala 186:22]
  assign cntr_wires_5 = _T_148[5:0]; // @[SDFChainRadix22.scala 48:24 SDFChainRadix22.scala 176:29]
  assign _GEN_132 = 3'h5 == _T_35[2:0] ? cntr_wires_5 : _GEN_131; // @[SDFChainRadix22.scala 186:22]
  assign _GEN_577 = {{1'd0}, _GEN_132}; // @[SDFChainRadix22.scala 186:22]
  assign _T_167 = _GEN_577 == _T_166; // @[SDFChainRadix22.scala 186:22]
  assign _GEN_134 = 3'h1 == _T_35[2:0] ? enableVector_1 : enableInit; // @[SDFChainRadix22.scala 186:44]
  assign _GEN_135 = 3'h2 == _T_35[2:0] ? enableVector_2 : _GEN_134; // @[SDFChainRadix22.scala 186:44]
  assign _GEN_136 = 3'h3 == _T_35[2:0] ? enableVector_3 : _GEN_135; // @[SDFChainRadix22.scala 186:44]
  assign _GEN_137 = 3'h4 == _T_35[2:0] ? enableVector_4 : _GEN_136; // @[SDFChainRadix22.scala 186:44]
  assign _GEN_138 = 3'h5 == _T_35[2:0] ? enableVector_5 : _GEN_137; // @[SDFChainRadix22.scala 186:44]
  assign _T_168 = _T_167 & _GEN_138; // @[SDFChainRadix22.scala 186:44]
  assign _GEN_139 = _T_47 ? 1'h0 : initialOutDone; // @[SDFChainRadix22.scala 189:36]
  assign _GEN_140 = _T_168 | _GEN_139; // @[SDFChainRadix22.scala 186:60]
  assign _T_170 = numPoints == 7'h2; // @[SDFChainRadix22.scala 193:43]
  assign _T_173 = _T_171 & _T_37; // @[SDFChainRadix22.scala 193:72]
  assign _T_174 = _GEN_138 & initialOutDone; // @[SDFChainRadix22.scala 193:101]
  assign input_data_real = activeStages_0 ? $signed(io_in_bits_real) : $signed(16'sh0); // @[SDFChainRadix22.scala 211:23]
  assign input_data_imag = activeStages_0 ? $signed(io_in_bits_imag) : $signed(16'sh0); // @[SDFChainRadix22.scala 211:23]
  assign _T_184 = 6'h0 < _T_67; // @[SDFChainRadix22.scala 214:67]
  assign _T_188 = 6'h0 - _T_67; // @[SDFChainRadix22.scala 215:63]
  assign _GEN_144 = 3'h1 == _T_188[2:0] ? enableVector_1 : enableInit; // @[SDFChainRadix22.scala 216:20]
  assign _GEN_145 = 3'h2 == _T_188[2:0] ? enableVector_2 : _GEN_144; // @[SDFChainRadix22.scala 216:20]
  assign _GEN_146 = 3'h3 == _T_188[2:0] ? enableVector_3 : _GEN_145; // @[SDFChainRadix22.scala 216:20]
  assign _GEN_147 = 3'h4 == _T_188[2:0] ? enableVector_4 : _GEN_146; // @[SDFChainRadix22.scala 216:20]
  assign _GEN_148 = 3'h5 == _T_188[2:0] ? enableVector_5 : _GEN_147; // @[SDFChainRadix22.scala 216:20]
  assign _T_193 = 6'h0 - cumulativeDelayWire; // @[SDFChainRadix22.scala 217:68]
  assign _GEN_150 = 3'h1 == _T_188[2:0] ? cntr_wires_1 : cntr_wires_0; // @[SDFChainRadix22.scala 217:38]
  assign _GEN_151 = 3'h2 == _T_188[2:0] ? cntr_wires_2 : _GEN_150; // @[SDFChainRadix22.scala 217:38]
  assign _GEN_152 = 3'h3 == _T_188[2:0] ? cntr_wires_3 : _GEN_151; // @[SDFChainRadix22.scala 217:38]
  assign _GEN_153 = 3'h4 == _T_188[2:0] ? cntr_wires_4 : _GEN_152; // @[SDFChainRadix22.scala 217:38]
  assign _GEN_154 = 3'h5 == _T_188[2:0] ? cntr_wires_5 : _GEN_153; // @[SDFChainRadix22.scala 217:38]
  assign _T_199 = 6'h1 < _T_67; // @[SDFChainRadix22.scala 214:67]
  assign _T_203 = 6'h1 - _T_67; // @[SDFChainRadix22.scala 215:63]
  assign _GEN_156 = 3'h1 == _T_203[2:0] ? enableVector_1 : enableInit; // @[SDFChainRadix22.scala 216:20]
  assign _GEN_157 = 3'h2 == _T_203[2:0] ? enableVector_2 : _GEN_156; // @[SDFChainRadix22.scala 216:20]
  assign _GEN_158 = 3'h3 == _T_203[2:0] ? enableVector_3 : _GEN_157; // @[SDFChainRadix22.scala 216:20]
  assign _GEN_159 = 3'h4 == _T_203[2:0] ? enableVector_4 : _GEN_158; // @[SDFChainRadix22.scala 216:20]
  assign _GEN_160 = 3'h5 == _T_203[2:0] ? enableVector_5 : _GEN_159; // @[SDFChainRadix22.scala 216:20]
  assign _T_208 = 6'h20 - cumulativeDelayWire; // @[SDFChainRadix22.scala 217:68]
  assign _GEN_162 = 3'h1 == _T_203[2:0] ? cntr_wires_1 : cntr_wires_0; // @[SDFChainRadix22.scala 217:38]
  assign _GEN_163 = 3'h2 == _T_203[2:0] ? cntr_wires_2 : _GEN_162; // @[SDFChainRadix22.scala 217:38]
  assign _GEN_164 = 3'h3 == _T_203[2:0] ? cntr_wires_3 : _GEN_163; // @[SDFChainRadix22.scala 217:38]
  assign _GEN_165 = 3'h4 == _T_203[2:0] ? cntr_wires_4 : _GEN_164; // @[SDFChainRadix22.scala 217:38]
  assign _GEN_166 = 3'h5 == _T_203[2:0] ? cntr_wires_5 : _GEN_165; // @[SDFChainRadix22.scala 217:38]
  assign _T_210 = _GEN_166 - _T_208; // @[SDFChainRadix22.scala 217:38]
  assign _T_214 = 6'h2 < _T_67; // @[SDFChainRadix22.scala 214:67]
  assign _T_218 = 6'h2 - _T_67; // @[SDFChainRadix22.scala 215:63]
  assign _GEN_168 = 3'h1 == _T_218[2:0] ? enableVector_1 : enableInit; // @[SDFChainRadix22.scala 216:20]
  assign _GEN_169 = 3'h2 == _T_218[2:0] ? enableVector_2 : _GEN_168; // @[SDFChainRadix22.scala 216:20]
  assign _GEN_170 = 3'h3 == _T_218[2:0] ? enableVector_3 : _GEN_169; // @[SDFChainRadix22.scala 216:20]
  assign _GEN_171 = 3'h4 == _T_218[2:0] ? enableVector_4 : _GEN_170; // @[SDFChainRadix22.scala 216:20]
  assign _GEN_172 = 3'h5 == _T_218[2:0] ? enableVector_5 : _GEN_171; // @[SDFChainRadix22.scala 216:20]
  assign _T_223 = 6'h30 - cumulativeDelayWire; // @[SDFChainRadix22.scala 217:68]
  assign _GEN_174 = 3'h1 == _T_218[2:0] ? cntr_wires_1 : cntr_wires_0; // @[SDFChainRadix22.scala 217:38]
  assign _GEN_175 = 3'h2 == _T_218[2:0] ? cntr_wires_2 : _GEN_174; // @[SDFChainRadix22.scala 217:38]
  assign _GEN_176 = 3'h3 == _T_218[2:0] ? cntr_wires_3 : _GEN_175; // @[SDFChainRadix22.scala 217:38]
  assign _GEN_177 = 3'h4 == _T_218[2:0] ? cntr_wires_4 : _GEN_176; // @[SDFChainRadix22.scala 217:38]
  assign _GEN_178 = 3'h5 == _T_218[2:0] ? cntr_wires_5 : _GEN_177; // @[SDFChainRadix22.scala 217:38]
  assign _T_225 = _GEN_178 - _T_223; // @[SDFChainRadix22.scala 217:38]
  assign _T_229 = 6'h3 < _T_67; // @[SDFChainRadix22.scala 214:67]
  assign _T_233 = 6'h3 - _T_67; // @[SDFChainRadix22.scala 215:63]
  assign _GEN_180 = 3'h1 == _T_233[2:0] ? enableVector_1 : enableInit; // @[SDFChainRadix22.scala 216:20]
  assign _GEN_181 = 3'h2 == _T_233[2:0] ? enableVector_2 : _GEN_180; // @[SDFChainRadix22.scala 216:20]
  assign _GEN_182 = 3'h3 == _T_233[2:0] ? enableVector_3 : _GEN_181; // @[SDFChainRadix22.scala 216:20]
  assign _GEN_183 = 3'h4 == _T_233[2:0] ? enableVector_4 : _GEN_182; // @[SDFChainRadix22.scala 216:20]
  assign _GEN_184 = 3'h5 == _T_233[2:0] ? enableVector_5 : _GEN_183; // @[SDFChainRadix22.scala 216:20]
  assign _T_238 = 6'h38 - cumulativeDelayWire; // @[SDFChainRadix22.scala 217:68]
  assign _GEN_186 = 3'h1 == _T_233[2:0] ? cntr_wires_1 : cntr_wires_0; // @[SDFChainRadix22.scala 217:38]
  assign _GEN_187 = 3'h2 == _T_233[2:0] ? cntr_wires_2 : _GEN_186; // @[SDFChainRadix22.scala 217:38]
  assign _GEN_188 = 3'h3 == _T_233[2:0] ? cntr_wires_3 : _GEN_187; // @[SDFChainRadix22.scala 217:38]
  assign _GEN_189 = 3'h4 == _T_233[2:0] ? cntr_wires_4 : _GEN_188; // @[SDFChainRadix22.scala 217:38]
  assign _GEN_190 = 3'h5 == _T_233[2:0] ? cntr_wires_5 : _GEN_189; // @[SDFChainRadix22.scala 217:38]
  assign _T_240 = _GEN_190 - _T_238; // @[SDFChainRadix22.scala 217:38]
  assign _T_244 = 6'h4 < _T_67; // @[SDFChainRadix22.scala 214:67]
  assign _T_248 = 6'h4 - _T_67; // @[SDFChainRadix22.scala 215:63]
  assign _GEN_192 = 3'h1 == _T_248[2:0] ? enableVector_1 : enableInit; // @[SDFChainRadix22.scala 216:20]
  assign _GEN_193 = 3'h2 == _T_248[2:0] ? enableVector_2 : _GEN_192; // @[SDFChainRadix22.scala 216:20]
  assign _GEN_194 = 3'h3 == _T_248[2:0] ? enableVector_3 : _GEN_193; // @[SDFChainRadix22.scala 216:20]
  assign _GEN_195 = 3'h4 == _T_248[2:0] ? enableVector_4 : _GEN_194; // @[SDFChainRadix22.scala 216:20]
  assign _GEN_196 = 3'h5 == _T_248[2:0] ? enableVector_5 : _GEN_195; // @[SDFChainRadix22.scala 216:20]
  assign _T_253 = 6'h3c - cumulativeDelayWire; // @[SDFChainRadix22.scala 217:68]
  assign _GEN_198 = 3'h1 == _T_248[2:0] ? cntr_wires_1 : cntr_wires_0; // @[SDFChainRadix22.scala 217:38]
  assign _GEN_199 = 3'h2 == _T_248[2:0] ? cntr_wires_2 : _GEN_198; // @[SDFChainRadix22.scala 217:38]
  assign _GEN_200 = 3'h3 == _T_248[2:0] ? cntr_wires_3 : _GEN_199; // @[SDFChainRadix22.scala 217:38]
  assign _GEN_201 = 3'h4 == _T_248[2:0] ? cntr_wires_4 : _GEN_200; // @[SDFChainRadix22.scala 217:38]
  assign _GEN_202 = 3'h5 == _T_248[2:0] ? cntr_wires_5 : _GEN_201; // @[SDFChainRadix22.scala 217:38]
  assign _T_255 = _GEN_202 - _T_253; // @[SDFChainRadix22.scala 217:38]
  assign _T_259 = 6'h5 < _T_67; // @[SDFChainRadix22.scala 214:67]
  assign _T_263 = 6'h5 - _T_67; // @[SDFChainRadix22.scala 215:63]
  assign _GEN_204 = 3'h1 == _T_263[2:0] ? enableVector_1 : enableInit; // @[SDFChainRadix22.scala 216:20]
  assign _GEN_205 = 3'h2 == _T_263[2:0] ? enableVector_2 : _GEN_204; // @[SDFChainRadix22.scala 216:20]
  assign _GEN_206 = 3'h3 == _T_263[2:0] ? enableVector_3 : _GEN_205; // @[SDFChainRadix22.scala 216:20]
  assign _GEN_207 = 3'h4 == _T_263[2:0] ? enableVector_4 : _GEN_206; // @[SDFChainRadix22.scala 216:20]
  assign _GEN_208 = 3'h5 == _T_263[2:0] ? enableVector_5 : _GEN_207; // @[SDFChainRadix22.scala 216:20]
  assign _T_268 = 6'h3e - cumulativeDelayWire; // @[SDFChainRadix22.scala 217:68]
  assign _GEN_210 = 3'h1 == _T_263[2:0] ? cntr_wires_1 : cntr_wires_0; // @[SDFChainRadix22.scala 217:38]
  assign _GEN_211 = 3'h2 == _T_263[2:0] ? cntr_wires_2 : _GEN_210; // @[SDFChainRadix22.scala 217:38]
  assign _GEN_212 = 3'h3 == _T_263[2:0] ? cntr_wires_3 : _GEN_211; // @[SDFChainRadix22.scala 217:38]
  assign _GEN_213 = 3'h4 == _T_263[2:0] ? cntr_wires_4 : _GEN_212; // @[SDFChainRadix22.scala 217:38]
  assign _GEN_214 = 3'h5 == _T_263[2:0] ? cntr_wires_5 : _GEN_213; // @[SDFChainRadix22.scala 217:38]
  assign _T_270 = _GEN_214 - _T_268; // @[SDFChainRadix22.scala 217:38]
  assign _T_277 = 6'h0 == _T_67; // @[SDFChainRadix22.scala 234:23]
  assign _GEN_215 = _T_277 ? $signed(io_in_bits_imag) : $signed(input_data_imag); // @[SDFChainRadix22.scala 234:55]
  assign _GEN_216 = _T_277 ? $signed(io_in_bits_real) : $signed(input_data_real); // @[SDFChainRadix22.scala 234:55]
  assign _T_278 = sdf_stages_0_io_cntr < 6'h20; // @[SDFChainRadix22.scala 320:98]
  assign _T_280 = sdf_stages_0_io_cntr < 6'h10; // @[SDFChainRadix22.scala 320:135]
  assign _T_281 = _T_280 ? 1'h0 : 1'h1; // @[SDFChainRadix22.scala 320:122]
  assign _T_289 = 16'sh0 - $signed(sdf_stages_0_io_out_real); // @[FixedPointTypeClass.scala 39:43]
  assign _T_286_real = sdf_stages_0_io_out_imag; // @[SDFChainRadix22.scala 322:32 SDFChainRadix22.scala 325:29]
  assign _T_307 = 6'h1 == _T_67; // @[SDFChainRadix22.scala 234:23]
  assign _GEN_226 = _T_307 ? $signed(io_in_bits_imag) : $signed(outputWires_0_imag); // @[SDFChainRadix22.scala 234:55]
  assign _GEN_227 = _T_307 ? $signed(io_in_bits_real) : $signed(outputWires_0_real); // @[SDFChainRadix22.scala 234:55]
  assign _T_475 = _GEN_166 + 6'h1; // @[SDFChainRadix22.scala 276:83]
  assign _T_479 = _T_475 - _T_223; // @[SDFChainRadix22.scala 276:89]
  assign _GEN_266 = 6'h11 == _T_481 ? 5'h2 : 5'h0; // @[Reg.scala 16:23]
  assign _GEN_267 = 6'h12 == _T_481 ? 5'h4 : _GEN_266; // @[Reg.scala 16:23]
  assign _GEN_268 = 6'h13 == _T_481 ? 5'h6 : _GEN_267; // @[Reg.scala 16:23]
  assign _GEN_269 = 6'h14 == _T_481 ? 5'h8 : _GEN_268; // @[Reg.scala 16:23]
  assign _GEN_270 = 6'h15 == _T_481 ? 5'ha : _GEN_269; // @[Reg.scala 16:23]
  assign _GEN_271 = 6'h16 == _T_481 ? 5'hc : _GEN_270; // @[Reg.scala 16:23]
  assign _GEN_272 = 6'h17 == _T_481 ? 5'he : _GEN_271; // @[Reg.scala 16:23]
  assign _GEN_273 = 6'h18 == _T_481 ? 5'h10 : _GEN_272; // @[Reg.scala 16:23]
  assign _GEN_274 = 6'h19 == _T_481 ? 5'h11 : _GEN_273; // @[Reg.scala 16:23]
  assign _GEN_275 = 6'h1a == _T_481 ? 5'h12 : _GEN_274; // @[Reg.scala 16:23]
  assign _GEN_276 = 6'h1b == _T_481 ? 5'h14 : _GEN_275; // @[Reg.scala 16:23]
  assign _GEN_277 = 6'h1c == _T_481 ? 5'h15 : _GEN_276; // @[Reg.scala 16:23]
  assign _GEN_278 = 6'h1d == _T_481 ? 5'h16 : _GEN_277; // @[Reg.scala 16:23]
  assign _GEN_279 = 6'h1e == _T_481 ? 5'h18 : _GEN_278; // @[Reg.scala 16:23]
  assign _GEN_280 = 6'h1f == _T_481 ? 5'h19 : _GEN_279; // @[Reg.scala 16:23]
  assign _GEN_281 = 6'h20 == _T_481 ? 5'h0 : _GEN_280; // @[Reg.scala 16:23]
  assign _GEN_282 = 6'h21 == _T_481 ? 5'h1 : _GEN_281; // @[Reg.scala 16:23]
  assign _GEN_283 = 6'h22 == _T_481 ? 5'h2 : _GEN_282; // @[Reg.scala 16:23]
  assign _GEN_284 = 6'h23 == _T_481 ? 5'h3 : _GEN_283; // @[Reg.scala 16:23]
  assign _GEN_285 = 6'h24 == _T_481 ? 5'h4 : _GEN_284; // @[Reg.scala 16:23]
  assign _GEN_286 = 6'h25 == _T_481 ? 5'h5 : _GEN_285; // @[Reg.scala 16:23]
  assign _GEN_287 = 6'h26 == _T_481 ? 5'h6 : _GEN_286; // @[Reg.scala 16:23]
  assign _GEN_288 = 6'h27 == _T_481 ? 5'h7 : _GEN_287; // @[Reg.scala 16:23]
  assign _GEN_289 = 6'h28 == _T_481 ? 5'h8 : _GEN_288; // @[Reg.scala 16:23]
  assign _GEN_290 = 6'h29 == _T_481 ? 5'h9 : _GEN_289; // @[Reg.scala 16:23]
  assign _GEN_291 = 6'h2a == _T_481 ? 5'ha : _GEN_290; // @[Reg.scala 16:23]
  assign _GEN_292 = 6'h2b == _T_481 ? 5'hb : _GEN_291; // @[Reg.scala 16:23]
  assign _GEN_293 = 6'h2c == _T_481 ? 5'hc : _GEN_292; // @[Reg.scala 16:23]
  assign _GEN_294 = 6'h2d == _T_481 ? 5'hd : _GEN_293; // @[Reg.scala 16:23]
  assign _GEN_295 = 6'h2e == _T_481 ? 5'he : _GEN_294; // @[Reg.scala 16:23]
  assign _GEN_296 = 6'h2f == _T_481 ? 5'hf : _GEN_295; // @[Reg.scala 16:23]
  assign _GEN_297 = 6'h30 == _T_481 ? 5'h0 : _GEN_296; // @[Reg.scala 16:23]
  assign _GEN_298 = 6'h31 == _T_481 ? 5'h3 : _GEN_297; // @[Reg.scala 16:23]
  assign _GEN_299 = 6'h32 == _T_481 ? 5'h6 : _GEN_298; // @[Reg.scala 16:23]
  assign _GEN_300 = 6'h33 == _T_481 ? 5'h9 : _GEN_299; // @[Reg.scala 16:23]
  assign _GEN_301 = 6'h34 == _T_481 ? 5'hc : _GEN_300; // @[Reg.scala 16:23]
  assign _GEN_302 = 6'h35 == _T_481 ? 5'hf : _GEN_301; // @[Reg.scala 16:23]
  assign _GEN_303 = 6'h36 == _T_481 ? 5'h11 : _GEN_302; // @[Reg.scala 16:23]
  assign _GEN_304 = 6'h37 == _T_481 ? 5'h13 : _GEN_303; // @[Reg.scala 16:23]
  assign _GEN_305 = 6'h38 == _T_481 ? 5'h15 : _GEN_304; // @[Reg.scala 16:23]
  assign _GEN_306 = 6'h39 == _T_481 ? 5'h17 : _GEN_305; // @[Reg.scala 16:23]
  assign _GEN_307 = 6'h3a == _T_481 ? 5'h19 : _GEN_306; // @[Reg.scala 16:23]
  assign _GEN_308 = 6'h3b == _T_481 ? 5'h1a : _GEN_307; // @[Reg.scala 16:23]
  assign _GEN_309 = 6'h3c == _T_481 ? 5'h1b : _GEN_308; // @[Reg.scala 16:23]
  assign _GEN_310 = 6'h3d == _T_481 ? 5'h1c : _GEN_309; // @[Reg.scala 16:23]
  assign _GEN_311 = 6'h3e == _T_481 ? 5'h1d : _GEN_310; // @[Reg.scala 16:23]
  assign _GEN_312 = 6'h3f == _T_481 ? 5'h1e : _GEN_311; // @[Reg.scala 16:23]
  assign _GEN_578 = {{1{_T_490[15]}},_T_490}; // @[FixedPointTypeClass.scala 211:35]
  assign _GEN_579 = {$signed(_T_500), 2'h0}; // @[FixedPointTypeClass.scala 20:58]
  assign _T_503 = $signed(_GEN_579) + 35'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign _T_504 = _T_503[34:1]; // @[FixedPointTypeClass.scala 176:41]
  assign _GEN_580 = {{1{_T_492[15]}},_T_492}; // @[FixedPointTypeClass.scala 211:35]
  assign _GEN_581 = {$signed(_T_506), 2'h0}; // @[FixedPointTypeClass.scala 20:58]
  assign _T_509 = $signed(_GEN_581) + 35'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign _T_510 = _T_509[34:1]; // @[FixedPointTypeClass.scala 176:41]
  assign _GEN_582 = {{1{_T_491[15]}},_T_491}; // @[FixedPointTypeClass.scala 211:35]
  assign _GEN_583 = {$signed(_T_512), 2'h0}; // @[FixedPointTypeClass.scala 20:58]
  assign _T_515 = $signed(_GEN_583) + 35'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign _T_516 = _T_515[34:1]; // @[FixedPointTypeClass.scala 176:41]
  assign _T_526 = $signed(_T_518) + 35'sh4000; // @[FixedPointTypeClass.scala 20:58]
  assign _T_527 = _T_526[34:15]; // @[FixedPointTypeClass.scala 176:41]
  assign _T_530 = $signed(_T_520) + 35'sh4000; // @[FixedPointTypeClass.scala 20:58]
  assign _T_531 = _T_530[34:15]; // @[FixedPointTypeClass.scala 176:41]
  assign _T_540 = 6'h2 == _T_67; // @[SDFChainRadix22.scala 234:23]
  assign outputWires_1_imag = _T_531[15:0]; // @[SDFChainRadix22.scala 286:27 SDFChainRadix22.scala 306:19]
  assign _GEN_450 = _T_540 ? $signed(io_in_bits_imag) : $signed(outputWires_1_imag); // @[SDFChainRadix22.scala 234:55]
  assign outputWires_1_real = _T_527[15:0]; // @[SDFChainRadix22.scala 286:27 SDFChainRadix22.scala 306:19]
  assign _GEN_451 = _T_540 ? $signed(io_in_bits_real) : $signed(outputWires_1_real); // @[SDFChainRadix22.scala 234:55]
  assign _T_541 = sdf_stages_2_io_cntr < 6'h8; // @[SDFChainRadix22.scala 320:98]
  assign _T_543 = sdf_stages_2_io_cntr < 6'h4; // @[SDFChainRadix22.scala 320:135]
  assign _T_544 = _T_543 ? 1'h0 : 1'h1; // @[SDFChainRadix22.scala 320:122]
  assign _T_552 = 16'sh0 - $signed(sdf_stages_2_io_out_real); // @[FixedPointTypeClass.scala 39:43]
  assign _T_549_real = sdf_stages_2_io_out_imag; // @[SDFChainRadix22.scala 322:32 SDFChainRadix22.scala 325:29]
  assign _T_570 = 6'h3 == _T_67; // @[SDFChainRadix22.scala 234:23]
  assign _GEN_461 = _T_570 ? $signed(io_in_bits_imag) : $signed(outputWires_2_imag); // @[SDFChainRadix22.scala 234:55]
  assign _GEN_462 = _T_570 ? $signed(io_in_bits_real) : $signed(outputWires_2_real); // @[SDFChainRadix22.scala 234:55]
  assign _T_618 = _GEN_190 + 6'h1; // @[SDFChainRadix22.scala 276:83]
  assign _T_622 = _T_618 - _T_253; // @[SDFChainRadix22.scala 276:89]
  assign _GEN_489 = 4'h5 == _T_624[3:0] ? 3'h2 : 3'h0; // @[Reg.scala 16:23]
  assign _GEN_490 = 4'h6 == _T_624[3:0] ? 3'h4 : _GEN_489; // @[Reg.scala 16:23]
  assign _GEN_491 = 4'h7 == _T_624[3:0] ? 3'h5 : _GEN_490; // @[Reg.scala 16:23]
  assign _GEN_492 = 4'h8 == _T_624[3:0] ? 3'h0 : _GEN_491; // @[Reg.scala 16:23]
  assign _GEN_493 = 4'h9 == _T_624[3:0] ? 3'h1 : _GEN_492; // @[Reg.scala 16:23]
  assign _GEN_494 = 4'ha == _T_624[3:0] ? 3'h2 : _GEN_493; // @[Reg.scala 16:23]
  assign _GEN_495 = 4'hb == _T_624[3:0] ? 3'h3 : _GEN_494; // @[Reg.scala 16:23]
  assign _GEN_496 = 4'hc == _T_624[3:0] ? 3'h0 : _GEN_495; // @[Reg.scala 16:23]
  assign _GEN_497 = 4'hd == _T_624[3:0] ? 3'h3 : _GEN_496; // @[Reg.scala 16:23]
  assign _GEN_498 = 4'he == _T_624[3:0] ? 3'h5 : _GEN_497; // @[Reg.scala 16:23]
  assign _GEN_499 = 4'hf == _T_624[3:0] ? 3'h6 : _GEN_498; // @[Reg.scala 16:23]
  assign _GEN_586 = {{1{_T_634[15]}},_T_634}; // @[FixedPointTypeClass.scala 211:35]
  assign _GEN_587 = {$signed(_T_644), 2'h0}; // @[FixedPointTypeClass.scala 20:58]
  assign _T_647 = $signed(_GEN_587) + 35'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign _T_648 = _T_647[34:1]; // @[FixedPointTypeClass.scala 176:41]
  assign _GEN_588 = {{1{_T_636[15]}},_T_636}; // @[FixedPointTypeClass.scala 211:35]
  assign _GEN_589 = {$signed(_T_650), 2'h0}; // @[FixedPointTypeClass.scala 20:58]
  assign _T_653 = $signed(_GEN_589) + 35'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign _T_654 = _T_653[34:1]; // @[FixedPointTypeClass.scala 176:41]
  assign _GEN_590 = {{1{_T_635[15]}},_T_635}; // @[FixedPointTypeClass.scala 211:35]
  assign _GEN_591 = {$signed(_T_656), 2'h0}; // @[FixedPointTypeClass.scala 20:58]
  assign _T_659 = $signed(_GEN_591) + 35'sh1; // @[FixedPointTypeClass.scala 20:58]
  assign _T_660 = _T_659[34:1]; // @[FixedPointTypeClass.scala 176:41]
  assign _T_670 = $signed(_T_662) + 35'sh4000; // @[FixedPointTypeClass.scala 20:58]
  assign _T_671 = _T_670[34:15]; // @[FixedPointTypeClass.scala 176:41]
  assign _T_674 = $signed(_T_664) + 35'sh4000; // @[FixedPointTypeClass.scala 20:58]
  assign _T_675 = _T_674[34:15]; // @[FixedPointTypeClass.scala 176:41]
  assign _T_684 = 6'h4 == _T_67; // @[SDFChainRadix22.scala 234:23]
  assign outputWires_3_imag = _T_675[15:0]; // @[SDFChainRadix22.scala 286:27 SDFChainRadix22.scala 306:19]
  assign _GEN_541 = _T_684 ? $signed(io_in_bits_imag) : $signed(outputWires_3_imag); // @[SDFChainRadix22.scala 234:55]
  assign outputWires_3_real = _T_671[15:0]; // @[SDFChainRadix22.scala 286:27 SDFChainRadix22.scala 306:19]
  assign _GEN_542 = _T_684 ? $signed(io_in_bits_real) : $signed(outputWires_3_real); // @[SDFChainRadix22.scala 234:55]
  assign _T_685 = sdf_stages_4_io_cntr < 6'h2; // @[SDFChainRadix22.scala 320:98]
  assign _T_687 = sdf_stages_4_io_cntr < 6'h1; // @[SDFChainRadix22.scala 320:135]
  assign _T_688 = _T_687 ? 1'h0 : 1'h1; // @[SDFChainRadix22.scala 320:122]
  assign _T_696 = 16'sh0 - $signed(sdf_stages_4_io_out_real); // @[FixedPointTypeClass.scala 39:43]
  assign _T_693_real = sdf_stages_4_io_out_imag; // @[SDFChainRadix22.scala 322:32 SDFChainRadix22.scala 325:29]
  assign _T_714 = 6'h5 == _T_67; // @[SDFChainRadix22.scala 234:23]
  assign _GEN_552 = _T_714 ? $signed(io_in_bits_imag) : $signed(outputWires_4_imag); // @[SDFChainRadix22.scala 234:55]
  assign _GEN_553 = _T_714 ? $signed(io_in_bits_real) : $signed(outputWires_4_real); // @[SDFChainRadix22.scala 234:55]
  assign _T_728 = ~initialOutDone; // @[SDFChainRadix22.scala 361:33]
  assign _T_733 = state != 2'h2; // @[SDFChainRadix22.scala 361:127]
  assign _T_734 = io_out_ready & _T_733; // @[SDFChainRadix22.scala 361:117]
  assign _GEN_594 = {$signed(outQueue_io_deq_bits_imag), 14'h0}; // @[SDFChainRadix22.scala 375:33]
  assign _GEN_574 = {{2{_GEN_594[29]}},_GEN_594}; // @[SDFChainRadix22.scala 375:33]
  assign _GEN_595 = {$signed(outQueue_io_deq_bits_real), 14'h0}; // @[SDFChainRadix22.scala 375:33]
  assign _GEN_575 = {{2{_GEN_595[29]}},_GEN_595}; // @[SDFChainRadix22.scala 375:33]
  assign _GEN_596 = _GEN_575[31:14]; // @[SDFChainRadix22.scala 59:26 SDFChainRadix22.scala 376:20 SDFChainRadix22.scala 379:25]
  assign _GEN_598 = _GEN_574[31:14]; // @[SDFChainRadix22.scala 59:26 SDFChainRadix22.scala 376:20 SDFChainRadix22.scala 380:25]
  assign io_in_ready = _T_732 | _T_734; // @[SDFChainRadix22.scala 361:15]
  assign io_out_valid = outQueue_io_deq_valid; // @[SDFChainRadix22.scala 383:18]
  assign io_out_bits_real = _GEN_596[15:0]; // @[SDFChainRadix22.scala 382:17]
  assign io_out_bits_imag = _GEN_598[15:0]; // @[SDFChainRadix22.scala 382:17]
  assign io_lastOut = lastWait ? _T_63 : _T_65; // @[SDFChainRadix22.scala 389:14]
  assign io_busy = state == 2'h2; // @[SDFChainRadix22.scala 390:11]
  assign sdf_stages_0_clock = clock;
  assign sdf_stages_0_reset = reset;
  assign sdf_stages_0_io_in_real = activeStages_0 ? $signed(_GEN_216) : $signed(16'sh0); // @[SDFChainRadix22.scala 245:21 SDFChainRadix22.scala 248:21]
  assign sdf_stages_0_io_in_imag = activeStages_0 ? $signed(_GEN_215) : $signed(16'sh0); // @[SDFChainRadix22.scala 245:21 SDFChainRadix22.scala 248:21]
  assign sdf_stages_0_io_cntr = _GEN_154 - _T_193; // @[SDFChainRadix22.scala 217:16]
  assign sdf_stages_0_io_en = _T_184 ? 1'h0 : _GEN_148; // @[SDFChainRadix22.scala 216:14]
  assign sdf_stages_1_clock = clock;
  assign sdf_stages_1_reset = reset;
  assign sdf_stages_1_io_in_real = activeStages_1 ? $signed(_GEN_227) : $signed(16'sh0); // @[SDFChainRadix22.scala 245:21 SDFChainRadix22.scala 248:21]
  assign sdf_stages_1_io_in_imag = activeStages_1 ? $signed(_GEN_226) : $signed(16'sh0); // @[SDFChainRadix22.scala 245:21 SDFChainRadix22.scala 248:21]
  assign sdf_stages_1_io_cntr = {{1'd0}, _T_210[4:0]}; // @[SDFChainRadix22.scala 217:16]
  assign sdf_stages_1_io_en = _T_199 ? 1'h0 : _GEN_160; // @[SDFChainRadix22.scala 216:14]
  assign sdf_stages_2_clock = clock;
  assign sdf_stages_2_reset = reset;
  assign sdf_stages_2_io_in_real = activeStages_2 ? $signed(_GEN_451) : $signed(16'sh0); // @[SDFChainRadix22.scala 245:21 SDFChainRadix22.scala 248:21]
  assign sdf_stages_2_io_in_imag = activeStages_2 ? $signed(_GEN_450) : $signed(16'sh0); // @[SDFChainRadix22.scala 245:21 SDFChainRadix22.scala 248:21]
  assign sdf_stages_2_io_cntr = {{2'd0}, _T_225[3:0]}; // @[SDFChainRadix22.scala 217:16]
  assign sdf_stages_2_io_en = _T_214 ? 1'h0 : _GEN_172; // @[SDFChainRadix22.scala 216:14]
  assign sdf_stages_3_clock = clock;
  assign sdf_stages_3_reset = reset;
  assign sdf_stages_3_io_in_real = activeStages_3 ? $signed(_GEN_462) : $signed(16'sh0); // @[SDFChainRadix22.scala 245:21 SDFChainRadix22.scala 248:21]
  assign sdf_stages_3_io_in_imag = activeStages_3 ? $signed(_GEN_461) : $signed(16'sh0); // @[SDFChainRadix22.scala 245:21 SDFChainRadix22.scala 248:21]
  assign sdf_stages_3_io_cntr = {{3'd0}, _T_240[2:0]}; // @[SDFChainRadix22.scala 217:16]
  assign sdf_stages_3_io_en = _T_229 ? 1'h0 : _GEN_184; // @[SDFChainRadix22.scala 216:14]
  assign sdf_stages_4_clock = clock;
  assign sdf_stages_4_reset = reset;
  assign sdf_stages_4_io_in_real = activeStages_4 ? $signed(_GEN_542) : $signed(16'sh0); // @[SDFChainRadix22.scala 245:21 SDFChainRadix22.scala 248:21]
  assign sdf_stages_4_io_in_imag = activeStages_4 ? $signed(_GEN_541) : $signed(16'sh0); // @[SDFChainRadix22.scala 245:21 SDFChainRadix22.scala 248:21]
  assign sdf_stages_4_io_cntr = {{4'd0}, _T_255[1:0]}; // @[SDFChainRadix22.scala 217:16]
  assign sdf_stages_4_io_en = _T_244 ? 1'h0 : _GEN_196; // @[SDFChainRadix22.scala 216:14]
  assign sdf_stages_5_clock = clock;
  assign sdf_stages_5_reset = reset;
  assign sdf_stages_5_io_in_real = activeStages_5 ? $signed(_GEN_553) : $signed(16'sh0); // @[SDFChainRadix22.scala 245:21 SDFChainRadix22.scala 248:21]
  assign sdf_stages_5_io_in_imag = activeStages_5 ? $signed(_GEN_552) : $signed(16'sh0); // @[SDFChainRadix22.scala 245:21 SDFChainRadix22.scala 248:21]
  assign sdf_stages_5_io_cntr = {{5'd0}, _T_270[0]}; // @[SDFChainRadix22.scala 217:16]
  assign sdf_stages_5_io_en = _T_259 ? 1'h0 : _GEN_208; // @[SDFChainRadix22.scala 216:14]
  assign outQueue_clock = clock;
  assign outQueue_reset = reset;
  assign outQueue_io_enq_valid = outValid; // @[SDFChainRadix22.scala 358:25]
  assign outQueue_io_enq_bits_real = outputWires_5_real; // @[SDFChainRadix22.scala 357:24]
  assign outQueue_io_enq_bits_imag = outputWires_5_imag; // @[SDFChainRadix22.scala 357:24]
  assign outQueue_io_deq_ready = io_out_ready; // @[SDFChainRadix22.scala 359:25]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regNumStages = _RAND_0[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  state = _RAND_1[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  initialOutDone = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  cnt = _RAND_3[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  cntValidOut = _RAND_4[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  lastWait = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  lastIndeed = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  initialInDone = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  initialInDonePrev = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_100 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_101 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_102 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  enableVector_1 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_105 = _RAND_13[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_106 = _RAND_14[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_107 = _RAND_15[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_108 = _RAND_16[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_110 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_111 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_112 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  enableVector_2 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_115 = _RAND_21[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_116 = _RAND_22[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_117 = _RAND_23[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_118 = _RAND_24[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_120 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_121 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T_122 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  enableVector_3 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_125 = _RAND_29[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_126 = _RAND_30[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T_127 = _RAND_31[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _T_128 = _RAND_32[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _T_130 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _T_131 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _T_132 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  enableVector_4 = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _T_135 = _RAND_37[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _T_136 = _RAND_38[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _T_137 = _RAND_39[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _T_138 = _RAND_40[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  _T_140 = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  _T_141 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  _T_142 = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  enableVector_5 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  _T_145 = _RAND_45[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  _T_146 = _RAND_46[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  _T_147 = _RAND_47[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  _T_148 = _RAND_48[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  _T_171 = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  _T_283 = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  _T_295_real = _RAND_51[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  _T_295_imag = _RAND_52[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  _T_298_real = _RAND_53[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  _T_298_imag = _RAND_54[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  outputWires_0_real = _RAND_55[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  outputWires_0_imag = _RAND_56[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  _T_481 = _RAND_57[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  twiddles_1_real = _RAND_58[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  twiddles_1_imag = _RAND_59[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  _T_490 = _RAND_60[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  _T_491 = _RAND_61[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  _T_492 = _RAND_62[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  _T_494 = _RAND_63[16:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  _T_496 = _RAND_64[16:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  _T_498 = _RAND_65[16:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {2{`RANDOM}};
  _T_500 = _RAND_66[32:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {2{`RANDOM}};
  _T_506 = _RAND_67[32:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {2{`RANDOM}};
  _T_512 = _RAND_68[32:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {2{`RANDOM}};
  _T_518 = _RAND_69[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {2{`RANDOM}};
  _T_520 = _RAND_70[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  _T_546 = _RAND_71[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  _T_558_real = _RAND_72[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  _T_558_imag = _RAND_73[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  _T_561_real = _RAND_74[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  _T_561_imag = _RAND_75[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  outputWires_2_real = _RAND_76[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  outputWires_2_imag = _RAND_77[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  _T_624 = _RAND_78[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  twiddles_3_real = _RAND_79[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  twiddles_3_imag = _RAND_80[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  _T_634 = _RAND_81[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  _T_635 = _RAND_82[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  _T_636 = _RAND_83[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  _T_638 = _RAND_84[16:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  _T_640 = _RAND_85[16:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  _T_642 = _RAND_86[16:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {2{`RANDOM}};
  _T_644 = _RAND_87[32:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {2{`RANDOM}};
  _T_650 = _RAND_88[32:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {2{`RANDOM}};
  _T_656 = _RAND_89[32:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {2{`RANDOM}};
  _T_662 = _RAND_90[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {2{`RANDOM}};
  _T_664 = _RAND_91[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  _T_690 = _RAND_92[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  _T_702_real = _RAND_93[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  _T_702_imag = _RAND_94[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  _T_705_real = _RAND_95[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  _T_705_imag = _RAND_96[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  outputWires_4_real = _RAND_97[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  outputWires_4_imag = _RAND_98[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  _T_717_real = _RAND_99[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  _T_717_imag = _RAND_100[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  _T_720_real = _RAND_101[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  _T_720_imag = _RAND_102[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  outputWires_5_real = _RAND_103[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  outputWires_5_imag = _RAND_104[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  _T_725 = _RAND_105[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  _T_726 = _RAND_106[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  _T_727 = _RAND_107[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  outValid = _RAND_108[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  _T_729 = _RAND_109[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  _T_730 = _RAND_110[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  _T_731 = _RAND_111[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  _T_732 = _RAND_112[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      regNumStages <= 6'h6;
    end else if (_T_38) begin
      regNumStages <= io_fftSize;
    end
    if (reset) begin
      state <= 2'h0;
    end else if (_T_38) begin
      if (_T_37) begin
        state <= 2'h1;
      end
    end else if (_T_41) begin
      if (fireLast) begin
        state <= 2'h2;
      end
    end else if (_T_42) begin
      if (io_lastOut) begin
        state <= 2'h0;
      end
    end
    if (reset) begin
      initialOutDone <= 1'h0;
    end else begin
      initialOutDone <= _GEN_140;
    end
    if (reset) begin
      cnt <= 7'h0;
    end else if (_T_47) begin
      cnt <= 7'h0;
    end else if (enableInit) begin
      cnt <= _T_98;
    end
    if (reset) begin
      cntValidOut <= 6'h0;
    end else if (_T_57) begin
      cntValidOut <= 6'h0;
    end else if (_T_46) begin
      cntValidOut <= _T_60;
    end
    if (reset) begin
      lastWait <= 1'h0;
    end else if (_T_47) begin
      lastWait <= 1'h0;
    end else begin
      lastWait <= _GEN_16;
    end
    if (reset) begin
      lastIndeed <= 1'h0;
    end else if (_T_47) begin
      lastIndeed <= 1'h0;
    end else begin
      lastIndeed <= _GEN_20;
    end
    if (reset) begin
      initialInDone <= 1'h0;
    end else if (_T_47) begin
      initialInDone <= 1'h0;
    end else begin
      initialInDone <= _GEN_14;
    end
    if (reset) begin
      initialInDonePrev <= 1'h0;
    end else begin
      initialInDonePrev <= initialInDone;
    end
    if (reset) begin
      _T_100 <= 1'h0;
    end else if (_T_47) begin
      _T_100 <= 1'h0;
    end else begin
      _T_100 <= enableInit;
    end
    if (reset) begin
      _T_101 <= 1'h0;
    end else if (_T_47) begin
      _T_101 <= 1'h0;
    end else begin
      _T_101 <= _T_100;
    end
    if (reset) begin
      _T_102 <= 1'h0;
    end else if (_T_47) begin
      _T_102 <= 1'h0;
    end else begin
      _T_102 <= _T_101;
    end
    if (reset) begin
      enableVector_1 <= 1'h0;
    end else if (_T_47) begin
      enableVector_1 <= 1'h0;
    end else begin
      enableVector_1 <= _T_102;
    end
    if (reset) begin
      _T_105 <= 7'h0;
    end else if (_T_47) begin
      _T_105 <= 7'h0;
    end else begin
      _T_105 <= cnt;
    end
    if (reset) begin
      _T_106 <= 7'h0;
    end else if (_T_47) begin
      _T_106 <= 7'h0;
    end else begin
      _T_106 <= _T_105;
    end
    if (reset) begin
      _T_107 <= 7'h0;
    end else if (_T_47) begin
      _T_107 <= 7'h0;
    end else begin
      _T_107 <= _T_106;
    end
    if (reset) begin
      _T_108 <= 7'h0;
    end else if (_T_47) begin
      _T_108 <= 7'h0;
    end else begin
      _T_108 <= _T_107;
    end
    if (reset) begin
      _T_110 <= 1'h0;
    end else if (_T_47) begin
      _T_110 <= 1'h0;
    end else begin
      _T_110 <= enableVector_1;
    end
    if (reset) begin
      _T_111 <= 1'h0;
    end else if (_T_47) begin
      _T_111 <= 1'h0;
    end else begin
      _T_111 <= _T_110;
    end
    if (reset) begin
      _T_112 <= 1'h0;
    end else if (_T_47) begin
      _T_112 <= 1'h0;
    end else begin
      _T_112 <= _T_111;
    end
    if (reset) begin
      enableVector_2 <= 1'h0;
    end else if (_T_47) begin
      enableVector_2 <= 1'h0;
    end else begin
      enableVector_2 <= _T_112;
    end
    if (reset) begin
      _T_115 <= 7'h0;
    end else if (_T_47) begin
      _T_115 <= 7'h0;
    end else begin
      _T_115 <= _T_108;
    end
    if (reset) begin
      _T_116 <= 7'h0;
    end else if (_T_47) begin
      _T_116 <= 7'h0;
    end else begin
      _T_116 <= _T_115;
    end
    if (reset) begin
      _T_117 <= 7'h0;
    end else if (_T_47) begin
      _T_117 <= 7'h0;
    end else begin
      _T_117 <= _T_116;
    end
    if (reset) begin
      _T_118 <= 7'h0;
    end else if (_T_47) begin
      _T_118 <= 7'h0;
    end else begin
      _T_118 <= _T_117;
    end
    if (reset) begin
      _T_120 <= 1'h0;
    end else if (_T_47) begin
      _T_120 <= 1'h0;
    end else begin
      _T_120 <= enableVector_2;
    end
    if (reset) begin
      _T_121 <= 1'h0;
    end else if (_T_47) begin
      _T_121 <= 1'h0;
    end else begin
      _T_121 <= _T_120;
    end
    if (reset) begin
      _T_122 <= 1'h0;
    end else if (_T_47) begin
      _T_122 <= 1'h0;
    end else begin
      _T_122 <= _T_121;
    end
    if (reset) begin
      enableVector_3 <= 1'h0;
    end else if (_T_47) begin
      enableVector_3 <= 1'h0;
    end else begin
      enableVector_3 <= _T_122;
    end
    if (reset) begin
      _T_125 <= 7'h0;
    end else if (_T_47) begin
      _T_125 <= 7'h0;
    end else begin
      _T_125 <= _T_118;
    end
    if (reset) begin
      _T_126 <= 7'h0;
    end else if (_T_47) begin
      _T_126 <= 7'h0;
    end else begin
      _T_126 <= _T_125;
    end
    if (reset) begin
      _T_127 <= 7'h0;
    end else if (_T_47) begin
      _T_127 <= 7'h0;
    end else begin
      _T_127 <= _T_126;
    end
    if (reset) begin
      _T_128 <= 7'h0;
    end else if (_T_47) begin
      _T_128 <= 7'h0;
    end else begin
      _T_128 <= _T_127;
    end
    if (reset) begin
      _T_130 <= 1'h0;
    end else if (_T_47) begin
      _T_130 <= 1'h0;
    end else begin
      _T_130 <= enableVector_3;
    end
    if (reset) begin
      _T_131 <= 1'h0;
    end else if (_T_47) begin
      _T_131 <= 1'h0;
    end else begin
      _T_131 <= _T_130;
    end
    if (reset) begin
      _T_132 <= 1'h0;
    end else if (_T_47) begin
      _T_132 <= 1'h0;
    end else begin
      _T_132 <= _T_131;
    end
    if (reset) begin
      enableVector_4 <= 1'h0;
    end else if (_T_47) begin
      enableVector_4 <= 1'h0;
    end else begin
      enableVector_4 <= _T_132;
    end
    if (reset) begin
      _T_135 <= 7'h0;
    end else if (_T_47) begin
      _T_135 <= 7'h0;
    end else begin
      _T_135 <= _T_128;
    end
    if (reset) begin
      _T_136 <= 7'h0;
    end else if (_T_47) begin
      _T_136 <= 7'h0;
    end else begin
      _T_136 <= _T_135;
    end
    if (reset) begin
      _T_137 <= 7'h0;
    end else if (_T_47) begin
      _T_137 <= 7'h0;
    end else begin
      _T_137 <= _T_136;
    end
    if (reset) begin
      _T_138 <= 7'h0;
    end else if (_T_47) begin
      _T_138 <= 7'h0;
    end else begin
      _T_138 <= _T_137;
    end
    if (reset) begin
      _T_140 <= 1'h0;
    end else if (_T_47) begin
      _T_140 <= 1'h0;
    end else begin
      _T_140 <= enableVector_4;
    end
    if (reset) begin
      _T_141 <= 1'h0;
    end else if (_T_47) begin
      _T_141 <= 1'h0;
    end else begin
      _T_141 <= _T_140;
    end
    if (reset) begin
      _T_142 <= 1'h0;
    end else if (_T_47) begin
      _T_142 <= 1'h0;
    end else begin
      _T_142 <= _T_141;
    end
    if (reset) begin
      enableVector_5 <= 1'h0;
    end else if (_T_47) begin
      enableVector_5 <= 1'h0;
    end else begin
      enableVector_5 <= _T_142;
    end
    if (reset) begin
      _T_145 <= 7'h0;
    end else if (_T_47) begin
      _T_145 <= 7'h0;
    end else begin
      _T_145 <= _T_138;
    end
    if (reset) begin
      _T_146 <= 7'h0;
    end else if (_T_47) begin
      _T_146 <= 7'h0;
    end else begin
      _T_146 <= _T_145;
    end
    if (reset) begin
      _T_147 <= 7'h0;
    end else if (_T_47) begin
      _T_147 <= 7'h0;
    end else begin
      _T_147 <= _T_146;
    end
    if (reset) begin
      _T_148 <= 7'h0;
    end else if (_T_47) begin
      _T_148 <= 7'h0;
    end else begin
      _T_148 <= _T_147;
    end
    _T_171 <= _T_37 | _T_95;
    _T_283 <= _T_278 & _T_281;
    if (_T_283) begin
      _T_295_real <= _T_286_real;
    end else begin
      _T_295_real <= sdf_stages_0_io_out_real;
    end
    if (_T_283) begin
      _T_295_imag <= _T_289;
    end else begin
      _T_295_imag <= sdf_stages_0_io_out_imag;
    end
    _T_298_real <= _T_295_real;
    _T_298_imag <= _T_295_imag;
    outputWires_0_real <= _T_298_real;
    outputWires_0_imag <= _T_298_imag;
    if (_GEN_160) begin
      _T_481 <= _T_479;
    end
    if (5'h1e == _GEN_312) begin
      twiddles_1_real <= -16'sh1294;
    end else if (5'h1d == _GEN_312) begin
      twiddles_1_real <= -16'sh238e;
    end else if (5'h1c == _GEN_312) begin
      twiddles_1_real <= -16'sh3179;
    end else if (5'h1b == _GEN_312) begin
      twiddles_1_real <= -16'sh3b21;
    end else if (5'h1a == _GEN_312) begin
      twiddles_1_real <= -16'sh3fb1;
    end else if (5'h19 == _GEN_312) begin
      twiddles_1_real <= -16'sh3ec5;
    end else if (5'h18 == _GEN_312) begin
      twiddles_1_real <= -16'sh3b21;
    end else if (5'h17 == _GEN_312) begin
      twiddles_1_real <= -16'sh3871;
    end else if (5'h16 == _GEN_312) begin
      twiddles_1_real <= -16'sh3537;
    end else if (5'h15 == _GEN_312) begin
      twiddles_1_real <= -16'sh2d41;
    end else if (5'h14 == _GEN_312) begin
      twiddles_1_real <= -16'sh238e;
    end else if (5'h13 == _GEN_312) begin
      twiddles_1_real <= -16'sh1e2b;
    end else if (5'h12 == _GEN_312) begin
      twiddles_1_real <= -16'sh187e;
    end else if (5'h11 == _GEN_312) begin
      twiddles_1_real <= -16'shc7c;
    end else if (5'h10 == _GEN_312) begin
      twiddles_1_real <= 16'sh0;
    end else if (5'hf == _GEN_312) begin
      twiddles_1_real <= 16'sh646;
    end else if (5'he == _GEN_312) begin
      twiddles_1_real <= 16'shc7c;
    end else if (5'hd == _GEN_312) begin
      twiddles_1_real <= 16'sh1294;
    end else if (5'hc == _GEN_312) begin
      twiddles_1_real <= 16'sh187e;
    end else if (5'hb == _GEN_312) begin
      twiddles_1_real <= 16'sh1e2b;
    end else if (5'ha == _GEN_312) begin
      twiddles_1_real <= 16'sh238e;
    end else if (5'h9 == _GEN_312) begin
      twiddles_1_real <= 16'sh289a;
    end else if (5'h8 == _GEN_312) begin
      twiddles_1_real <= 16'sh2d41;
    end else if (5'h7 == _GEN_312) begin
      twiddles_1_real <= 16'sh3179;
    end else if (5'h6 == _GEN_312) begin
      twiddles_1_real <= 16'sh3537;
    end else if (5'h5 == _GEN_312) begin
      twiddles_1_real <= 16'sh3871;
    end else if (5'h4 == _GEN_312) begin
      twiddles_1_real <= 16'sh3b21;
    end else if (5'h3 == _GEN_312) begin
      twiddles_1_real <= 16'sh3d3f;
    end else if (5'h2 == _GEN_312) begin
      twiddles_1_real <= 16'sh3ec5;
    end else if (5'h1 == _GEN_312) begin
      twiddles_1_real <= 16'sh3fb1;
    end else begin
      twiddles_1_real <= 16'sh4000;
    end
    if (5'h1e == _GEN_312) begin
      twiddles_1_imag <= 16'sh3d3f;
    end else if (5'h1d == _GEN_312) begin
      twiddles_1_imag <= 16'sh3537;
    end else if (5'h1c == _GEN_312) begin
      twiddles_1_imag <= 16'sh289a;
    end else if (5'h1b == _GEN_312) begin
      twiddles_1_imag <= 16'sh187e;
    end else if (5'h1a == _GEN_312) begin
      twiddles_1_imag <= 16'sh646;
    end else if (5'h19 == _GEN_312) begin
      twiddles_1_imag <= -16'shc7c;
    end else if (5'h18 == _GEN_312) begin
      twiddles_1_imag <= -16'sh187e;
    end else if (5'h17 == _GEN_312) begin
      twiddles_1_imag <= -16'sh1e2b;
    end else if (5'h16 == _GEN_312) begin
      twiddles_1_imag <= -16'sh238e;
    end else if (5'h15 == _GEN_312) begin
      twiddles_1_imag <= -16'sh2d41;
    end else if (5'h14 == _GEN_312) begin
      twiddles_1_imag <= -16'sh3537;
    end else if (5'h13 == _GEN_312) begin
      twiddles_1_imag <= -16'sh3871;
    end else if (5'h12 == _GEN_312) begin
      twiddles_1_imag <= -16'sh3b21;
    end else if (5'h11 == _GEN_312) begin
      twiddles_1_imag <= -16'sh3ec5;
    end else if (5'h10 == _GEN_312) begin
      twiddles_1_imag <= -16'sh4000;
    end else if (5'hf == _GEN_312) begin
      twiddles_1_imag <= -16'sh3fb1;
    end else if (5'he == _GEN_312) begin
      twiddles_1_imag <= -16'sh3ec5;
    end else if (5'hd == _GEN_312) begin
      twiddles_1_imag <= -16'sh3d3f;
    end else if (5'hc == _GEN_312) begin
      twiddles_1_imag <= -16'sh3b21;
    end else if (5'hb == _GEN_312) begin
      twiddles_1_imag <= -16'sh3871;
    end else if (5'ha == _GEN_312) begin
      twiddles_1_imag <= -16'sh3537;
    end else if (5'h9 == _GEN_312) begin
      twiddles_1_imag <= -16'sh3179;
    end else if (5'h8 == _GEN_312) begin
      twiddles_1_imag <= -16'sh2d41;
    end else if (5'h7 == _GEN_312) begin
      twiddles_1_imag <= -16'sh289a;
    end else if (5'h6 == _GEN_312) begin
      twiddles_1_imag <= -16'sh238e;
    end else if (5'h5 == _GEN_312) begin
      twiddles_1_imag <= -16'sh1e2b;
    end else if (5'h4 == _GEN_312) begin
      twiddles_1_imag <= -16'sh187e;
    end else if (5'h3 == _GEN_312) begin
      twiddles_1_imag <= -16'sh1294;
    end else if (5'h2 == _GEN_312) begin
      twiddles_1_imag <= -16'shc7c;
    end else if (5'h1 == _GEN_312) begin
      twiddles_1_imag <= -16'sh646;
    end else begin
      twiddles_1_imag <= 16'sh0;
    end
    _T_490 <= sdf_stages_1_io_out_real;
    _T_491 <= twiddles_1_real;
    _T_492 <= twiddles_1_imag;
    _T_494 <= $signed(twiddles_1_real) + $signed(twiddles_1_imag);
    _T_496 <= $signed(sdf_stages_1_io_out_real) + $signed(sdf_stages_1_io_out_imag);
    _T_498 <= $signed(sdf_stages_1_io_out_imag) - $signed(sdf_stages_1_io_out_real);
    _T_500 <= $signed(_GEN_578) * $signed(_T_494);
    _T_506 <= $signed(_T_496) * $signed(_GEN_580);
    _T_512 <= $signed(_T_498) * $signed(_GEN_582);
    _T_518 <= $signed(_T_504) - $signed(_T_510);
    _T_520 <= $signed(_T_504) + $signed(_T_516);
    _T_546 <= _T_541 & _T_544;
    if (_T_546) begin
      _T_558_real <= _T_549_real;
    end else begin
      _T_558_real <= sdf_stages_2_io_out_real;
    end
    if (_T_546) begin
      _T_558_imag <= _T_552;
    end else begin
      _T_558_imag <= sdf_stages_2_io_out_imag;
    end
    _T_561_real <= _T_558_real;
    _T_561_imag <= _T_558_imag;
    outputWires_2_real <= _T_561_real;
    outputWires_2_imag <= _T_561_imag;
    if (_GEN_184) begin
      _T_624 <= _T_622;
    end
    if (3'h6 == _GEN_499) begin
      twiddles_3_real <= -16'sh3b21;
    end else if (3'h5 == _GEN_499) begin
      twiddles_3_real <= -16'sh2d41;
    end else if (3'h4 == _GEN_499) begin
      twiddles_3_real <= 16'sh0;
    end else if (3'h3 == _GEN_499) begin
      twiddles_3_real <= 16'sh187e;
    end else if (3'h2 == _GEN_499) begin
      twiddles_3_real <= 16'sh2d41;
    end else if (3'h1 == _GEN_499) begin
      twiddles_3_real <= 16'sh3b21;
    end else begin
      twiddles_3_real <= 16'sh4000;
    end
    if (3'h6 == _GEN_499) begin
      twiddles_3_imag <= 16'sh187e;
    end else if (3'h5 == _GEN_499) begin
      twiddles_3_imag <= -16'sh2d41;
    end else if (3'h4 == _GEN_499) begin
      twiddles_3_imag <= -16'sh4000;
    end else if (3'h3 == _GEN_499) begin
      twiddles_3_imag <= -16'sh3b21;
    end else if (3'h2 == _GEN_499) begin
      twiddles_3_imag <= -16'sh2d41;
    end else if (3'h1 == _GEN_499) begin
      twiddles_3_imag <= -16'sh187e;
    end else begin
      twiddles_3_imag <= 16'sh0;
    end
    _T_634 <= sdf_stages_3_io_out_real;
    _T_635 <= twiddles_3_real;
    _T_636 <= twiddles_3_imag;
    _T_638 <= $signed(twiddles_3_real) + $signed(twiddles_3_imag);
    _T_640 <= $signed(sdf_stages_3_io_out_real) + $signed(sdf_stages_3_io_out_imag);
    _T_642 <= $signed(sdf_stages_3_io_out_imag) - $signed(sdf_stages_3_io_out_real);
    _T_644 <= $signed(_GEN_586) * $signed(_T_638);
    _T_650 <= $signed(_T_640) * $signed(_GEN_588);
    _T_656 <= $signed(_T_642) * $signed(_GEN_590);
    _T_662 <= $signed(_T_648) - $signed(_T_654);
    _T_664 <= $signed(_T_648) + $signed(_T_660);
    _T_690 <= _T_685 & _T_688;
    if (_T_690) begin
      _T_702_real <= _T_693_real;
    end else begin
      _T_702_real <= sdf_stages_4_io_out_real;
    end
    if (_T_690) begin
      _T_702_imag <= _T_696;
    end else begin
      _T_702_imag <= sdf_stages_4_io_out_imag;
    end
    _T_705_real <= _T_702_real;
    _T_705_imag <= _T_702_imag;
    outputWires_4_real <= _T_705_real;
    outputWires_4_imag <= _T_705_imag;
    _T_717_real <= sdf_stages_5_io_out_real;
    _T_717_imag <= sdf_stages_5_io_out_imag;
    _T_720_real <= _T_717_real;
    _T_720_imag <= _T_717_imag;
    outputWires_5_real <= _T_720_real;
    outputWires_5_imag <= _T_720_imag;
    if (reset) begin
      _T_725 <= 1'h0;
    end else if (_T_47) begin
      _T_725 <= 1'h0;
    end else if (_T_170) begin
      _T_725 <= _T_173;
    end else begin
      _T_725 <= _T_174;
    end
    if (reset) begin
      _T_726 <= 1'h0;
    end else if (_T_47) begin
      _T_726 <= 1'h0;
    end else begin
      _T_726 <= _T_725;
    end
    if (reset) begin
      _T_727 <= 1'h0;
    end else if (_T_47) begin
      _T_727 <= 1'h0;
    end else begin
      _T_727 <= _T_726;
    end
    if (reset) begin
      outValid <= 1'h0;
    end else if (_T_47) begin
      outValid <= 1'h0;
    end else begin
      outValid <= _T_727;
    end
    if (reset) begin
      _T_729 <= 1'h0;
    end else begin
      _T_729 <= _T_728;
    end
    if (reset) begin
      _T_730 <= 1'h0;
    end else begin
      _T_730 <= _T_729;
    end
    if (reset) begin
      _T_731 <= 1'h0;
    end else begin
      _T_731 <= _T_730;
    end
    if (reset) begin
      _T_732 <= 1'h0;
    end else begin
      _T_732 <= _T_731;
    end
  end
endmodule
module SDFFFT_64_16(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [15:0] io_in_bits_real,
  input  [15:0] io_in_bits_imag,
  input         io_out_ready,
  output        io_out_valid,
  output [15:0] io_out_bits_real,
  output [15:0] io_out_bits_imag,
  output        io_lastOut,
  input         io_lastIn,
  input  [5:0]  io_fftSize,
  output        io_busy
);
  wire  SDFChainRadix22_clock; // @[SDFFFT.scala 418:119]
  wire  SDFChainRadix22_reset; // @[SDFFFT.scala 418:119]
  wire  SDFChainRadix22_io_in_ready; // @[SDFFFT.scala 418:119]
  wire  SDFChainRadix22_io_in_valid; // @[SDFFFT.scala 418:119]
  wire [15:0] SDFChainRadix22_io_in_bits_real; // @[SDFFFT.scala 418:119]
  wire [15:0] SDFChainRadix22_io_in_bits_imag; // @[SDFFFT.scala 418:119]
  wire  SDFChainRadix22_io_out_ready; // @[SDFFFT.scala 418:119]
  wire  SDFChainRadix22_io_out_valid; // @[SDFFFT.scala 418:119]
  wire [15:0] SDFChainRadix22_io_out_bits_real; // @[SDFFFT.scala 418:119]
  wire [15:0] SDFChainRadix22_io_out_bits_imag; // @[SDFFFT.scala 418:119]
  wire  SDFChainRadix22_io_lastOut; // @[SDFFFT.scala 418:119]
  wire  SDFChainRadix22_io_lastIn; // @[SDFFFT.scala 418:119]
  wire [5:0] SDFChainRadix22_io_fftSize; // @[SDFFFT.scala 418:119]
  wire  SDFChainRadix22_io_busy; // @[SDFFFT.scala 418:119]
  reg [5:0] cntWin; // @[SDFFFT.scala 265:23]
  reg [31:0] _RAND_0;
  wire [5:0] _T_5; // @[SDFFFT.scala 269:41]
  wire [64:0] _T_6; // @[SDFFFT.scala 269:23]
  wire  _T_7; // @[Decoupled.scala 40:37]
  wire [5:0] _T_9; // @[SDFFFT.scala 274:22]
  wire [5:0] numPoints; // @[SDFFFT.scala 266:23 SDFFFT.scala 269:15]
  wire [5:0] _T_11; // @[SDFFFT.scala 276:44]
  wire  _T_12; // @[SDFFFT.scala 276:29]
  wire  _T_13; // @[SDFFFT.scala 276:19]
  wire [31:0] _T_65; // @[FixedPointTypeClass.scala 42:59]
  wire [31:0] _T_66; // @[FixedPointTypeClass.scala 42:59]
  wire [29:0] _GEN_74; // @[SDFFFT.scala 500:56]
  wire [31:0] _GEN_70; // @[SDFFFT.scala 500:56]
  wire [29:0] _GEN_75; // @[SDFFFT.scala 500:56]
  wire [31:0] _GEN_71; // @[SDFFFT.scala 500:56]
  wire [17:0] _GEN_76; // @[SDFFFT.scala 508:18 SDFFFT.scala 513:28]
  wire [17:0] _GEN_78; // @[SDFFFT.scala 508:18 SDFFFT.scala 514:28]
  wire [17:0] _GEN_80; // @[SDFFFT.scala 503:31 SDFFFT.scala 511:21]
  wire [17:0] _GEN_82; // @[SDFFFT.scala 504:31 SDFFFT.scala 511:21]
  SDFChainRadix22 SDFChainRadix22 ( // @[SDFFFT.scala 418:119]
    .clock(SDFChainRadix22_clock),
    .reset(SDFChainRadix22_reset),
    .io_in_ready(SDFChainRadix22_io_in_ready),
    .io_in_valid(SDFChainRadix22_io_in_valid),
    .io_in_bits_real(SDFChainRadix22_io_in_bits_real),
    .io_in_bits_imag(SDFChainRadix22_io_in_bits_imag),
    .io_out_ready(SDFChainRadix22_io_out_ready),
    .io_out_valid(SDFChainRadix22_io_out_valid),
    .io_out_bits_real(SDFChainRadix22_io_out_bits_real),
    .io_out_bits_imag(SDFChainRadix22_io_out_bits_imag),
    .io_lastOut(SDFChainRadix22_io_lastOut),
    .io_lastIn(SDFChainRadix22_io_lastIn),
    .io_fftSize(SDFChainRadix22_io_fftSize),
    .io_busy(SDFChainRadix22_io_busy)
  );
  assign _T_5 = io_fftSize - 6'h1; // @[SDFFFT.scala 269:41]
  assign _T_6 = 65'h2 << _T_5; // @[SDFFFT.scala 269:23]
  assign _T_7 = io_in_ready & io_in_valid; // @[Decoupled.scala 40:37]
  assign _T_9 = cntWin + 6'h1; // @[SDFFFT.scala 274:22]
  assign numPoints = _T_6[5:0]; // @[SDFFFT.scala 266:23 SDFFFT.scala 269:15]
  assign _T_11 = numPoints - 6'h1; // @[SDFFFT.scala 276:44]
  assign _T_12 = cntWin == _T_11; // @[SDFFFT.scala 276:29]
  assign _T_13 = io_lastIn | _T_12; // @[SDFFFT.scala 276:19]
  assign _T_65 = $signed(io_in_bits_real) * 16'sh4000; // @[FixedPointTypeClass.scala 42:59]
  assign _T_66 = $signed(io_in_bits_imag) * 16'sh4000; // @[FixedPointTypeClass.scala 42:59]
  assign _GEN_74 = {$signed(SDFChainRadix22_io_out_bits_imag), 14'h0}; // @[SDFFFT.scala 500:56]
  assign _GEN_70 = {{2{_GEN_74[29]}},_GEN_74}; // @[SDFFFT.scala 500:56]
  assign _GEN_75 = {$signed(SDFChainRadix22_io_out_bits_real), 14'h0}; // @[SDFFFT.scala 500:56]
  assign _GEN_71 = {{2{_GEN_75[29]}},_GEN_75}; // @[SDFFFT.scala 500:56]
  assign io_in_ready = SDFChainRadix22_io_in_ready; // @[SDFFFT.scala 507:23 SDFFFT.scala 511:21]
  assign io_out_valid = SDFChainRadix22_io_out_valid; // @[SDFFFT.scala 508:18 SDFFFT.scala 516:24]
  assign _GEN_76 = _GEN_71[31:14]; // @[SDFFFT.scala 508:18 SDFFFT.scala 513:28]
  assign io_out_bits_real = _GEN_76[15:0]; // @[SDFFFT.scala 508:18 SDFFFT.scala 513:28]
  assign _GEN_78 = _GEN_70[31:14]; // @[SDFFFT.scala 508:18 SDFFFT.scala 514:28]
  assign io_out_bits_imag = _GEN_78[15:0]; // @[SDFFFT.scala 508:18 SDFFFT.scala 514:28]
  assign io_lastOut = SDFChainRadix22_io_lastOut; // @[SDFFFT.scala 520:20]
  assign io_busy = SDFChainRadix22_io_busy; // @[SDFFFT.scala 523:15]
  assign SDFChainRadix22_clock = clock;
  assign SDFChainRadix22_reset = reset;
  assign SDFChainRadix22_io_in_valid = io_in_valid; // @[SDFFFT.scala 506:27 SDFFFT.scala 511:21]
  assign _GEN_80 = _T_65[31:14]; // @[SDFFFT.scala 503:31 SDFFFT.scala 511:21]
  assign SDFChainRadix22_io_in_bits_real = _GEN_80[15:0]; // @[SDFFFT.scala 503:31 SDFFFT.scala 511:21]
  assign _GEN_82 = _T_66[31:14]; // @[SDFFFT.scala 504:31 SDFFFT.scala 511:21]
  assign SDFChainRadix22_io_in_bits_imag = _GEN_82[15:0]; // @[SDFFFT.scala 504:31 SDFFFT.scala 511:21]
  assign SDFChainRadix22_io_out_ready = io_out_ready; // @[SDFFFT.scala 508:18 SDFFFT.scala 517:28]
  assign SDFChainRadix22_io_lastIn = io_lastIn; // @[SDFFFT.scala 519:23]
  assign SDFChainRadix22_io_fftSize = io_fftSize; // @[SDFFFT.scala 526:28]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cntWin = _RAND_0[5:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      cntWin <= 6'h0;
    end else if (_T_13) begin
      cntWin <= 6'h0;
    end else if (_T_7) begin
      cntWin <= _T_9;
    end
  end
endmodule
module AXI4FFTBlock(
  input         clock,
  input         reset,
  output        auto_mem_in_aw_ready,
  input         auto_mem_in_aw_valid,
  input         auto_mem_in_aw_bits_id,
  input  [29:0] auto_mem_in_aw_bits_addr,
  output        auto_mem_in_w_ready,
  input         auto_mem_in_w_valid,
  input  [31:0] auto_mem_in_w_bits_data,
  input  [3:0]  auto_mem_in_w_bits_strb,
  input         auto_mem_in_b_ready,
  output        auto_mem_in_b_valid,
  output        auto_mem_in_b_bits_id,
  output        auto_mem_in_ar_ready,
  input         auto_mem_in_ar_valid,
  input         auto_mem_in_ar_bits_id,
  input  [29:0] auto_mem_in_ar_bits_addr,
  input  [2:0]  auto_mem_in_ar_bits_size,
  input         auto_mem_in_r_ready,
  output        auto_mem_in_r_valid,
  output        auto_mem_in_r_bits_id,
  output [31:0] auto_mem_in_r_bits_data,
  output        auto_stream_in_ready,
  input         auto_stream_in_valid,
  input  [31:0] auto_stream_in_bits_data,
  input         auto_stream_in_bits_last,
  input         auto_stream_out_ready,
  output        auto_stream_out_valid,
  output [31:0] auto_stream_out_bits_data,
  output        auto_stream_out_bits_last
);
  wire  fft_clock; // @[FFTBlock.scala 53:21]
  wire  fft_reset; // @[FFTBlock.scala 53:21]
  wire  fft_io_in_ready; // @[FFTBlock.scala 53:21]
  wire  fft_io_in_valid; // @[FFTBlock.scala 53:21]
  wire [15:0] fft_io_in_bits_real; // @[FFTBlock.scala 53:21]
  wire [15:0] fft_io_in_bits_imag; // @[FFTBlock.scala 53:21]
  wire  fft_io_out_ready; // @[FFTBlock.scala 53:21]
  wire  fft_io_out_valid; // @[FFTBlock.scala 53:21]
  wire [15:0] fft_io_out_bits_real; // @[FFTBlock.scala 53:21]
  wire [15:0] fft_io_out_bits_imag; // @[FFTBlock.scala 53:21]
  wire  fft_io_lastOut; // @[FFTBlock.scala 53:21]
  wire  fft_io_lastIn; // @[FFTBlock.scala 53:21]
  wire [5:0] fft_io_fftSize; // @[FFTBlock.scala 53:21]
  wire  fft_io_busy; // @[FFTBlock.scala 53:21]
  wire  Queue_clock; // @[Decoupled.scala 287:21]
  wire  Queue_reset; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_read; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_enq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_extra; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_read; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_deq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_extra; // @[Decoupled.scala 287:21]
  reg [2:0] fftSize; // @[FFTBlock.scala 59:34]
  reg [31:0] _RAND_0;
  reg  fftDir; // @[FFTBlock.scala 60:34]
  reg [31:0] _RAND_1;
  reg [5:0] keepMSBorLSBReg; // @[FFTBlock.scala 61:34]
  reg [31:0] _RAND_2;
  reg  busy; // @[FFTBlock.scala 64:34]
  reg [31:0] _RAND_3;
  wire  _T_2; // @[RegisterRouter.scala 40:39]
  wire  _T_3; // @[RegisterRouter.scala 40:26]
  wire  _T_4; // @[RegisterRouter.scala 42:29]
  wire  _T_47_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 290:17]
  wire [29:0] _T_11; // @[RegisterRouter.scala 48:19]
  wire [2:0] _T_226; // @[Cat.scala 29:58]
  wire [5:0] _T_51; // @[RegisterRouter.scala 59:16]
  wire  _T_61; // @[RegisterRouter.scala 59:16]
  wire  _T_5; // @[RegisterRouter.scala 42:26]
  wire [1:0] _T_14; // @[OneHot.scala 65:12]
  wire [1:0] _T_16; // @[Misc.scala 200:81]
  wire  _T_17; // @[Misc.scala 204:21]
  wire  _T_20; // @[Misc.scala 209:20]
  wire  _T_22; // @[Misc.scala 213:38]
  wire  _T_23; // @[Misc.scala 213:29]
  wire  _T_25; // @[Misc.scala 213:38]
  wire  _T_26; // @[Misc.scala 213:29]
  wire  _T_29; // @[Misc.scala 209:20]
  wire  _T_30; // @[Misc.scala 212:27]
  wire  _T_31; // @[Misc.scala 213:38]
  wire  _T_32; // @[Misc.scala 213:29]
  wire  _T_33; // @[Misc.scala 212:27]
  wire  _T_34; // @[Misc.scala 213:38]
  wire  _T_35; // @[Misc.scala 213:29]
  wire  _T_36; // @[Misc.scala 212:27]
  wire  _T_37; // @[Misc.scala 213:38]
  wire  _T_38; // @[Misc.scala 213:29]
  wire  _T_39; // @[Misc.scala 212:27]
  wire  _T_40; // @[Misc.scala 213:38]
  wire  _T_41; // @[Misc.scala 213:29]
  wire [3:0] _T_44; // @[Cat.scala 29:58]
  wire [3:0] _T_46; // @[RegisterRouter.scala 54:25]
  wire [7:0] _T_71; // @[Bitwise.scala 72:12]
  wire [7:0] _T_73; // @[Bitwise.scala 72:12]
  wire [7:0] _T_75; // @[Bitwise.scala 72:12]
  wire [7:0] _T_77; // @[Bitwise.scala 72:12]
  wire [31:0] _T_80; // @[Cat.scala 29:58]
  wire  _T_99; // @[RegisterRouter.scala 59:16]
  wire  _T_245; // @[RegisterRouter.scala 59:16]
  wire [7:0] _T_227; // @[OneHot.scala 58:35]
  wire  _T_292; // @[RegisterRouter.scala 59:16]
  wire  _T_294; // @[RegisterRouter.scala 59:16]
  wire  _T_295; // @[RegisterRouter.scala 59:16]
  wire  _T_106; // @[RegisterRouter.scala 59:16]
  wire  _T_299; // @[RegisterRouter.scala 59:16]
  wire  _T_300; // @[RegisterRouter.scala 59:16]
  wire  _T_129; // @[RegisterRouter.scala 59:16]
  wire  _GEN_1; // @[RegField.scala 134:88]
  wire  _T_145; // @[RegisterRouter.scala 59:16]
  wire  _T_304; // @[RegisterRouter.scala 59:16]
  wire  _T_305; // @[RegisterRouter.scala 59:16]
  wire  _T_152; // @[RegisterRouter.scala 59:16]
  wire  _GEN_36; // @[MuxLiteral.scala 48:10]
  wire  _GEN_37; // @[MuxLiteral.scala 48:10]
  wire  _GEN_38; // @[MuxLiteral.scala 48:10]
  wire  _GEN_39; // @[MuxLiteral.scala 48:10]
  wire  _GEN_51; // @[MuxLiteral.scala 48:10]
  wire  _GEN_40; // @[MuxLiteral.scala 48:10]
  wire  _GEN_52; // @[MuxLiteral.scala 48:10]
  wire  _GEN_41; // @[MuxLiteral.scala 48:10]
  wire  _GEN_53; // @[MuxLiteral.scala 48:10]
  wire  _GEN_42; // @[MuxLiteral.scala 48:10]
  wire [5:0] _T_437_0; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [5:0] _T_437_1; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [5:0] _GEN_44; // @[MuxLiteral.scala 48:10]
  wire [5:0] _GEN_45; // @[MuxLiteral.scala 48:10]
  wire [5:0] _T_437_3; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [5:0] _GEN_46; // @[MuxLiteral.scala 48:10]
  wire [5:0] _GEN_47; // @[MuxLiteral.scala 48:10]
  wire [5:0] _GEN_48; // @[MuxLiteral.scala 48:10]
  wire [5:0] _GEN_49; // @[MuxLiteral.scala 48:10]
  wire [5:0] _GEN_50; // @[MuxLiteral.scala 48:10]
  wire [5:0] _T_439; // @[RegisterRouter.scala 59:16]
  wire  _T_440_bits_read; // @[Decoupled.scala 308:19 Decoupled.scala 309:14]
  wire  _T_440_valid; // @[Decoupled.scala 308:19 Decoupled.scala 310:15]
  wire  _T_443; // @[RegisterRouter.scala 65:29]
  SDFFFT_64_16 fft ( // @[FFTBlock.scala 53:21]
    .clock(fft_clock),
    .reset(fft_reset),
    .io_in_ready(fft_io_in_ready),
    .io_in_valid(fft_io_in_valid),
    .io_in_bits_real(fft_io_in_bits_real),
    .io_in_bits_imag(fft_io_in_bits_imag),
    .io_out_ready(fft_io_out_ready),
    .io_out_valid(fft_io_out_valid),
    .io_out_bits_real(fft_io_out_bits_real),
    .io_out_bits_imag(fft_io_out_bits_imag),
    .io_lastOut(fft_io_lastOut),
    .io_lastIn(fft_io_lastIn),
    .io_fftSize(fft_io_fftSize),
    .io_busy(fft_io_busy)
  );
  Queue Queue ( // @[Decoupled.scala 287:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_read(Queue_io_enq_bits_read),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_extra(Queue_io_enq_bits_extra),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_read(Queue_io_deq_bits_read),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_extra(Queue_io_deq_bits_extra)
  );
  assign _T_2 = auto_mem_in_aw_valid & auto_mem_in_w_valid; // @[RegisterRouter.scala 40:39]
  assign _T_3 = auto_mem_in_ar_valid | _T_2; // @[RegisterRouter.scala 40:26]
  assign _T_4 = ~auto_mem_in_ar_valid; // @[RegisterRouter.scala 42:29]
  assign _T_47_ready = Queue_io_enq_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 290:17]
  assign _T_11 = auto_mem_in_ar_valid ? auto_mem_in_ar_bits_addr : auto_mem_in_aw_bits_addr; // @[RegisterRouter.scala 48:19]
  assign _T_226 = {_T_11[4],_T_11[3],_T_11[2]}; // @[Cat.scala 29:58]
  assign _T_51 = _T_11[7:2] & 6'h38; // @[RegisterRouter.scala 59:16]
  assign _T_61 = _T_51 == 6'h0; // @[RegisterRouter.scala 59:16]
  assign _T_5 = _T_47_ready & _T_4; // @[RegisterRouter.scala 42:26]
  assign _T_14 = 2'h1 << auto_mem_in_ar_bits_size[0]; // @[OneHot.scala 65:12]
  assign _T_16 = _T_14 | 2'h1; // @[Misc.scala 200:81]
  assign _T_17 = auto_mem_in_ar_bits_size >= 3'h2; // @[Misc.scala 204:21]
  assign _T_20 = ~auto_mem_in_ar_bits_addr[1]; // @[Misc.scala 209:20]
  assign _T_22 = _T_16[1] & _T_20; // @[Misc.scala 213:38]
  assign _T_23 = _T_17 | _T_22; // @[Misc.scala 213:29]
  assign _T_25 = _T_16[1] & auto_mem_in_ar_bits_addr[1]; // @[Misc.scala 213:38]
  assign _T_26 = _T_17 | _T_25; // @[Misc.scala 213:29]
  assign _T_29 = ~auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 209:20]
  assign _T_30 = _T_20 & _T_29; // @[Misc.scala 212:27]
  assign _T_31 = _T_16[0] & _T_30; // @[Misc.scala 213:38]
  assign _T_32 = _T_23 | _T_31; // @[Misc.scala 213:29]
  assign _T_33 = _T_20 & auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  assign _T_34 = _T_16[0] & _T_33; // @[Misc.scala 213:38]
  assign _T_35 = _T_23 | _T_34; // @[Misc.scala 213:29]
  assign _T_36 = auto_mem_in_ar_bits_addr[1] & _T_29; // @[Misc.scala 212:27]
  assign _T_37 = _T_16[0] & _T_36; // @[Misc.scala 213:38]
  assign _T_38 = _T_26 | _T_37; // @[Misc.scala 213:29]
  assign _T_39 = auto_mem_in_ar_bits_addr[1] & auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  assign _T_40 = _T_16[0] & _T_39; // @[Misc.scala 213:38]
  assign _T_41 = _T_26 | _T_40; // @[Misc.scala 213:29]
  assign _T_44 = {_T_41,_T_38,_T_35,_T_32}; // @[Cat.scala 29:58]
  assign _T_46 = auto_mem_in_ar_valid ? _T_44 : auto_mem_in_w_bits_strb; // @[RegisterRouter.scala 54:25]
  assign _T_71 = _T_46[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_73 = _T_46[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_75 = _T_46[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_77 = _T_46[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_80 = {_T_77,_T_75,_T_73,_T_71}; // @[Cat.scala 29:58]
  assign _T_99 = _T_80[2:0] == 3'h7; // @[RegisterRouter.scala 59:16]
  assign _T_245 = _T_3 & _T_47_ready; // @[RegisterRouter.scala 59:16]
  assign _T_227 = 8'h1 << _T_226; // @[OneHot.scala 58:35]
  assign _T_292 = _T_245 & _T_4; // @[RegisterRouter.scala 59:16]
  assign _T_294 = _T_292 & _T_227[0]; // @[RegisterRouter.scala 59:16]
  assign _T_295 = _T_294 & _T_61; // @[RegisterRouter.scala 59:16]
  assign _T_106 = _T_295 & _T_99; // @[RegisterRouter.scala 59:16]
  assign _T_299 = _T_292 & _T_227[1]; // @[RegisterRouter.scala 59:16]
  assign _T_300 = _T_299 & _T_61; // @[RegisterRouter.scala 59:16]
  assign _T_129 = _T_300 & _T_80[0]; // @[RegisterRouter.scala 59:16]
  assign _GEN_1 = _T_129 ? auto_mem_in_w_bits_data[0] : fftDir; // @[RegField.scala 134:88]
  assign _T_145 = _T_80[5:0] == 6'h3f; // @[RegisterRouter.scala 59:16]
  assign _T_304 = _T_292 & _T_227[2]; // @[RegisterRouter.scala 59:16]
  assign _T_305 = _T_304 & _T_61; // @[RegisterRouter.scala 59:16]
  assign _T_152 = _T_305 & _T_145; // @[RegisterRouter.scala 59:16]
  assign _GEN_36 = 3'h1 == _T_226 ? _T_61 : _T_61; // @[MuxLiteral.scala 48:10]
  assign _GEN_37 = 3'h2 == _T_226 ? _T_61 : _GEN_36; // @[MuxLiteral.scala 48:10]
  assign _GEN_38 = 3'h3 == _T_226 ? _T_61 : _GEN_37; // @[MuxLiteral.scala 48:10]
  assign _GEN_39 = 3'h4 == _T_226 ? _T_61 : _GEN_38; // @[MuxLiteral.scala 48:10]
  assign _GEN_51 = 3'h5 == _T_226; // @[MuxLiteral.scala 48:10]
  assign _GEN_40 = _GEN_51 | _GEN_39; // @[MuxLiteral.scala 48:10]
  assign _GEN_52 = 3'h6 == _T_226; // @[MuxLiteral.scala 48:10]
  assign _GEN_41 = _GEN_52 | _GEN_40; // @[MuxLiteral.scala 48:10]
  assign _GEN_53 = 3'h7 == _T_226; // @[MuxLiteral.scala 48:10]
  assign _GEN_42 = _GEN_53 | _GEN_41; // @[MuxLiteral.scala 48:10]
  assign _T_437_0 = {{3'd0}, fftSize}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  assign _T_437_1 = {{5'd0}, fftDir}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  assign _GEN_44 = 3'h1 == _T_226 ? _T_437_1 : _T_437_0; // @[MuxLiteral.scala 48:10]
  assign _GEN_45 = 3'h2 == _T_226 ? keepMSBorLSBReg : _GEN_44; // @[MuxLiteral.scala 48:10]
  assign _T_437_3 = {{5'd0}, busy}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  assign _GEN_46 = 3'h3 == _T_226 ? _T_437_3 : _GEN_45; // @[MuxLiteral.scala 48:10]
  assign _GEN_47 = 3'h4 == _T_226 ? 6'h0 : _GEN_46; // @[MuxLiteral.scala 48:10]
  assign _GEN_48 = 3'h5 == _T_226 ? 6'h0 : _GEN_47; // @[MuxLiteral.scala 48:10]
  assign _GEN_49 = 3'h6 == _T_226 ? 6'h0 : _GEN_48; // @[MuxLiteral.scala 48:10]
  assign _GEN_50 = 3'h7 == _T_226 ? 6'h0 : _GEN_49; // @[MuxLiteral.scala 48:10]
  assign _T_439 = _GEN_42 ? _GEN_50 : 6'h0; // @[RegisterRouter.scala 59:16]
  assign _T_440_bits_read = Queue_io_deq_bits_read; // @[Decoupled.scala 308:19 Decoupled.scala 309:14]
  assign _T_440_valid = Queue_io_deq_valid; // @[Decoupled.scala 308:19 Decoupled.scala 310:15]
  assign _T_443 = ~_T_440_bits_read; // @[RegisterRouter.scala 65:29]
  assign auto_mem_in_aw_ready = _T_5 & auto_mem_in_w_valid; // @[LazyModule.scala 173:31]
  assign auto_mem_in_w_ready = _T_5 & auto_mem_in_aw_valid; // @[LazyModule.scala 173:31]
  assign auto_mem_in_b_valid = _T_440_valid & _T_443; // @[LazyModule.scala 173:31]
  assign auto_mem_in_b_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_mem_in_ar_ready = Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_valid = _T_440_valid & _T_440_bits_read; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 173:31]
  assign auto_stream_in_ready = fft_io_in_ready; // @[LazyModule.scala 173:31]
  assign auto_stream_out_valid = fft_io_out_valid; // @[LazyModule.scala 173:49]
  assign auto_stream_out_bits_data = {fft_io_out_bits_real,fft_io_out_bits_imag}; // @[LazyModule.scala 173:49]
  assign auto_stream_out_bits_last = fft_io_lastOut; // @[LazyModule.scala 173:49]
  assign fft_clock = clock;
  assign fft_reset = reset;
  assign fft_io_in_valid = auto_stream_in_valid; // @[FFTBlock.scala 103:24]
  assign fft_io_in_bits_real = auto_stream_in_bits_data[31:16]; // @[FFTBlock.scala 104:24]
  assign fft_io_in_bits_imag = auto_stream_in_bits_data[15:0]; // @[FFTBlock.scala 104:24]
  assign fft_io_out_ready = auto_stream_out_ready; // @[FFTBlock.scala 111:22]
  assign fft_io_lastIn = auto_stream_in_bits_last; // @[FFTBlock.scala 106:24]
  assign fft_io_fftSize = {{3'd0}, fftSize}; // @[FFTBlock.scala 71:26]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_mem_in_ar_valid | _T_2; // @[Decoupled.scala 288:22]
  assign Queue_io_enq_bits_read = auto_mem_in_ar_valid; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_data = {{26'd0}, _T_439}; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_extra = auto_mem_in_ar_valid ? auto_mem_in_ar_bits_id : auto_mem_in_aw_bits_id; // @[Decoupled.scala 289:21]
  assign Queue_io_deq_ready = _T_440_bits_read ? auto_mem_in_r_ready : auto_mem_in_b_ready; // @[Decoupled.scala 311:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  fftSize = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  fftDir = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  keepMSBorLSBReg = _RAND_2[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  busy = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      fftSize <= 3'h6;
    end else if (_T_106) begin
      fftSize <= auto_mem_in_w_bits_data[2:0];
    end
    fftDir <= reset | _GEN_1;
    if (reset) begin
      keepMSBorLSBReg <= 6'h0;
    end else if (_T_152) begin
      keepMSBorLSBReg <= auto_mem_in_w_bits_data[5:0];
    end
    if (reset) begin
      busy <= 1'h0;
    end else begin
      busy <= fft_io_busy;
    end
  end
endmodule
module AXI4Splitter_3(
  input         clock,
  input         reset,
  output        auto_mem_in_aw_ready,
  input         auto_mem_in_aw_valid,
  input         auto_mem_in_aw_bits_id,
  input  [29:0] auto_mem_in_aw_bits_addr,
  output        auto_mem_in_w_ready,
  input         auto_mem_in_w_valid,
  input  [31:0] auto_mem_in_w_bits_data,
  input  [3:0]  auto_mem_in_w_bits_strb,
  input         auto_mem_in_b_ready,
  output        auto_mem_in_b_valid,
  output        auto_mem_in_b_bits_id,
  output        auto_mem_in_ar_ready,
  input         auto_mem_in_ar_valid,
  input         auto_mem_in_ar_bits_id,
  input  [29:0] auto_mem_in_ar_bits_addr,
  input  [2:0]  auto_mem_in_ar_bits_size,
  input         auto_mem_in_r_ready,
  output        auto_mem_in_r_valid,
  output        auto_mem_in_r_bits_id,
  output [31:0] auto_mem_in_r_bits_data,
  output        auto_stream_in_ready,
  input         auto_stream_in_valid,
  input  [31:0] auto_stream_in_bits_data,
  input         auto_stream_in_bits_last,
  input         auto_stream_out_1_ready,
  output        auto_stream_out_1_valid,
  output [31:0] auto_stream_out_1_bits_data,
  output        auto_stream_out_1_bits_last,
  input         auto_stream_out_0_ready,
  output        auto_stream_out_0_valid,
  output [31:0] auto_stream_out_0_bits_data,
  output        auto_stream_out_0_bits_last
);
  wire  Queue_clock; // @[Decoupled.scala 287:21]
  wire  Queue_reset; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_read; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_enq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_extra; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_read; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_deq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_extra; // @[Decoupled.scala 287:21]
  reg [31:0] ctrlReg; // @[Splitter.scala 27:26]
  reg [31:0] _RAND_0;
  reg [31:0] maskReg; // @[Splitter.scala 28:26]
  reg [31:0] _RAND_1;
  wire  _T_4; // @[RegisterRouter.scala 40:39]
  wire  _T_5; // @[RegisterRouter.scala 40:26]
  wire  _T_6; // @[RegisterRouter.scala 42:29]
  wire  _T_49_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 290:17]
  wire [29:0] _T_13; // @[RegisterRouter.scala 48:19]
  wire [1:0] _T_53; // @[RegisterRouter.scala 59:16]
  wire  _T_55; // @[RegisterRouter.scala 59:16]
  wire  _T_7; // @[RegisterRouter.scala 42:26]
  wire [1:0] _T_16; // @[OneHot.scala 65:12]
  wire [1:0] _T_18; // @[Misc.scala 200:81]
  wire  _T_19; // @[Misc.scala 204:21]
  wire  _T_22; // @[Misc.scala 209:20]
  wire  _T_24; // @[Misc.scala 213:38]
  wire  _T_25; // @[Misc.scala 213:29]
  wire  _T_27; // @[Misc.scala 213:38]
  wire  _T_28; // @[Misc.scala 213:29]
  wire  _T_31; // @[Misc.scala 209:20]
  wire  _T_32; // @[Misc.scala 212:27]
  wire  _T_33; // @[Misc.scala 213:38]
  wire  _T_34; // @[Misc.scala 213:29]
  wire  _T_35; // @[Misc.scala 212:27]
  wire  _T_36; // @[Misc.scala 213:38]
  wire  _T_37; // @[Misc.scala 213:29]
  wire  _T_38; // @[Misc.scala 212:27]
  wire  _T_39; // @[Misc.scala 213:38]
  wire  _T_40; // @[Misc.scala 213:29]
  wire  _T_41; // @[Misc.scala 212:27]
  wire  _T_42; // @[Misc.scala 213:38]
  wire  _T_43; // @[Misc.scala 213:29]
  wire [3:0] _T_46; // @[Cat.scala 29:58]
  wire [3:0] _T_48; // @[RegisterRouter.scala 54:25]
  wire [7:0] _T_67; // @[Bitwise.scala 72:12]
  wire [7:0] _T_69; // @[Bitwise.scala 72:12]
  wire [7:0] _T_71; // @[Bitwise.scala 72:12]
  wire [7:0] _T_73; // @[Bitwise.scala 72:12]
  wire [31:0] _T_76; // @[Cat.scala 29:58]
  wire  _T_95; // @[RegisterRouter.scala 59:16]
  wire  _T_148; // @[RegisterRouter.scala 59:16]
  wire [1:0] _T_142; // @[OneHot.scala 58:35]
  wire  _T_165; // @[RegisterRouter.scala 59:16]
  wire  _T_172; // @[RegisterRouter.scala 59:16]
  wire  _T_173; // @[RegisterRouter.scala 59:16]
  wire  _T_102; // @[RegisterRouter.scala 59:16]
  wire  _T_167; // @[RegisterRouter.scala 59:16]
  wire  _T_168; // @[RegisterRouter.scala 59:16]
  wire  _T_125; // @[RegisterRouter.scala 59:16]
  wire  _GEN_11; // @[MuxLiteral.scala 48:10]
  wire [31:0] _GEN_13; // @[MuxLiteral.scala 48:10]
  wire  _T_223_bits_read; // @[Decoupled.scala 308:19 Decoupled.scala 309:14]
  wire  _T_223_valid; // @[Decoupled.scala 308:19 Decoupled.scala 310:15]
  wire  _T_226; // @[RegisterRouter.scala 65:29]
  wire  readyOR; // @[Splitter.scala 45:34]
  wire  readyAND; // @[Splitter.scala 46:34]
  wire  _T_229; // @[Splitter.scala 49:19]
  wire  _T_230; // @[Splitter.scala 52:24]
  wire  _GEN_14; // @[Splitter.scala 52:33]
  wire  _T_233; // @[Splitter.scala 62:34]
  wire  _T_237; // @[Splitter.scala 62:34]
  Queue Queue ( // @[Decoupled.scala 287:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_read(Queue_io_enq_bits_read),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_extra(Queue_io_enq_bits_extra),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_read(Queue_io_deq_bits_read),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_extra(Queue_io_deq_bits_extra)
  );
  assign _T_4 = auto_mem_in_aw_valid & auto_mem_in_w_valid; // @[RegisterRouter.scala 40:39]
  assign _T_5 = auto_mem_in_ar_valid | _T_4; // @[RegisterRouter.scala 40:26]
  assign _T_6 = ~auto_mem_in_ar_valid; // @[RegisterRouter.scala 42:29]
  assign _T_49_ready = Queue_io_enq_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 290:17]
  assign _T_13 = auto_mem_in_ar_valid ? auto_mem_in_ar_bits_addr : auto_mem_in_aw_bits_addr; // @[RegisterRouter.scala 48:19]
  assign _T_53 = _T_13[3:2] & 2'h2; // @[RegisterRouter.scala 59:16]
  assign _T_55 = _T_53 == 2'h0; // @[RegisterRouter.scala 59:16]
  assign _T_7 = _T_49_ready & _T_6; // @[RegisterRouter.scala 42:26]
  assign _T_16 = 2'h1 << auto_mem_in_ar_bits_size[0]; // @[OneHot.scala 65:12]
  assign _T_18 = _T_16 | 2'h1; // @[Misc.scala 200:81]
  assign _T_19 = auto_mem_in_ar_bits_size >= 3'h2; // @[Misc.scala 204:21]
  assign _T_22 = ~auto_mem_in_ar_bits_addr[1]; // @[Misc.scala 209:20]
  assign _T_24 = _T_18[1] & _T_22; // @[Misc.scala 213:38]
  assign _T_25 = _T_19 | _T_24; // @[Misc.scala 213:29]
  assign _T_27 = _T_18[1] & auto_mem_in_ar_bits_addr[1]; // @[Misc.scala 213:38]
  assign _T_28 = _T_19 | _T_27; // @[Misc.scala 213:29]
  assign _T_31 = ~auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 209:20]
  assign _T_32 = _T_22 & _T_31; // @[Misc.scala 212:27]
  assign _T_33 = _T_18[0] & _T_32; // @[Misc.scala 213:38]
  assign _T_34 = _T_25 | _T_33; // @[Misc.scala 213:29]
  assign _T_35 = _T_22 & auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  assign _T_36 = _T_18[0] & _T_35; // @[Misc.scala 213:38]
  assign _T_37 = _T_25 | _T_36; // @[Misc.scala 213:29]
  assign _T_38 = auto_mem_in_ar_bits_addr[1] & _T_31; // @[Misc.scala 212:27]
  assign _T_39 = _T_18[0] & _T_38; // @[Misc.scala 213:38]
  assign _T_40 = _T_28 | _T_39; // @[Misc.scala 213:29]
  assign _T_41 = auto_mem_in_ar_bits_addr[1] & auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  assign _T_42 = _T_18[0] & _T_41; // @[Misc.scala 213:38]
  assign _T_43 = _T_28 | _T_42; // @[Misc.scala 213:29]
  assign _T_46 = {_T_43,_T_40,_T_37,_T_34}; // @[Cat.scala 29:58]
  assign _T_48 = auto_mem_in_ar_valid ? _T_46 : auto_mem_in_w_bits_strb; // @[RegisterRouter.scala 54:25]
  assign _T_67 = _T_48[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_69 = _T_48[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_71 = _T_48[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_73 = _T_48[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_76 = {_T_73,_T_71,_T_69,_T_67}; // @[Cat.scala 29:58]
  assign _T_95 = _T_76 == 32'hffffffff; // @[RegisterRouter.scala 59:16]
  assign _T_148 = _T_5 & _T_49_ready; // @[RegisterRouter.scala 59:16]
  assign _T_142 = 2'h1 << _T_13[2]; // @[OneHot.scala 58:35]
  assign _T_165 = _T_148 & _T_6; // @[RegisterRouter.scala 59:16]
  assign _T_172 = _T_165 & _T_142[1]; // @[RegisterRouter.scala 59:16]
  assign _T_173 = _T_172 & _T_55; // @[RegisterRouter.scala 59:16]
  assign _T_102 = _T_173 & _T_95; // @[RegisterRouter.scala 59:16]
  assign _T_167 = _T_165 & _T_142[0]; // @[RegisterRouter.scala 59:16]
  assign _T_168 = _T_167 & _T_55; // @[RegisterRouter.scala 59:16]
  assign _T_125 = _T_168 & _T_95; // @[RegisterRouter.scala 59:16]
  assign _GEN_11 = _T_13[2] ? _T_55 : _T_55; // @[MuxLiteral.scala 48:10]
  assign _GEN_13 = _T_13[2] ? maskReg : ctrlReg; // @[MuxLiteral.scala 48:10]
  assign _T_223_bits_read = Queue_io_deq_bits_read; // @[Decoupled.scala 308:19 Decoupled.scala 309:14]
  assign _T_223_valid = Queue_io_deq_valid; // @[Decoupled.scala 308:19 Decoupled.scala 310:15]
  assign _T_226 = ~_T_223_bits_read; // @[RegisterRouter.scala 65:29]
  assign readyOR = auto_stream_out_0_ready | auto_stream_out_1_ready; // @[Splitter.scala 45:34]
  assign readyAND = auto_stream_out_0_ready & auto_stream_out_1_ready; // @[Splitter.scala 46:34]
  assign _T_229 = ctrlReg == 32'h0; // @[Splitter.scala 49:19]
  assign _T_230 = ctrlReg == 32'h1; // @[Splitter.scala 52:24]
  assign _GEN_14 = _T_230 & readyOR; // @[Splitter.scala 52:33]
  assign _T_233 = ~maskReg[0]; // @[Splitter.scala 62:34]
  assign _T_237 = ~maskReg[1]; // @[Splitter.scala 62:34]
  assign auto_mem_in_aw_ready = _T_7 & auto_mem_in_w_valid; // @[LazyModule.scala 173:31]
  assign auto_mem_in_w_ready = _T_7 & auto_mem_in_aw_valid; // @[LazyModule.scala 173:31]
  assign auto_mem_in_b_valid = _T_223_valid & _T_226; // @[LazyModule.scala 173:31]
  assign auto_mem_in_b_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_mem_in_ar_ready = Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_valid = _T_223_valid & _T_223_bits_read; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 173:31]
  assign auto_stream_in_ready = _T_229 ? readyAND : _GEN_14; // @[LazyModule.scala 173:31]
  assign auto_stream_out_1_valid = auto_stream_in_valid & _T_237; // @[LazyModule.scala 173:49]
  assign auto_stream_out_1_bits_data = auto_stream_in_bits_data; // @[LazyModule.scala 173:49]
  assign auto_stream_out_1_bits_last = auto_stream_in_bits_last; // @[LazyModule.scala 173:49]
  assign auto_stream_out_0_valid = auto_stream_in_valid & _T_233; // @[LazyModule.scala 173:49]
  assign auto_stream_out_0_bits_data = auto_stream_in_bits_data; // @[LazyModule.scala 173:49]
  assign auto_stream_out_0_bits_last = auto_stream_in_bits_last; // @[LazyModule.scala 173:49]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_mem_in_ar_valid | _T_4; // @[Decoupled.scala 288:22]
  assign Queue_io_enq_bits_read = auto_mem_in_ar_valid; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_data = _GEN_11 ? _GEN_13 : 32'h0; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_extra = auto_mem_in_ar_valid ? auto_mem_in_ar_bits_id : auto_mem_in_aw_bits_id; // @[Decoupled.scala 289:21]
  assign Queue_io_deq_ready = _T_223_bits_read ? auto_mem_in_r_ready : auto_mem_in_b_ready; // @[Decoupled.scala 311:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ctrlReg = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  maskReg = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      ctrlReg <= 32'h0;
    end else if (_T_125) begin
      ctrlReg <= auto_mem_in_w_bits_data;
    end
    if (reset) begin
      maskReg <= 32'h0;
    end else if (_T_102) begin
      maskReg <= auto_mem_in_w_bits_data;
    end
  end
endmodule
module AXI4StreamMux_4(
  input         clock,
  input         reset,
  output        auto_register_in_aw_ready,
  input         auto_register_in_aw_valid,
  input         auto_register_in_aw_bits_id,
  input  [29:0] auto_register_in_aw_bits_addr,
  output        auto_register_in_w_ready,
  input         auto_register_in_w_valid,
  input  [31:0] auto_register_in_w_bits_data,
  input  [3:0]  auto_register_in_w_bits_strb,
  input         auto_register_in_b_ready,
  output        auto_register_in_b_valid,
  output        auto_register_in_b_bits_id,
  output        auto_register_in_ar_ready,
  input         auto_register_in_ar_valid,
  input         auto_register_in_ar_bits_id,
  input  [29:0] auto_register_in_ar_bits_addr,
  input  [2:0]  auto_register_in_ar_bits_size,
  input         auto_register_in_r_ready,
  output        auto_register_in_r_valid,
  output        auto_register_in_r_bits_id,
  output [31:0] auto_register_in_r_bits_data,
  output        auto_stream_in_2_ready,
  input         auto_stream_in_2_valid,
  input  [31:0] auto_stream_in_2_bits_data,
  input         auto_stream_in_2_bits_last,
  output        auto_stream_in_1_ready,
  input         auto_stream_in_1_valid,
  input  [31:0] auto_stream_in_1_bits_data,
  input         auto_stream_in_1_bits_last,
  output        auto_stream_in_0_ready,
  input         auto_stream_in_0_valid,
  input  [31:0] auto_stream_in_0_bits_data,
  input         auto_stream_in_0_bits_last,
  input         auto_stream_out_0_ready,
  output        auto_stream_out_0_valid,
  output [31:0] auto_stream_out_0_bits_data,
  output        auto_stream_out_0_bits_last
);
  wire  Queue_clock; // @[Decoupled.scala 287:21]
  wire  Queue_reset; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_read; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_enq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_extra; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_read; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_deq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_extra; // @[Decoupled.scala 287:21]
  reg [2:0] sels_0; // @[Mux.scala 32:23]
  reg [31:0] _RAND_0;
  reg [2:0] sels_1; // @[Mux.scala 32:23]
  reg [31:0] _RAND_1;
  wire  _T_3; // @[Mux.scala 45:28]
  wire  _GEN_7; // @[Mux.scala 45:41]
  wire  _GEN_8; // @[Mux.scala 45:41]
  wire  _T_4; // @[Mux.scala 45:28]
  wire  _GEN_12; // @[Mux.scala 45:41]
  wire [31:0] _GEN_15; // @[Mux.scala 45:41]
  wire  _GEN_16; // @[Mux.scala 45:41]
  wire  _GEN_17; // @[Mux.scala 45:41]
  wire  _T_5; // @[Mux.scala 45:28]
  wire  _GEN_21; // @[Mux.scala 45:41]
  wire [31:0] _GEN_24; // @[Mux.scala 45:41]
  wire  _GEN_25; // @[Mux.scala 45:41]
  wire  _GEN_26; // @[Mux.scala 45:41]
  wire  _T_6; // @[Mux.scala 45:28]
  wire  _GEN_30; // @[Mux.scala 45:41]
  wire [31:0] _GEN_33; // @[Mux.scala 45:41]
  wire  _GEN_34; // @[Mux.scala 45:41]
  wire  _T_7; // @[Mux.scala 45:28]
  wire  _T_8; // @[Mux.scala 40:46]
  wire [2:0] _T_10; // @[Mux.scala 41:29]
  wire  _T_11; // @[Mux.scala 45:28]
  wire  _T_12; // @[Mux.scala 45:28]
  wire  _T_13; // @[Mux.scala 45:28]
  wire  _T_17; // @[RegisterRouter.scala 40:39]
  wire  _T_18; // @[RegisterRouter.scala 40:26]
  wire  _T_19; // @[RegisterRouter.scala 42:29]
  wire  _T_62_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 290:17]
  wire [29:0] _T_26; // @[RegisterRouter.scala 48:19]
  wire [1:0] _T_66; // @[RegisterRouter.scala 59:16]
  wire  _T_68; // @[RegisterRouter.scala 59:16]
  wire  _T_20; // @[RegisterRouter.scala 42:26]
  wire [1:0] _T_29; // @[OneHot.scala 65:12]
  wire [1:0] _T_31; // @[Misc.scala 200:81]
  wire  _T_32; // @[Misc.scala 204:21]
  wire  _T_35; // @[Misc.scala 209:20]
  wire  _T_37; // @[Misc.scala 213:38]
  wire  _T_38; // @[Misc.scala 213:29]
  wire  _T_40; // @[Misc.scala 213:38]
  wire  _T_41; // @[Misc.scala 213:29]
  wire  _T_44; // @[Misc.scala 209:20]
  wire  _T_45; // @[Misc.scala 212:27]
  wire  _T_46; // @[Misc.scala 213:38]
  wire  _T_47; // @[Misc.scala 213:29]
  wire  _T_48; // @[Misc.scala 212:27]
  wire  _T_49; // @[Misc.scala 213:38]
  wire  _T_50; // @[Misc.scala 213:29]
  wire  _T_51; // @[Misc.scala 212:27]
  wire  _T_52; // @[Misc.scala 213:38]
  wire  _T_53; // @[Misc.scala 213:29]
  wire  _T_54; // @[Misc.scala 212:27]
  wire  _T_55; // @[Misc.scala 213:38]
  wire  _T_56; // @[Misc.scala 213:29]
  wire [3:0] _T_59; // @[Cat.scala 29:58]
  wire [3:0] _T_61; // @[RegisterRouter.scala 54:25]
  wire [7:0] _T_80; // @[Bitwise.scala 72:12]
  wire [7:0] _T_82; // @[Bitwise.scala 72:12]
  wire [7:0] _T_84; // @[Bitwise.scala 72:12]
  wire [7:0] _T_86; // @[Bitwise.scala 72:12]
  wire [31:0] _T_89; // @[Cat.scala 29:58]
  wire  _T_108; // @[RegisterRouter.scala 59:16]
  wire  _T_161; // @[RegisterRouter.scala 59:16]
  wire [1:0] _T_155; // @[OneHot.scala 58:35]
  wire  _T_178; // @[RegisterRouter.scala 59:16]
  wire  _T_185; // @[RegisterRouter.scala 59:16]
  wire  _T_186; // @[RegisterRouter.scala 59:16]
  wire  _T_115; // @[RegisterRouter.scala 59:16]
  wire  _T_180; // @[RegisterRouter.scala 59:16]
  wire  _T_181; // @[RegisterRouter.scala 59:16]
  wire  _T_138; // @[RegisterRouter.scala 59:16]
  wire  _GEN_101; // @[MuxLiteral.scala 48:10]
  wire [2:0] _GEN_103; // @[MuxLiteral.scala 48:10]
  wire [2:0] _T_235; // @[RegisterRouter.scala 59:16]
  wire  _T_236_bits_read; // @[Decoupled.scala 308:19 Decoupled.scala 309:14]
  wire  _T_236_valid; // @[Decoupled.scala 308:19 Decoupled.scala 310:15]
  wire  _T_239; // @[RegisterRouter.scala 65:29]
  Queue Queue ( // @[Decoupled.scala 287:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_read(Queue_io_enq_bits_read),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_extra(Queue_io_enq_bits_extra),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_read(Queue_io_deq_bits_read),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_extra(Queue_io_deq_bits_extra)
  );
  assign _T_3 = sels_0 == 3'h0; // @[Mux.scala 45:28]
  assign _GEN_7 = _T_3 & auto_stream_in_0_valid; // @[Mux.scala 45:41]
  assign _GEN_8 = _T_3 & auto_stream_out_0_ready; // @[Mux.scala 45:41]
  assign _T_4 = sels_0 == 3'h1; // @[Mux.scala 45:28]
  assign _GEN_12 = _T_4 ? auto_stream_in_1_bits_last : auto_stream_in_0_bits_last; // @[Mux.scala 45:41]
  assign _GEN_15 = _T_4 ? auto_stream_in_1_bits_data : auto_stream_in_0_bits_data; // @[Mux.scala 45:41]
  assign _GEN_16 = _T_4 ? auto_stream_in_1_valid : _GEN_7; // @[Mux.scala 45:41]
  assign _GEN_17 = _T_4 & auto_stream_out_0_ready; // @[Mux.scala 45:41]
  assign _T_5 = sels_0 == 3'h2; // @[Mux.scala 45:28]
  assign _GEN_21 = _T_5 ? auto_stream_in_2_bits_last : _GEN_12; // @[Mux.scala 45:41]
  assign _GEN_24 = _T_5 ? auto_stream_in_2_bits_data : _GEN_15; // @[Mux.scala 45:41]
  assign _GEN_25 = _T_5 ? auto_stream_in_2_valid : _GEN_16; // @[Mux.scala 45:41]
  assign _GEN_26 = _T_5 & auto_stream_out_0_ready; // @[Mux.scala 45:41]
  assign _T_6 = sels_0 == 3'h3; // @[Mux.scala 45:28]
  assign _GEN_30 = _T_6 ? 1'h0 : _GEN_21; // @[Mux.scala 45:41]
  assign _GEN_33 = _T_6 ? 32'hffffffff : _GEN_24; // @[Mux.scala 45:41]
  assign _GEN_34 = _T_6 | _GEN_25; // @[Mux.scala 45:41]
  assign _T_7 = sels_0 == 3'h4; // @[Mux.scala 45:28]
  assign _T_8 = sels_0 == sels_1; // @[Mux.scala 40:46]
  assign _T_10 = _T_8 ? 3'h5 : sels_1; // @[Mux.scala 41:29]
  assign _T_11 = _T_10 == 3'h0; // @[Mux.scala 45:28]
  assign _T_12 = _T_10 == 3'h1; // @[Mux.scala 45:28]
  assign _T_13 = _T_10 == 3'h2; // @[Mux.scala 45:28]
  assign _T_17 = auto_register_in_aw_valid & auto_register_in_w_valid; // @[RegisterRouter.scala 40:39]
  assign _T_18 = auto_register_in_ar_valid | _T_17; // @[RegisterRouter.scala 40:26]
  assign _T_19 = ~auto_register_in_ar_valid; // @[RegisterRouter.scala 42:29]
  assign _T_62_ready = Queue_io_enq_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 290:17]
  assign _T_26 = auto_register_in_ar_valid ? auto_register_in_ar_bits_addr : auto_register_in_aw_bits_addr; // @[RegisterRouter.scala 48:19]
  assign _T_66 = _T_26[3:2] & 2'h2; // @[RegisterRouter.scala 59:16]
  assign _T_68 = _T_66 == 2'h0; // @[RegisterRouter.scala 59:16]
  assign _T_20 = _T_62_ready & _T_19; // @[RegisterRouter.scala 42:26]
  assign _T_29 = 2'h1 << auto_register_in_ar_bits_size[0]; // @[OneHot.scala 65:12]
  assign _T_31 = _T_29 | 2'h1; // @[Misc.scala 200:81]
  assign _T_32 = auto_register_in_ar_bits_size >= 3'h2; // @[Misc.scala 204:21]
  assign _T_35 = ~auto_register_in_ar_bits_addr[1]; // @[Misc.scala 209:20]
  assign _T_37 = _T_31[1] & _T_35; // @[Misc.scala 213:38]
  assign _T_38 = _T_32 | _T_37; // @[Misc.scala 213:29]
  assign _T_40 = _T_31[1] & auto_register_in_ar_bits_addr[1]; // @[Misc.scala 213:38]
  assign _T_41 = _T_32 | _T_40; // @[Misc.scala 213:29]
  assign _T_44 = ~auto_register_in_ar_bits_addr[0]; // @[Misc.scala 209:20]
  assign _T_45 = _T_35 & _T_44; // @[Misc.scala 212:27]
  assign _T_46 = _T_31[0] & _T_45; // @[Misc.scala 213:38]
  assign _T_47 = _T_38 | _T_46; // @[Misc.scala 213:29]
  assign _T_48 = _T_35 & auto_register_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  assign _T_49 = _T_31[0] & _T_48; // @[Misc.scala 213:38]
  assign _T_50 = _T_38 | _T_49; // @[Misc.scala 213:29]
  assign _T_51 = auto_register_in_ar_bits_addr[1] & _T_44; // @[Misc.scala 212:27]
  assign _T_52 = _T_31[0] & _T_51; // @[Misc.scala 213:38]
  assign _T_53 = _T_41 | _T_52; // @[Misc.scala 213:29]
  assign _T_54 = auto_register_in_ar_bits_addr[1] & auto_register_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  assign _T_55 = _T_31[0] & _T_54; // @[Misc.scala 213:38]
  assign _T_56 = _T_41 | _T_55; // @[Misc.scala 213:29]
  assign _T_59 = {_T_56,_T_53,_T_50,_T_47}; // @[Cat.scala 29:58]
  assign _T_61 = auto_register_in_ar_valid ? _T_59 : auto_register_in_w_bits_strb; // @[RegisterRouter.scala 54:25]
  assign _T_80 = _T_61[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_82 = _T_61[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_84 = _T_61[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_86 = _T_61[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_89 = {_T_86,_T_84,_T_82,_T_80}; // @[Cat.scala 29:58]
  assign _T_108 = _T_89[2:0] == 3'h7; // @[RegisterRouter.scala 59:16]
  assign _T_161 = _T_18 & _T_62_ready; // @[RegisterRouter.scala 59:16]
  assign _T_155 = 2'h1 << _T_26[2]; // @[OneHot.scala 58:35]
  assign _T_178 = _T_161 & _T_19; // @[RegisterRouter.scala 59:16]
  assign _T_185 = _T_178 & _T_155[1]; // @[RegisterRouter.scala 59:16]
  assign _T_186 = _T_185 & _T_68; // @[RegisterRouter.scala 59:16]
  assign _T_115 = _T_186 & _T_108; // @[RegisterRouter.scala 59:16]
  assign _T_180 = _T_178 & _T_155[0]; // @[RegisterRouter.scala 59:16]
  assign _T_181 = _T_180 & _T_68; // @[RegisterRouter.scala 59:16]
  assign _T_138 = _T_181 & _T_108; // @[RegisterRouter.scala 59:16]
  assign _GEN_101 = _T_26[2] ? _T_68 : _T_68; // @[MuxLiteral.scala 48:10]
  assign _GEN_103 = _T_26[2] ? sels_1 : sels_0; // @[MuxLiteral.scala 48:10]
  assign _T_235 = _GEN_101 ? _GEN_103 : 3'h0; // @[RegisterRouter.scala 59:16]
  assign _T_236_bits_read = Queue_io_deq_bits_read; // @[Decoupled.scala 308:19 Decoupled.scala 309:14]
  assign _T_236_valid = Queue_io_deq_valid; // @[Decoupled.scala 308:19 Decoupled.scala 310:15]
  assign _T_239 = ~_T_236_bits_read; // @[RegisterRouter.scala 65:29]
  assign auto_register_in_aw_ready = _T_20 & auto_register_in_w_valid; // @[LazyModule.scala 173:31]
  assign auto_register_in_w_ready = _T_20 & auto_register_in_aw_valid; // @[LazyModule.scala 173:31]
  assign auto_register_in_b_valid = _T_236_valid & _T_239; // @[LazyModule.scala 173:31]
  assign auto_register_in_b_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_register_in_ar_ready = Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_register_in_r_valid = _T_236_valid & _T_236_bits_read; // @[LazyModule.scala 173:31]
  assign auto_register_in_r_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_register_in_r_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 173:31]
  assign auto_stream_in_2_ready = _T_13 | _GEN_26; // @[LazyModule.scala 173:31]
  assign auto_stream_in_1_ready = _T_12 | _GEN_17; // @[LazyModule.scala 173:31]
  assign auto_stream_in_0_ready = _T_11 | _GEN_8; // @[LazyModule.scala 173:31]
  assign auto_stream_out_0_valid = _T_7 | _GEN_34; // @[LazyModule.scala 173:49]
  assign auto_stream_out_0_bits_data = _T_7 ? 32'h0 : _GEN_33; // @[LazyModule.scala 173:49]
  assign auto_stream_out_0_bits_last = _T_7 ? 1'h0 : _GEN_30; // @[LazyModule.scala 173:49]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_register_in_ar_valid | _T_17; // @[Decoupled.scala 288:22]
  assign Queue_io_enq_bits_read = auto_register_in_ar_valid; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_data = {{29'd0}, _T_235}; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_extra = auto_register_in_ar_valid ? auto_register_in_ar_bits_id : auto_register_in_aw_bits_id; // @[Decoupled.scala 289:21]
  assign Queue_io_deq_ready = _T_236_bits_read ? auto_register_in_r_ready : auto_register_in_b_ready; // @[Decoupled.scala 311:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  sels_0 = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  sels_1 = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      sels_0 <= 3'h5;
    end else if (_T_138) begin
      sels_0 <= auto_register_in_w_bits_data[2:0];
    end
    if (reset) begin
      sels_1 <= 3'h5;
    end else if (_T_115) begin
      sels_1 <= auto_register_in_w_bits_data[2:0];
    end
  end
endmodule
module AXI4StreamMux_5(
  input         clock,
  input         reset,
  output        auto_register_in_aw_ready,
  input         auto_register_in_aw_valid,
  input         auto_register_in_aw_bits_id,
  input  [29:0] auto_register_in_aw_bits_addr,
  output        auto_register_in_w_ready,
  input         auto_register_in_w_valid,
  input  [31:0] auto_register_in_w_bits_data,
  input  [3:0]  auto_register_in_w_bits_strb,
  input         auto_register_in_b_ready,
  output        auto_register_in_b_valid,
  output        auto_register_in_b_bits_id,
  output        auto_register_in_ar_ready,
  input         auto_register_in_ar_valid,
  input         auto_register_in_ar_bits_id,
  input  [29:0] auto_register_in_ar_bits_addr,
  input  [2:0]  auto_register_in_ar_bits_size,
  input         auto_register_in_r_ready,
  output        auto_register_in_r_valid,
  output        auto_register_in_r_bits_id,
  output [31:0] auto_register_in_r_bits_data,
  output        auto_stream_in_ready,
  input         auto_stream_in_valid,
  input  [31:0] auto_stream_in_bits_data,
  input         auto_stream_in_bits_last,
  input         auto_stream_out_1_ready,
  output        auto_stream_out_1_valid,
  output [31:0] auto_stream_out_1_bits_data,
  output        auto_stream_out_1_bits_last
);
  wire  Queue_clock; // @[Decoupled.scala 287:21]
  wire  Queue_reset; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_read; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_enq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_extra; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_read; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_deq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_extra; // @[Decoupled.scala 287:21]
  reg  sels_0; // @[Mux.scala 32:23]
  reg [31:0] _RAND_0;
  reg  sels_1; // @[Mux.scala 32:23]
  reg [31:0] _RAND_1;
  wire  _T_3; // @[Mux.scala 45:28]
  wire  _T_4; // @[Mux.scala 40:46]
  wire  _T_6; // @[Mux.scala 41:29]
  wire  _T_7; // @[Mux.scala 45:28]
  wire  _T_9; // @[RegisterRouter.scala 40:39]
  wire  _T_10; // @[RegisterRouter.scala 40:26]
  wire  _T_11; // @[RegisterRouter.scala 42:29]
  wire  _T_54_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 290:17]
  wire [29:0] _T_18; // @[RegisterRouter.scala 48:19]
  wire [1:0] _T_58; // @[RegisterRouter.scala 59:16]
  wire  _T_60; // @[RegisterRouter.scala 59:16]
  wire  _T_12; // @[RegisterRouter.scala 42:26]
  wire [1:0] _T_21; // @[OneHot.scala 65:12]
  wire [1:0] _T_23; // @[Misc.scala 200:81]
  wire  _T_24; // @[Misc.scala 204:21]
  wire  _T_27; // @[Misc.scala 209:20]
  wire  _T_29; // @[Misc.scala 213:38]
  wire  _T_30; // @[Misc.scala 213:29]
  wire  _T_32; // @[Misc.scala 213:38]
  wire  _T_33; // @[Misc.scala 213:29]
  wire  _T_36; // @[Misc.scala 209:20]
  wire  _T_37; // @[Misc.scala 212:27]
  wire  _T_38; // @[Misc.scala 213:38]
  wire  _T_39; // @[Misc.scala 213:29]
  wire  _T_40; // @[Misc.scala 212:27]
  wire  _T_41; // @[Misc.scala 213:38]
  wire  _T_42; // @[Misc.scala 213:29]
  wire  _T_43; // @[Misc.scala 212:27]
  wire  _T_44; // @[Misc.scala 213:38]
  wire  _T_45; // @[Misc.scala 213:29]
  wire  _T_46; // @[Misc.scala 212:27]
  wire  _T_47; // @[Misc.scala 213:38]
  wire  _T_48; // @[Misc.scala 213:29]
  wire [3:0] _T_51; // @[Cat.scala 29:58]
  wire [3:0] _T_53; // @[RegisterRouter.scala 54:25]
  wire [7:0] _T_72; // @[Bitwise.scala 72:12]
  wire [7:0] _T_74; // @[Bitwise.scala 72:12]
  wire [7:0] _T_76; // @[Bitwise.scala 72:12]
  wire [7:0] _T_78; // @[Bitwise.scala 72:12]
  wire [31:0] _T_81; // @[Cat.scala 29:58]
  wire  _T_153; // @[RegisterRouter.scala 59:16]
  wire [1:0] _T_147; // @[OneHot.scala 58:35]
  wire  _T_170; // @[RegisterRouter.scala 59:16]
  wire  _T_177; // @[RegisterRouter.scala 59:16]
  wire  _T_178; // @[RegisterRouter.scala 59:16]
  wire  _T_107; // @[RegisterRouter.scala 59:16]
  wire  _GEN_18; // @[RegField.scala 134:88]
  wire  _T_172; // @[RegisterRouter.scala 59:16]
  wire  _T_173; // @[RegisterRouter.scala 59:16]
  wire  _T_130; // @[RegisterRouter.scala 59:16]
  wire  _GEN_19; // @[RegField.scala 134:88]
  wire  _GEN_29; // @[MuxLiteral.scala 48:10]
  wire  _GEN_31; // @[MuxLiteral.scala 48:10]
  wire  _T_227; // @[RegisterRouter.scala 59:16]
  wire  _T_228_bits_read; // @[Decoupled.scala 308:19 Decoupled.scala 309:14]
  wire  _T_228_valid; // @[Decoupled.scala 308:19 Decoupled.scala 310:15]
  wire  _T_231; // @[RegisterRouter.scala 65:29]
  Queue Queue ( // @[Decoupled.scala 287:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_read(Queue_io_enq_bits_read),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_extra(Queue_io_enq_bits_extra),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_read(Queue_io_deq_bits_read),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_extra(Queue_io_deq_bits_extra)
  );
  assign _T_3 = ~sels_0; // @[Mux.scala 45:28]
  assign _T_4 = sels_0 == sels_1; // @[Mux.scala 40:46]
  assign _T_6 = _T_4 | sels_1; // @[Mux.scala 41:29]
  assign _T_7 = ~_T_6; // @[Mux.scala 45:28]
  assign _T_9 = auto_register_in_aw_valid & auto_register_in_w_valid; // @[RegisterRouter.scala 40:39]
  assign _T_10 = auto_register_in_ar_valid | _T_9; // @[RegisterRouter.scala 40:26]
  assign _T_11 = ~auto_register_in_ar_valid; // @[RegisterRouter.scala 42:29]
  assign _T_54_ready = Queue_io_enq_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 290:17]
  assign _T_18 = auto_register_in_ar_valid ? auto_register_in_ar_bits_addr : auto_register_in_aw_bits_addr; // @[RegisterRouter.scala 48:19]
  assign _T_58 = _T_18[3:2] & 2'h2; // @[RegisterRouter.scala 59:16]
  assign _T_60 = _T_58 == 2'h0; // @[RegisterRouter.scala 59:16]
  assign _T_12 = _T_54_ready & _T_11; // @[RegisterRouter.scala 42:26]
  assign _T_21 = 2'h1 << auto_register_in_ar_bits_size[0]; // @[OneHot.scala 65:12]
  assign _T_23 = _T_21 | 2'h1; // @[Misc.scala 200:81]
  assign _T_24 = auto_register_in_ar_bits_size >= 3'h2; // @[Misc.scala 204:21]
  assign _T_27 = ~auto_register_in_ar_bits_addr[1]; // @[Misc.scala 209:20]
  assign _T_29 = _T_23[1] & _T_27; // @[Misc.scala 213:38]
  assign _T_30 = _T_24 | _T_29; // @[Misc.scala 213:29]
  assign _T_32 = _T_23[1] & auto_register_in_ar_bits_addr[1]; // @[Misc.scala 213:38]
  assign _T_33 = _T_24 | _T_32; // @[Misc.scala 213:29]
  assign _T_36 = ~auto_register_in_ar_bits_addr[0]; // @[Misc.scala 209:20]
  assign _T_37 = _T_27 & _T_36; // @[Misc.scala 212:27]
  assign _T_38 = _T_23[0] & _T_37; // @[Misc.scala 213:38]
  assign _T_39 = _T_30 | _T_38; // @[Misc.scala 213:29]
  assign _T_40 = _T_27 & auto_register_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  assign _T_41 = _T_23[0] & _T_40; // @[Misc.scala 213:38]
  assign _T_42 = _T_30 | _T_41; // @[Misc.scala 213:29]
  assign _T_43 = auto_register_in_ar_bits_addr[1] & _T_36; // @[Misc.scala 212:27]
  assign _T_44 = _T_23[0] & _T_43; // @[Misc.scala 213:38]
  assign _T_45 = _T_33 | _T_44; // @[Misc.scala 213:29]
  assign _T_46 = auto_register_in_ar_bits_addr[1] & auto_register_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  assign _T_47 = _T_23[0] & _T_46; // @[Misc.scala 213:38]
  assign _T_48 = _T_33 | _T_47; // @[Misc.scala 213:29]
  assign _T_51 = {_T_48,_T_45,_T_42,_T_39}; // @[Cat.scala 29:58]
  assign _T_53 = auto_register_in_ar_valid ? _T_51 : auto_register_in_w_bits_strb; // @[RegisterRouter.scala 54:25]
  assign _T_72 = _T_53[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_74 = _T_53[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_76 = _T_53[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_78 = _T_53[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_81 = {_T_78,_T_76,_T_74,_T_72}; // @[Cat.scala 29:58]
  assign _T_153 = _T_10 & _T_54_ready; // @[RegisterRouter.scala 59:16]
  assign _T_147 = 2'h1 << _T_18[2]; // @[OneHot.scala 58:35]
  assign _T_170 = _T_153 & _T_11; // @[RegisterRouter.scala 59:16]
  assign _T_177 = _T_170 & _T_147[1]; // @[RegisterRouter.scala 59:16]
  assign _T_178 = _T_177 & _T_60; // @[RegisterRouter.scala 59:16]
  assign _T_107 = _T_178 & _T_81[0]; // @[RegisterRouter.scala 59:16]
  assign _GEN_18 = _T_107 ? auto_register_in_w_bits_data[0] : sels_1; // @[RegField.scala 134:88]
  assign _T_172 = _T_170 & _T_147[0]; // @[RegisterRouter.scala 59:16]
  assign _T_173 = _T_172 & _T_60; // @[RegisterRouter.scala 59:16]
  assign _T_130 = _T_173 & _T_81[0]; // @[RegisterRouter.scala 59:16]
  assign _GEN_19 = _T_130 ? auto_register_in_w_bits_data[0] : sels_0; // @[RegField.scala 134:88]
  assign _GEN_29 = _T_18[2] ? _T_60 : _T_60; // @[MuxLiteral.scala 48:10]
  assign _GEN_31 = _T_18[2] ? sels_1 : sels_0; // @[MuxLiteral.scala 48:10]
  assign _T_227 = _GEN_29 & _GEN_31; // @[RegisterRouter.scala 59:16]
  assign _T_228_bits_read = Queue_io_deq_bits_read; // @[Decoupled.scala 308:19 Decoupled.scala 309:14]
  assign _T_228_valid = Queue_io_deq_valid; // @[Decoupled.scala 308:19 Decoupled.scala 310:15]
  assign _T_231 = ~_T_228_bits_read; // @[RegisterRouter.scala 65:29]
  assign auto_register_in_aw_ready = _T_12 & auto_register_in_w_valid; // @[LazyModule.scala 173:31]
  assign auto_register_in_w_ready = _T_12 & auto_register_in_aw_valid; // @[LazyModule.scala 173:31]
  assign auto_register_in_b_valid = _T_228_valid & _T_231; // @[LazyModule.scala 173:31]
  assign auto_register_in_b_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_register_in_ar_ready = Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_register_in_r_valid = _T_228_valid & _T_228_bits_read; // @[LazyModule.scala 173:31]
  assign auto_register_in_r_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_register_in_r_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 173:31]
  assign auto_stream_in_ready = _T_7 ? auto_stream_out_1_ready : _T_3; // @[LazyModule.scala 173:31]
  assign auto_stream_out_1_valid = _T_7 & auto_stream_in_valid; // @[LazyModule.scala 173:49]
  assign auto_stream_out_1_bits_data = auto_stream_in_bits_data; // @[LazyModule.scala 173:49]
  assign auto_stream_out_1_bits_last = auto_stream_in_bits_last; // @[LazyModule.scala 173:49]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_register_in_ar_valid | _T_9; // @[Decoupled.scala 288:22]
  assign Queue_io_enq_bits_read = auto_register_in_ar_valid; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_data = {{31'd0}, _T_227}; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_extra = auto_register_in_ar_valid ? auto_register_in_ar_bits_id : auto_register_in_aw_bits_id; // @[Decoupled.scala 289:21]
  assign Queue_io_deq_ready = _T_228_bits_read ? auto_register_in_r_ready : auto_register_in_b_ready; // @[Decoupled.scala 311:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  sels_0 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  sels_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    sels_0 <= reset | _GEN_19;
    sels_1 <= reset | _GEN_18;
  end
endmodule
module Queue_15(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [15:0] io_enq_bits_real,
  input  [15:0] io_enq_bits_imag,
  input         io_deq_ready,
  output        io_deq_valid,
  output [15:0] io_deq_bits_real,
  output [15:0] io_deq_bits_imag
);
  reg [15:0] _T_4_real [0:4]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_0;
  wire [15:0] _T_4_real__T_26_data; // @[Decoupled.scala 209:24]
  wire [2:0] _T_4_real__T_26_addr; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_1;
  wire [15:0] _T_4_real__T_16_data; // @[Decoupled.scala 209:24]
  wire [2:0] _T_4_real__T_16_addr; // @[Decoupled.scala 209:24]
  wire  _T_4_real__T_16_mask; // @[Decoupled.scala 209:24]
  wire  _T_4_real__T_16_en; // @[Decoupled.scala 209:24]
  reg [15:0] _T_4_imag [0:4]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_2;
  wire [15:0] _T_4_imag__T_26_data; // @[Decoupled.scala 209:24]
  wire [2:0] _T_4_imag__T_26_addr; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_3;
  wire [15:0] _T_4_imag__T_16_data; // @[Decoupled.scala 209:24]
  wire [2:0] _T_4_imag__T_16_addr; // @[Decoupled.scala 209:24]
  wire  _T_4_imag__T_16_mask; // @[Decoupled.scala 209:24]
  wire  _T_4_imag__T_16_en; // @[Decoupled.scala 209:24]
  reg [2:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_4;
  reg [2:0] value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  reg  _T_5; // @[Decoupled.scala 212:35]
  reg [31:0] _RAND_6;
  wire  _T_6; // @[Decoupled.scala 214:41]
  wire  _T_7; // @[Decoupled.scala 215:36]
  wire  _T_8; // @[Decoupled.scala 215:33]
  wire  _T_9; // @[Decoupled.scala 216:32]
  wire  _T_10; // @[Decoupled.scala 40:37]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  wrap; // @[Counter.scala 38:24]
  wire [2:0] _T_18; // @[Counter.scala 39:22]
  wire  wrap_1; // @[Counter.scala 38:24]
  wire [2:0] _T_20; // @[Counter.scala 39:22]
  wire  _T_21; // @[Decoupled.scala 227:16]
  assign _T_4_real__T_26_addr = value_1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_4_real__T_26_data = _T_4_real[_T_4_real__T_26_addr]; // @[Decoupled.scala 209:24]
  `else
  assign _T_4_real__T_26_data = _T_4_real__T_26_addr >= 3'h5 ? _RAND_1[15:0] : _T_4_real[_T_4_real__T_26_addr]; // @[Decoupled.scala 209:24]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_4_real__T_16_data = io_enq_bits_real;
  assign _T_4_real__T_16_addr = value;
  assign _T_4_real__T_16_mask = 1'h1;
  assign _T_4_real__T_16_en = io_enq_ready & io_enq_valid;
  assign _T_4_imag__T_26_addr = value_1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_4_imag__T_26_data = _T_4_imag[_T_4_imag__T_26_addr]; // @[Decoupled.scala 209:24]
  `else
  assign _T_4_imag__T_26_data = _T_4_imag__T_26_addr >= 3'h5 ? _RAND_3[15:0] : _T_4_imag[_T_4_imag__T_26_addr]; // @[Decoupled.scala 209:24]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_4_imag__T_16_data = io_enq_bits_imag;
  assign _T_4_imag__T_16_addr = value;
  assign _T_4_imag__T_16_mask = 1'h1;
  assign _T_4_imag__T_16_en = io_enq_ready & io_enq_valid;
  assign _T_6 = value == value_1; // @[Decoupled.scala 214:41]
  assign _T_7 = ~_T_5; // @[Decoupled.scala 215:36]
  assign _T_8 = _T_6 & _T_7; // @[Decoupled.scala 215:33]
  assign _T_9 = _T_6 & _T_5; // @[Decoupled.scala 216:32]
  assign _T_10 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  assign _T_12 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  assign wrap = value == 3'h4; // @[Counter.scala 38:24]
  assign _T_18 = value + 3'h1; // @[Counter.scala 39:22]
  assign wrap_1 = value_1 == 3'h4; // @[Counter.scala 38:24]
  assign _T_20 = value_1 + 3'h1; // @[Counter.scala 39:22]
  assign _T_21 = _T_10 != _T_12; // @[Decoupled.scala 227:16]
  assign io_enq_ready = ~_T_9; // @[Decoupled.scala 232:16]
  assign io_deq_valid = ~_T_8; // @[Decoupled.scala 231:16]
  assign io_deq_bits_real = _T_4_real__T_26_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_imag = _T_4_imag__T_26_data; // @[Decoupled.scala 233:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 5; initvar = initvar+1)
    _T_4_real[initvar] = _RAND_0[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  _RAND_2 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 5; initvar = initvar+1)
    _T_4_imag[initvar] = _RAND_2[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  value = _RAND_4[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value_1 = _RAND_5[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_5 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T_4_real__T_16_en & _T_4_real__T_16_mask) begin
      _T_4_real[_T_4_real__T_16_addr] <= _T_4_real__T_16_data; // @[Decoupled.scala 209:24]
    end
    if(_T_4_imag__T_16_en & _T_4_imag__T_16_mask) begin
      _T_4_imag[_T_4_imag__T_16_addr] <= _T_4_imag__T_16_data; // @[Decoupled.scala 209:24]
    end
    if (reset) begin
      value <= 3'h0;
    end else if (_T_10) begin
      if (wrap) begin
        value <= 3'h0;
      end else begin
        value <= _T_18;
      end
    end
    if (reset) begin
      value_1 <= 3'h0;
    end else if (_T_12) begin
      if (wrap_1) begin
        value_1 <= 3'h0;
      end else begin
        value_1 <= _T_20;
      end
    end
    if (reset) begin
      _T_5 <= 1'h0;
    end else if (_T_21) begin
      _T_5 <= _T_10;
    end
  end
endmodule
module Queue_16(
  input   clock,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input   io_enq_bits,
  input   io_deq_ready,
  output  io_deq_valid,
  output  io_deq_bits
);
  reg  _T [0:4]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_0;
  wire  _T__T_18_data; // @[Decoupled.scala 209:24]
  wire [2:0] _T__T_18_addr; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_1;
  wire  _T__T_10_data; // @[Decoupled.scala 209:24]
  wire [2:0] _T__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T__T_10_en; // @[Decoupled.scala 209:24]
  reg [2:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_2;
  reg [2:0] value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_3;
  reg  _T_1; // @[Decoupled.scala 212:35]
  reg [31:0] _RAND_4;
  wire  _T_2; // @[Decoupled.scala 214:41]
  wire  _T_3; // @[Decoupled.scala 215:36]
  wire  _T_4; // @[Decoupled.scala 215:33]
  wire  _T_5; // @[Decoupled.scala 216:32]
  wire  _T_6; // @[Decoupled.scala 40:37]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  wrap; // @[Counter.scala 38:24]
  wire [2:0] _T_12; // @[Counter.scala 39:22]
  wire  wrap_1; // @[Counter.scala 38:24]
  wire [2:0] _T_14; // @[Counter.scala 39:22]
  wire  _T_15; // @[Decoupled.scala 227:16]
  assign _T__T_18_addr = value_1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__T_18_data = _T[_T__T_18_addr]; // @[Decoupled.scala 209:24]
  `else
  assign _T__T_18_data = _T__T_18_addr >= 3'h5 ? _RAND_1[0:0] : _T[_T__T_18_addr]; // @[Decoupled.scala 209:24]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__T_10_data = io_enq_bits;
  assign _T__T_10_addr = value;
  assign _T__T_10_mask = 1'h1;
  assign _T__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_2 = value == value_1; // @[Decoupled.scala 214:41]
  assign _T_3 = ~_T_1; // @[Decoupled.scala 215:36]
  assign _T_4 = _T_2 & _T_3; // @[Decoupled.scala 215:33]
  assign _T_5 = _T_2 & _T_1; // @[Decoupled.scala 216:32]
  assign _T_6 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  assign _T_8 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  assign wrap = value == 3'h4; // @[Counter.scala 38:24]
  assign _T_12 = value + 3'h1; // @[Counter.scala 39:22]
  assign wrap_1 = value_1 == 3'h4; // @[Counter.scala 38:24]
  assign _T_14 = value_1 + 3'h1; // @[Counter.scala 39:22]
  assign _T_15 = _T_6 != _T_8; // @[Decoupled.scala 227:16]
  assign io_enq_ready = ~_T_5; // @[Decoupled.scala 232:16]
  assign io_deq_valid = ~_T_4; // @[Decoupled.scala 231:16]
  assign io_deq_bits = _T__T_18_data; // @[Decoupled.scala 233:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 5; initvar = initvar+1)
    _T[initvar] = _RAND_0[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  value = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  value_1 = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T__T_10_en & _T__T_10_mask) begin
      _T[_T__T_10_addr] <= _T__T_10_data; // @[Decoupled.scala 209:24]
    end
    if (reset) begin
      value <= 3'h0;
    end else if (_T_6) begin
      if (wrap) begin
        value <= 3'h0;
      end else begin
        value <= _T_12;
      end
    end
    if (reset) begin
      value_1 <= 3'h0;
    end else if (_T_8) begin
      if (wrap_1) begin
        value_1 <= 3'h0;
      end else begin
        value_1 <= _T_14;
      end
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else if (_T_15) begin
      _T_1 <= _T_6;
    end
  end
endmodule
module LogMagMux(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [15:0] io_in_bits_real,
  input  [15:0] io_in_bits_imag,
  input         io_lastIn,
  input         io_out_ready,
  output        io_out_valid,
  output [15:0] io_out_bits_real,
  output [15:0] io_out_bits_imag,
  input  [1:0]  io_sel,
  output        io_lastOut
);
  wire  Queue_clock; // @[Skid.scala 21:23]
  wire  Queue_reset; // @[Skid.scala 21:23]
  wire  Queue_io_enq_ready; // @[Skid.scala 21:23]
  wire  Queue_io_enq_valid; // @[Skid.scala 21:23]
  wire [15:0] Queue_io_enq_bits_real; // @[Skid.scala 21:23]
  wire [15:0] Queue_io_enq_bits_imag; // @[Skid.scala 21:23]
  wire  Queue_io_deq_ready; // @[Skid.scala 21:23]
  wire  Queue_io_deq_valid; // @[Skid.scala 21:23]
  wire [15:0] Queue_io_deq_bits_real; // @[Skid.scala 21:23]
  wire [15:0] Queue_io_deq_bits_imag; // @[Skid.scala 21:23]
  wire  Queue_1_clock; // @[Skid.scala 21:23]
  wire  Queue_1_reset; // @[Skid.scala 21:23]
  wire  Queue_1_io_enq_ready; // @[Skid.scala 21:23]
  wire  Queue_1_io_enq_valid; // @[Skid.scala 21:23]
  wire  Queue_1_io_enq_bits; // @[Skid.scala 21:23]
  wire  Queue_1_io_deq_ready; // @[Skid.scala 21:23]
  wire  Queue_1_io_deq_valid; // @[Skid.scala 21:23]
  wire  Queue_1_io_deq_bits; // @[Skid.scala 21:23]
  wire [15:0] _T_7; // @[FixedPointTypeClass.scala 30:68]
  wire [15:0] absInReal; // @[FixedPointTypeClass.scala 247:8]
  wire [15:0] _T_11; // @[FixedPointTypeClass.scala 30:68]
  wire [15:0] absInImag; // @[FixedPointTypeClass.scala 247:8]
  wire  _T_12; // @[FixedPointTypeClass.scala 55:59]
  wire [15:0] u; // @[Order.scala 56:31]
  wire  _T_13; // @[FixedPointTypeClass.scala 53:59]
  wire [15:0] v; // @[Order.scala 55:31]
  wire [12:0] _T_14; // @[FixedPointTypeClass.scala 117:50]
  wire [15:0] _GEN_559; // @[FixedPointTypeClass.scala 24:22]
  reg [16:0] _T_16; // @[Reg.scala 15:16]
  reg [31:0] _RAND_0;
  reg [16:0] jplMagOp1; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1;
  wire [12:0] _T_17; // @[FixedPointTypeClass.scala 117:50]
  wire [15:0] _GEN_560; // @[FixedPointTypeClass.scala 33:22]
  reg [16:0] tmpOp2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2;
  reg [14:0] _T_20; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3;
  wire [16:0] _GEN_561; // @[FixedPointTypeClass.scala 24:22]
  reg [17:0] jplMagOp2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4;
  reg [31:0] _T_23; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5;
  wire [32:0] _T_24; // @[FixedPointTypeClass.scala 153:43]
  reg [31:0] _T_26; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6;
  wire [32:0] _T_27; // @[FixedPointTypeClass.scala 153:43]
  reg [33:0] _T_29; // @[Reg.scala 15:16]
  reg [63:0] _RAND_7;
  reg [33:0] _T_30; // @[Reg.scala 15:16]
  reg [63:0] _RAND_8;
  reg [33:0] _T_31; // @[Reg.scala 15:16]
  reg [63:0] _RAND_9;
  wire [17:0] _GEN_562; // @[FixedPointTypeClass.scala 55:59]
  wire  _T_32; // @[FixedPointTypeClass.scala 55:59]
  reg [17:0] _T_33; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10;
  reg [17:0] jplMag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11;
  wire [17:0] _T_34; // @[LogMagMux.scala 113:35]
  wire  _T_37; // @[CircuitMath.scala 37:22]
  wire  _T_41; // @[CircuitMath.scala 37:22]
  wire  _T_44; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_48; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_49; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_53; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_54; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_55; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_56; // @[Cat.scala 29:58]
  wire  _T_59; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_63; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_64; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_68; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_69; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_70; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_71; // @[Cat.scala 29:58]
  wire [2:0] _T_72; // @[CircuitMath.scala 38:21]
  wire [3:0] _T_73; // @[Cat.scala 29:58]
  wire [3:0] _T_74; // @[CircuitMath.scala 38:21]
  wire [4:0] logUInt; // @[Cat.scala 29:58]
  wire [17:0] _T_589; // @[LogMagMux.scala 131:50]
  wire [31:0] _T_590; // @[UIntTypeClass.scala 124:39]
  reg [17:0] noLeadOne; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12;
  wire [4:0] _T_596; // @[LogMagMux.scala 132:44]
  reg [4:0] shiftNum; // @[Reg.scala 15:16]
  reg [31:0] _RAND_13;
  wire [48:0] _GEN_563; // @[UIntTypeClass.scala 124:39]
  wire [48:0] _T_599; // @[UIntTypeClass.scala 124:39]
  wire [8:0] logLookUpAddr; // @[LogMagMux.scala 134:74]
  wire [9:0] _GEN_15; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_16; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_17; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_18; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_19; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_20; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_21; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_22; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_23; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_24; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_25; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_26; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_27; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_28; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_29; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_30; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_31; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_32; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_33; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_34; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_35; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_36; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_37; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_38; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_39; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_40; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_41; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_42; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_43; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_44; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_45; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_46; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_47; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_48; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_49; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_50; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_51; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_52; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_53; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_54; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_55; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_56; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_57; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_58; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_59; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_60; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_61; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_62; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_63; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_64; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_65; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_66; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_67; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_68; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_69; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_70; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_71; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_72; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_73; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_74; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_75; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_76; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_77; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_78; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_79; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_80; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_81; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_82; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_83; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_84; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_85; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_86; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_87; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_88; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_89; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_90; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_91; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_92; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_93; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_94; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_95; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_96; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_97; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_98; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_99; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_100; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_101; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_102; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_103; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_104; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_105; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_106; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_107; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_108; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_109; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_110; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_111; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_112; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_113; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_114; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_115; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_116; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_117; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_118; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_119; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_120; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_121; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_122; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_123; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_124; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_125; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_126; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_127; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_128; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_129; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_130; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_131; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_132; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_133; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_134; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_135; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_136; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_137; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_138; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_139; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_140; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_141; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_142; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_143; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_144; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_145; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_146; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_147; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_148; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_149; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_150; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_151; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_152; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_153; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_154; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_155; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_156; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_157; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_158; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_159; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_160; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_161; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_162; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_163; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_164; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_165; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_166; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_167; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_168; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_169; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_170; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_171; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_172; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_173; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_174; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_175; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_176; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_177; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_178; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_179; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_180; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_181; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_182; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_183; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_184; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_185; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_186; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_187; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_188; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_189; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_190; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_191; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_192; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_193; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_194; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_195; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_196; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_197; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_198; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_199; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_200; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_201; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_202; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_203; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_204; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_205; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_206; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_207; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_208; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_209; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_210; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_211; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_212; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_213; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_214; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_215; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_216; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_217; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_218; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_219; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_220; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_221; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_222; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_223; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_224; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_225; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_226; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_227; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_228; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_229; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_230; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_231; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_232; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_233; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_234; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_235; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_236; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_237; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_238; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_239; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_240; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_241; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_242; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_243; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_244; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_245; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_246; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_247; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_248; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_249; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_250; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_251; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_252; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_253; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_254; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_255; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_256; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_257; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_258; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_259; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_260; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_261; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_262; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_263; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_264; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_265; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_266; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_267; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_268; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_269; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_270; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_271; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_272; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_273; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_274; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_275; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_276; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_277; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_278; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_279; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_280; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_281; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_282; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_283; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_284; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_285; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_286; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_287; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_288; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_289; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_290; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_291; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_292; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_293; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_294; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_295; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_296; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_297; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_298; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_299; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_300; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_301; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_302; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_303; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_304; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_305; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_306; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_307; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_308; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_309; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_310; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_311; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_312; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_313; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_314; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_315; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_316; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_317; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_318; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_319; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_320; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_321; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_322; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_323; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_324; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_325; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_326; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_327; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_328; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_329; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_330; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_331; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_332; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_333; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_334; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_335; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_336; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_337; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_338; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_339; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_340; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_341; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_342; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_343; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_344; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_345; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_346; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_347; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_348; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_349; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_350; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_351; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_352; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_353; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_354; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_355; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_356; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_357; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_358; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_359; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_360; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_361; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_362; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_363; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_364; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_365; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_366; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_367; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_368; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_369; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_370; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_371; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_372; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_373; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_374; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_375; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_376; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_377; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_378; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_379; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_380; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_381; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_382; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_383; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_384; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_385; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_386; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_387; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_388; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_389; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_390; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_391; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_392; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_393; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_394; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_395; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_396; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_397; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_398; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_399; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_400; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_401; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_402; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_403; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_404; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_405; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_406; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_407; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_408; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_409; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_410; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_411; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_412; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_413; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_414; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_415; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_416; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_417; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_418; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_419; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_420; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_421; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_422; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_423; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_424; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_425; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_426; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_427; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_428; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_429; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_430; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_431; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_432; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_433; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_434; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_435; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_436; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_437; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_438; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_439; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_440; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_441; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_442; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_443; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_444; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_445; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_446; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_447; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_448; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_449; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_450; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_451; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_452; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_453; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_454; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_455; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_456; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_457; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_458; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_459; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_460; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_461; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_462; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_463; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_464; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_465; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_466; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_467; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_468; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_469; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_470; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_471; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_472; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_473; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_474; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_475; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_476; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_477; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_478; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_479; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_480; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_481; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_482; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_483; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_484; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_485; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_486; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_487; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_488; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_489; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_490; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_491; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_492; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_493; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_494; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_495; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_496; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_497; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_498; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_499; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_500; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_501; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_502; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_503; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_504; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_505; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_506; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_507; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_508; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_509; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_510; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_511; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_512; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_513; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_514; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_515; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_516; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_517; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_518; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_519; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_520; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_521; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_522; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_523; // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_524; // @[LogMagMux.scala 136:11]
  wire [9:0] logFrac; // @[LogMagMux.scala 136:11]
  reg [4:0] _T_601; // @[Reg.scala 15:16]
  reg [31:0] _RAND_14;
  wire [13:0] _GEN_564; // @[LogMagMux.scala 141:91]
  wire [13:0] _GEN_565; // @[LogMagMux.scala 141:91]
  wire [13:0] _T_604; // @[LogMagMux.scala 141:91]
  wire [15:0] log2MagOut_imag; // @[LogMagMux.scala 160:38]
  reg [1:0] _T_614; // @[Reg.scala 15:16]
  reg [31:0] _RAND_15;
  reg [1:0] _T_615; // @[Reg.scala 15:16]
  reg [31:0] _RAND_16;
  reg [1:0] _T_616; // @[Reg.scala 15:16]
  reg [31:0] _RAND_17;
  reg [1:0] _T_617; // @[Reg.scala 15:16]
  reg [31:0] _RAND_18;
  reg [15:0] _T_620_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_19;
  reg [15:0] _T_620_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_20;
  reg [15:0] _T_623_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_21;
  reg [15:0] _T_623_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_22;
  reg [15:0] _T_626_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_23;
  reg [15:0] _T_626_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_24;
  reg [15:0] _T_629_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_25;
  reg [15:0] _T_629_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_26;
  wire  _T_630; // @[Mux.scala 68:19]
  wire [15:0] _T_633_real; // @[Mux.scala 68:16]
  wire [15:0] _T_633_imag; // @[Mux.scala 68:16]
  wire  _T_634; // @[Mux.scala 68:19]
  wire [15:0] _T_637_real; // @[Mux.scala 68:16]
  wire [15:0] jplMagOut_imag; // @[LogMagMux.scala 151:23 LogMagMux.scala 154:18]
  wire [15:0] _T_637_imag; // @[Mux.scala 68:16]
  wire  _T_638; // @[Mux.scala 68:19]
  wire [15:0] _T_641_real; // @[Mux.scala 68:16]
  wire [32:0] _GEN_567; // @[LogMagMux.scala 95:20 LogMagMux.scala 105:10]
  wire [15:0] magSqr; // @[LogMagMux.scala 95:20 LogMagMux.scala 105:10]
  wire [15:0] _T_641_imag; // @[Mux.scala 68:16]
  wire  _T_642; // @[Mux.scala 68:19]
  wire [15:0] output_mux_real; // @[Mux.scala 68:16]
  wire [15:0] output_mux_imag; // @[Mux.scala 68:16]
  wire  _T_645; // @[Decoupled.scala 40:37]
  reg  initialInDone; // @[LogMagMux.scala 187:30]
  reg [31:0] _RAND_27;
  reg [2:0] _T_653; // @[LogMagMux.scala 190:24]
  reg [31:0] _RAND_28;
  wire [2:0] _T_656; // @[LogMagMux.scala 193:22]
  wire  _T_657; // @[LogMagMux.scala 196:18]
  wire  _T_659; // @[LogMagMux.scala 196:39]
  wire  _GEN_544; // @[LogMagMux.scala 196:56]
  wire  _T_667; // @[Skid.scala 29:30]
  wire  _T_668; // @[Skid.scala 29:27]
  wire  skidInData_ready; // @[LogMagMux.scala 205:24 Skid.scala 29:14]
  wire  skidInData_valid; // @[LogMagMux.scala 205:24 LogMagMux.scala 207:20]
  wire  _T_662; // @[Decoupled.scala 40:37]
  reg  _T_663; // @[Reg.scala 27:20]
  reg [31:0] _RAND_29;
  reg  _T_664; // @[Reg.scala 27:20]
  reg [31:0] _RAND_30;
  reg  _T_665; // @[Reg.scala 27:20]
  reg [31:0] _RAND_31;
  reg  _T_666; // @[Reg.scala 27:20]
  reg [31:0] _RAND_32;
  reg  _T_673; // @[Reg.scala 15:16]
  reg [31:0] _RAND_33;
  reg  _T_674; // @[Reg.scala 15:16]
  reg [31:0] _RAND_34;
  reg  _T_675; // @[Reg.scala 15:16]
  reg [31:0] _RAND_35;
  reg  _T_676; // @[Reg.scala 15:16]
  reg [31:0] _RAND_36;
  wire  _T_677; // @[Decoupled.scala 40:37]
  reg  _T_678; // @[Reg.scala 27:20]
  reg [31:0] _RAND_37;
  reg  _T_679; // @[Reg.scala 27:20]
  reg [31:0] _RAND_38;
  reg  _T_680; // @[Reg.scala 27:20]
  reg [31:0] _RAND_39;
  reg  _T_681; // @[Reg.scala 27:20]
  reg [31:0] _RAND_40;
  wire [15:0] skidInData_bits_real; // @[LogMagMux.scala 205:24 LogMagMux.scala 206:19]
  wire [15:0] skidInData_bits_imag; // @[LogMagMux.scala 205:24 LogMagMux.scala 206:19]
  Queue_15 Queue ( // @[Skid.scala 21:23]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_real(Queue_io_enq_bits_real),
    .io_enq_bits_imag(Queue_io_enq_bits_imag),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_real(Queue_io_deq_bits_real),
    .io_deq_bits_imag(Queue_io_deq_bits_imag)
  );
  Queue_16 Queue_1 ( // @[Skid.scala 21:23]
    .clock(Queue_1_clock),
    .reset(Queue_1_reset),
    .io_enq_ready(Queue_1_io_enq_ready),
    .io_enq_valid(Queue_1_io_enq_valid),
    .io_enq_bits(Queue_1_io_enq_bits),
    .io_deq_ready(Queue_1_io_deq_ready),
    .io_deq_valid(Queue_1_io_deq_valid),
    .io_deq_bits(Queue_1_io_deq_bits)
  );
  assign _T_7 = 16'sh0 - $signed(io_in_bits_real); // @[FixedPointTypeClass.scala 30:68]
  assign absInReal = io_in_bits_real[15] ? $signed(_T_7) : $signed(io_in_bits_real); // @[FixedPointTypeClass.scala 247:8]
  assign _T_11 = 16'sh0 - $signed(io_in_bits_imag); // @[FixedPointTypeClass.scala 30:68]
  assign absInImag = io_in_bits_imag[15] ? $signed(_T_11) : $signed(io_in_bits_imag); // @[FixedPointTypeClass.scala 247:8]
  assign _T_12 = $signed(absInReal) > $signed(absInImag); // @[FixedPointTypeClass.scala 55:59]
  assign u = _T_12 ? $signed(absInReal) : $signed(absInImag); // @[Order.scala 56:31]
  assign _T_13 = $signed(absInReal) < $signed(absInImag); // @[FixedPointTypeClass.scala 53:59]
  assign v = _T_13 ? $signed(absInReal) : $signed(absInImag); // @[Order.scala 55:31]
  assign _T_14 = v[15:3]; // @[FixedPointTypeClass.scala 117:50]
  assign _GEN_559 = {{3{_T_14[12]}},_T_14}; // @[FixedPointTypeClass.scala 24:22]
  assign _T_17 = u[15:3]; // @[FixedPointTypeClass.scala 117:50]
  assign _GEN_560 = {{3{_T_17[12]}},_T_17}; // @[FixedPointTypeClass.scala 33:22]
  assign _GEN_561 = {{2{_T_20[14]}},_T_20}; // @[FixedPointTypeClass.scala 24:22]
  assign _T_24 = {$signed(_T_23), 1'h0}; // @[FixedPointTypeClass.scala 153:43]
  assign _T_27 = {$signed(_T_26), 1'h0}; // @[FixedPointTypeClass.scala 153:43]
  assign _GEN_562 = {{1{jplMagOp1[16]}},jplMagOp1}; // @[FixedPointTypeClass.scala 55:59]
  assign _T_32 = $signed(_GEN_562) > $signed(jplMagOp2); // @[FixedPointTypeClass.scala 55:59]
  assign _T_34 = jplMag; // @[LogMagMux.scala 113:35]
  assign _T_37 = _T_34[17:16] != 2'h0; // @[CircuitMath.scala 37:22]
  assign _T_41 = _T_34[15:8] != 8'h0; // @[CircuitMath.scala 37:22]
  assign _T_44 = _T_34[15:12] != 4'h0; // @[CircuitMath.scala 37:22]
  assign _T_48 = _T_34[14] ? 2'h2 : {{1'd0}, _T_34[13]}; // @[CircuitMath.scala 32:10]
  assign _T_49 = _T_34[15] ? 2'h3 : _T_48; // @[CircuitMath.scala 32:10]
  assign _T_53 = _T_34[10] ? 2'h2 : {{1'd0}, _T_34[9]}; // @[CircuitMath.scala 32:10]
  assign _T_54 = _T_34[11] ? 2'h3 : _T_53; // @[CircuitMath.scala 32:10]
  assign _T_55 = _T_44 ? _T_49 : _T_54; // @[CircuitMath.scala 38:21]
  assign _T_56 = {_T_44,_T_55}; // @[Cat.scala 29:58]
  assign _T_59 = _T_34[7:4] != 4'h0; // @[CircuitMath.scala 37:22]
  assign _T_63 = _T_34[6] ? 2'h2 : {{1'd0}, _T_34[5]}; // @[CircuitMath.scala 32:10]
  assign _T_64 = _T_34[7] ? 2'h3 : _T_63; // @[CircuitMath.scala 32:10]
  assign _T_68 = _T_34[2] ? 2'h2 : {{1'd0}, _T_34[1]}; // @[CircuitMath.scala 32:10]
  assign _T_69 = _T_34[3] ? 2'h3 : _T_68; // @[CircuitMath.scala 32:10]
  assign _T_70 = _T_59 ? _T_64 : _T_69; // @[CircuitMath.scala 38:21]
  assign _T_71 = {_T_59,_T_70}; // @[Cat.scala 29:58]
  assign _T_72 = _T_41 ? _T_56 : _T_71; // @[CircuitMath.scala 38:21]
  assign _T_73 = {_T_41,_T_72}; // @[Cat.scala 29:58]
  assign _T_74 = _T_37 ? {{3'd0}, _T_34[17]} : _T_73; // @[CircuitMath.scala 38:21]
  assign logUInt = {_T_37,_T_74}; // @[Cat.scala 29:58]
  assign _T_589 = _T_32 ? $signed({{1{jplMagOp1[16]}},jplMagOp1}) : $signed(jplMagOp2); // @[LogMagMux.scala 131:50]
  assign _T_590 = 32'h1 << logUInt; // @[UIntTypeClass.scala 124:39]
  assign _T_596 = 5'h10 - logUInt; // @[LogMagMux.scala 132:44]
  assign _GEN_563 = {{31'd0}, noLeadOne}; // @[UIntTypeClass.scala 124:39]
  assign _T_599 = _GEN_563 << shiftNum; // @[UIntTypeClass.scala 124:39]
  assign logLookUpAddr = _T_599[14:6]; // @[LogMagMux.scala 134:74]
  assign _GEN_15 = 9'h1 == logLookUpAddr ? $signed(10'sh1) : $signed(10'sh0); // @[LogMagMux.scala 136:11]
  assign _GEN_16 = 9'h2 == logLookUpAddr ? $signed(10'sh3) : $signed(_GEN_15); // @[LogMagMux.scala 136:11]
  assign _GEN_17 = 9'h3 == logLookUpAddr ? $signed(10'sh4) : $signed(_GEN_16); // @[LogMagMux.scala 136:11]
  assign _GEN_18 = 9'h4 == logLookUpAddr ? $signed(10'sh6) : $signed(_GEN_17); // @[LogMagMux.scala 136:11]
  assign _GEN_19 = 9'h5 == logLookUpAddr ? $signed(10'sh7) : $signed(_GEN_18); // @[LogMagMux.scala 136:11]
  assign _GEN_20 = 9'h6 == logLookUpAddr ? $signed(10'sh9) : $signed(_GEN_19); // @[LogMagMux.scala 136:11]
  assign _GEN_21 = 9'h7 == logLookUpAddr ? $signed(10'sha) : $signed(_GEN_20); // @[LogMagMux.scala 136:11]
  assign _GEN_22 = 9'h8 == logLookUpAddr ? $signed(10'shb) : $signed(_GEN_21); // @[LogMagMux.scala 136:11]
  assign _GEN_23 = 9'h9 == logLookUpAddr ? $signed(10'shd) : $signed(_GEN_22); // @[LogMagMux.scala 136:11]
  assign _GEN_24 = 9'ha == logLookUpAddr ? $signed(10'she) : $signed(_GEN_23); // @[LogMagMux.scala 136:11]
  assign _GEN_25 = 9'hb == logLookUpAddr ? $signed(10'sh10) : $signed(_GEN_24); // @[LogMagMux.scala 136:11]
  assign _GEN_26 = 9'hc == logLookUpAddr ? $signed(10'sh11) : $signed(_GEN_25); // @[LogMagMux.scala 136:11]
  assign _GEN_27 = 9'hd == logLookUpAddr ? $signed(10'sh13) : $signed(_GEN_26); // @[LogMagMux.scala 136:11]
  assign _GEN_28 = 9'he == logLookUpAddr ? $signed(10'sh14) : $signed(_GEN_27); // @[LogMagMux.scala 136:11]
  assign _GEN_29 = 9'hf == logLookUpAddr ? $signed(10'sh15) : $signed(_GEN_28); // @[LogMagMux.scala 136:11]
  assign _GEN_30 = 9'h10 == logLookUpAddr ? $signed(10'sh17) : $signed(_GEN_29); // @[LogMagMux.scala 136:11]
  assign _GEN_31 = 9'h11 == logLookUpAddr ? $signed(10'sh18) : $signed(_GEN_30); // @[LogMagMux.scala 136:11]
  assign _GEN_32 = 9'h12 == logLookUpAddr ? $signed(10'sh1a) : $signed(_GEN_31); // @[LogMagMux.scala 136:11]
  assign _GEN_33 = 9'h13 == logLookUpAddr ? $signed(10'sh1b) : $signed(_GEN_32); // @[LogMagMux.scala 136:11]
  assign _GEN_34 = 9'h14 == logLookUpAddr ? $signed(10'sh1c) : $signed(_GEN_33); // @[LogMagMux.scala 136:11]
  assign _GEN_35 = 9'h15 == logLookUpAddr ? $signed(10'sh1e) : $signed(_GEN_34); // @[LogMagMux.scala 136:11]
  assign _GEN_36 = 9'h16 == logLookUpAddr ? $signed(10'sh1f) : $signed(_GEN_35); // @[LogMagMux.scala 136:11]
  assign _GEN_37 = 9'h17 == logLookUpAddr ? $signed(10'sh20) : $signed(_GEN_36); // @[LogMagMux.scala 136:11]
  assign _GEN_38 = 9'h18 == logLookUpAddr ? $signed(10'sh22) : $signed(_GEN_37); // @[LogMagMux.scala 136:11]
  assign _GEN_39 = 9'h19 == logLookUpAddr ? $signed(10'sh23) : $signed(_GEN_38); // @[LogMagMux.scala 136:11]
  assign _GEN_40 = 9'h1a == logLookUpAddr ? $signed(10'sh25) : $signed(_GEN_39); // @[LogMagMux.scala 136:11]
  assign _GEN_41 = 9'h1b == logLookUpAddr ? $signed(10'sh26) : $signed(_GEN_40); // @[LogMagMux.scala 136:11]
  assign _GEN_42 = 9'h1c == logLookUpAddr ? $signed(10'sh27) : $signed(_GEN_41); // @[LogMagMux.scala 136:11]
  assign _GEN_43 = 9'h1d == logLookUpAddr ? $signed(10'sh29) : $signed(_GEN_42); // @[LogMagMux.scala 136:11]
  assign _GEN_44 = 9'h1e == logLookUpAddr ? $signed(10'sh2a) : $signed(_GEN_43); // @[LogMagMux.scala 136:11]
  assign _GEN_45 = 9'h1f == logLookUpAddr ? $signed(10'sh2b) : $signed(_GEN_44); // @[LogMagMux.scala 136:11]
  assign _GEN_46 = 9'h20 == logLookUpAddr ? $signed(10'sh2d) : $signed(_GEN_45); // @[LogMagMux.scala 136:11]
  assign _GEN_47 = 9'h21 == logLookUpAddr ? $signed(10'sh2e) : $signed(_GEN_46); // @[LogMagMux.scala 136:11]
  assign _GEN_48 = 9'h22 == logLookUpAddr ? $signed(10'sh2f) : $signed(_GEN_47); // @[LogMagMux.scala 136:11]
  assign _GEN_49 = 9'h23 == logLookUpAddr ? $signed(10'sh31) : $signed(_GEN_48); // @[LogMagMux.scala 136:11]
  assign _GEN_50 = 9'h24 == logLookUpAddr ? $signed(10'sh32) : $signed(_GEN_49); // @[LogMagMux.scala 136:11]
  assign _GEN_51 = 9'h25 == logLookUpAddr ? $signed(10'sh34) : $signed(_GEN_50); // @[LogMagMux.scala 136:11]
  assign _GEN_52 = 9'h26 == logLookUpAddr ? $signed(10'sh35) : $signed(_GEN_51); // @[LogMagMux.scala 136:11]
  assign _GEN_53 = 9'h27 == logLookUpAddr ? $signed(10'sh36) : $signed(_GEN_52); // @[LogMagMux.scala 136:11]
  assign _GEN_54 = 9'h28 == logLookUpAddr ? $signed(10'sh38) : $signed(_GEN_53); // @[LogMagMux.scala 136:11]
  assign _GEN_55 = 9'h29 == logLookUpAddr ? $signed(10'sh39) : $signed(_GEN_54); // @[LogMagMux.scala 136:11]
  assign _GEN_56 = 9'h2a == logLookUpAddr ? $signed(10'sh3a) : $signed(_GEN_55); // @[LogMagMux.scala 136:11]
  assign _GEN_57 = 9'h2b == logLookUpAddr ? $signed(10'sh3c) : $signed(_GEN_56); // @[LogMagMux.scala 136:11]
  assign _GEN_58 = 9'h2c == logLookUpAddr ? $signed(10'sh3d) : $signed(_GEN_57); // @[LogMagMux.scala 136:11]
  assign _GEN_59 = 9'h2d == logLookUpAddr ? $signed(10'sh3e) : $signed(_GEN_58); // @[LogMagMux.scala 136:11]
  assign _GEN_60 = 9'h2e == logLookUpAddr ? $signed(10'sh40) : $signed(_GEN_59); // @[LogMagMux.scala 136:11]
  assign _GEN_61 = 9'h2f == logLookUpAddr ? $signed(10'sh41) : $signed(_GEN_60); // @[LogMagMux.scala 136:11]
  assign _GEN_62 = 9'h30 == logLookUpAddr ? $signed(10'sh42) : $signed(_GEN_61); // @[LogMagMux.scala 136:11]
  assign _GEN_63 = 9'h31 == logLookUpAddr ? $signed(10'sh44) : $signed(_GEN_62); // @[LogMagMux.scala 136:11]
  assign _GEN_64 = 9'h32 == logLookUpAddr ? $signed(10'sh45) : $signed(_GEN_63); // @[LogMagMux.scala 136:11]
  assign _GEN_65 = 9'h33 == logLookUpAddr ? $signed(10'sh46) : $signed(_GEN_64); // @[LogMagMux.scala 136:11]
  assign _GEN_66 = 9'h34 == logLookUpAddr ? $signed(10'sh47) : $signed(_GEN_65); // @[LogMagMux.scala 136:11]
  assign _GEN_67 = 9'h35 == logLookUpAddr ? $signed(10'sh49) : $signed(_GEN_66); // @[LogMagMux.scala 136:11]
  assign _GEN_68 = 9'h36 == logLookUpAddr ? $signed(10'sh4a) : $signed(_GEN_67); // @[LogMagMux.scala 136:11]
  assign _GEN_69 = 9'h37 == logLookUpAddr ? $signed(10'sh4b) : $signed(_GEN_68); // @[LogMagMux.scala 136:11]
  assign _GEN_70 = 9'h38 == logLookUpAddr ? $signed(10'sh4d) : $signed(_GEN_69); // @[LogMagMux.scala 136:11]
  assign _GEN_71 = 9'h39 == logLookUpAddr ? $signed(10'sh4e) : $signed(_GEN_70); // @[LogMagMux.scala 136:11]
  assign _GEN_72 = 9'h3a == logLookUpAddr ? $signed(10'sh4f) : $signed(_GEN_71); // @[LogMagMux.scala 136:11]
  assign _GEN_73 = 9'h3b == logLookUpAddr ? $signed(10'sh51) : $signed(_GEN_72); // @[LogMagMux.scala 136:11]
  assign _GEN_74 = 9'h3c == logLookUpAddr ? $signed(10'sh52) : $signed(_GEN_73); // @[LogMagMux.scala 136:11]
  assign _GEN_75 = 9'h3d == logLookUpAddr ? $signed(10'sh53) : $signed(_GEN_74); // @[LogMagMux.scala 136:11]
  assign _GEN_76 = 9'h3e == logLookUpAddr ? $signed(10'sh54) : $signed(_GEN_75); // @[LogMagMux.scala 136:11]
  assign _GEN_77 = 9'h3f == logLookUpAddr ? $signed(10'sh56) : $signed(_GEN_76); // @[LogMagMux.scala 136:11]
  assign _GEN_78 = 9'h40 == logLookUpAddr ? $signed(10'sh57) : $signed(_GEN_77); // @[LogMagMux.scala 136:11]
  assign _GEN_79 = 9'h41 == logLookUpAddr ? $signed(10'sh58) : $signed(_GEN_78); // @[LogMagMux.scala 136:11]
  assign _GEN_80 = 9'h42 == logLookUpAddr ? $signed(10'sh5a) : $signed(_GEN_79); // @[LogMagMux.scala 136:11]
  assign _GEN_81 = 9'h43 == logLookUpAddr ? $signed(10'sh5b) : $signed(_GEN_80); // @[LogMagMux.scala 136:11]
  assign _GEN_82 = 9'h44 == logLookUpAddr ? $signed(10'sh5c) : $signed(_GEN_81); // @[LogMagMux.scala 136:11]
  assign _GEN_83 = 9'h45 == logLookUpAddr ? $signed(10'sh5d) : $signed(_GEN_82); // @[LogMagMux.scala 136:11]
  assign _GEN_84 = 9'h46 == logLookUpAddr ? $signed(10'sh5f) : $signed(_GEN_83); // @[LogMagMux.scala 136:11]
  assign _GEN_85 = 9'h47 == logLookUpAddr ? $signed(10'sh60) : $signed(_GEN_84); // @[LogMagMux.scala 136:11]
  assign _GEN_86 = 9'h48 == logLookUpAddr ? $signed(10'sh61) : $signed(_GEN_85); // @[LogMagMux.scala 136:11]
  assign _GEN_87 = 9'h49 == logLookUpAddr ? $signed(10'sh62) : $signed(_GEN_86); // @[LogMagMux.scala 136:11]
  assign _GEN_88 = 9'h4a == logLookUpAddr ? $signed(10'sh64) : $signed(_GEN_87); // @[LogMagMux.scala 136:11]
  assign _GEN_89 = 9'h4b == logLookUpAddr ? $signed(10'sh65) : $signed(_GEN_88); // @[LogMagMux.scala 136:11]
  assign _GEN_90 = 9'h4c == logLookUpAddr ? $signed(10'sh66) : $signed(_GEN_89); // @[LogMagMux.scala 136:11]
  assign _GEN_91 = 9'h4d == logLookUpAddr ? $signed(10'sh67) : $signed(_GEN_90); // @[LogMagMux.scala 136:11]
  assign _GEN_92 = 9'h4e == logLookUpAddr ? $signed(10'sh69) : $signed(_GEN_91); // @[LogMagMux.scala 136:11]
  assign _GEN_93 = 9'h4f == logLookUpAddr ? $signed(10'sh6a) : $signed(_GEN_92); // @[LogMagMux.scala 136:11]
  assign _GEN_94 = 9'h50 == logLookUpAddr ? $signed(10'sh6b) : $signed(_GEN_93); // @[LogMagMux.scala 136:11]
  assign _GEN_95 = 9'h51 == logLookUpAddr ? $signed(10'sh6c) : $signed(_GEN_94); // @[LogMagMux.scala 136:11]
  assign _GEN_96 = 9'h52 == logLookUpAddr ? $signed(10'sh6e) : $signed(_GEN_95); // @[LogMagMux.scala 136:11]
  assign _GEN_97 = 9'h53 == logLookUpAddr ? $signed(10'sh6f) : $signed(_GEN_96); // @[LogMagMux.scala 136:11]
  assign _GEN_98 = 9'h54 == logLookUpAddr ? $signed(10'sh70) : $signed(_GEN_97); // @[LogMagMux.scala 136:11]
  assign _GEN_99 = 9'h55 == logLookUpAddr ? $signed(10'sh71) : $signed(_GEN_98); // @[LogMagMux.scala 136:11]
  assign _GEN_100 = 9'h56 == logLookUpAddr ? $signed(10'sh73) : $signed(_GEN_99); // @[LogMagMux.scala 136:11]
  assign _GEN_101 = 9'h57 == logLookUpAddr ? $signed(10'sh74) : $signed(_GEN_100); // @[LogMagMux.scala 136:11]
  assign _GEN_102 = 9'h58 == logLookUpAddr ? $signed(10'sh75) : $signed(_GEN_101); // @[LogMagMux.scala 136:11]
  assign _GEN_103 = 9'h59 == logLookUpAddr ? $signed(10'sh76) : $signed(_GEN_102); // @[LogMagMux.scala 136:11]
  assign _GEN_104 = 9'h5a == logLookUpAddr ? $signed(10'sh78) : $signed(_GEN_103); // @[LogMagMux.scala 136:11]
  assign _GEN_105 = 9'h5b == logLookUpAddr ? $signed(10'sh79) : $signed(_GEN_104); // @[LogMagMux.scala 136:11]
  assign _GEN_106 = 9'h5c == logLookUpAddr ? $signed(10'sh7a) : $signed(_GEN_105); // @[LogMagMux.scala 136:11]
  assign _GEN_107 = 9'h5d == logLookUpAddr ? $signed(10'sh7b) : $signed(_GEN_106); // @[LogMagMux.scala 136:11]
  assign _GEN_108 = 9'h5e == logLookUpAddr ? $signed(10'sh7d) : $signed(_GEN_107); // @[LogMagMux.scala 136:11]
  assign _GEN_109 = 9'h5f == logLookUpAddr ? $signed(10'sh7e) : $signed(_GEN_108); // @[LogMagMux.scala 136:11]
  assign _GEN_110 = 9'h60 == logLookUpAddr ? $signed(10'sh7f) : $signed(_GEN_109); // @[LogMagMux.scala 136:11]
  assign _GEN_111 = 9'h61 == logLookUpAddr ? $signed(10'sh80) : $signed(_GEN_110); // @[LogMagMux.scala 136:11]
  assign _GEN_112 = 9'h62 == logLookUpAddr ? $signed(10'sh81) : $signed(_GEN_111); // @[LogMagMux.scala 136:11]
  assign _GEN_113 = 9'h63 == logLookUpAddr ? $signed(10'sh83) : $signed(_GEN_112); // @[LogMagMux.scala 136:11]
  assign _GEN_114 = 9'h64 == logLookUpAddr ? $signed(10'sh84) : $signed(_GEN_113); // @[LogMagMux.scala 136:11]
  assign _GEN_115 = 9'h65 == logLookUpAddr ? $signed(10'sh85) : $signed(_GEN_114); // @[LogMagMux.scala 136:11]
  assign _GEN_116 = 9'h66 == logLookUpAddr ? $signed(10'sh86) : $signed(_GEN_115); // @[LogMagMux.scala 136:11]
  assign _GEN_117 = 9'h67 == logLookUpAddr ? $signed(10'sh87) : $signed(_GEN_116); // @[LogMagMux.scala 136:11]
  assign _GEN_118 = 9'h68 == logLookUpAddr ? $signed(10'sh89) : $signed(_GEN_117); // @[LogMagMux.scala 136:11]
  assign _GEN_119 = 9'h69 == logLookUpAddr ? $signed(10'sh8a) : $signed(_GEN_118); // @[LogMagMux.scala 136:11]
  assign _GEN_120 = 9'h6a == logLookUpAddr ? $signed(10'sh8b) : $signed(_GEN_119); // @[LogMagMux.scala 136:11]
  assign _GEN_121 = 9'h6b == logLookUpAddr ? $signed(10'sh8c) : $signed(_GEN_120); // @[LogMagMux.scala 136:11]
  assign _GEN_122 = 9'h6c == logLookUpAddr ? $signed(10'sh8d) : $signed(_GEN_121); // @[LogMagMux.scala 136:11]
  assign _GEN_123 = 9'h6d == logLookUpAddr ? $signed(10'sh8f) : $signed(_GEN_122); // @[LogMagMux.scala 136:11]
  assign _GEN_124 = 9'h6e == logLookUpAddr ? $signed(10'sh90) : $signed(_GEN_123); // @[LogMagMux.scala 136:11]
  assign _GEN_125 = 9'h6f == logLookUpAddr ? $signed(10'sh91) : $signed(_GEN_124); // @[LogMagMux.scala 136:11]
  assign _GEN_126 = 9'h70 == logLookUpAddr ? $signed(10'sh92) : $signed(_GEN_125); // @[LogMagMux.scala 136:11]
  assign _GEN_127 = 9'h71 == logLookUpAddr ? $signed(10'sh93) : $signed(_GEN_126); // @[LogMagMux.scala 136:11]
  assign _GEN_128 = 9'h72 == logLookUpAddr ? $signed(10'sh94) : $signed(_GEN_127); // @[LogMagMux.scala 136:11]
  assign _GEN_129 = 9'h73 == logLookUpAddr ? $signed(10'sh96) : $signed(_GEN_128); // @[LogMagMux.scala 136:11]
  assign _GEN_130 = 9'h74 == logLookUpAddr ? $signed(10'sh97) : $signed(_GEN_129); // @[LogMagMux.scala 136:11]
  assign _GEN_131 = 9'h75 == logLookUpAddr ? $signed(10'sh98) : $signed(_GEN_130); // @[LogMagMux.scala 136:11]
  assign _GEN_132 = 9'h76 == logLookUpAddr ? $signed(10'sh99) : $signed(_GEN_131); // @[LogMagMux.scala 136:11]
  assign _GEN_133 = 9'h77 == logLookUpAddr ? $signed(10'sh9a) : $signed(_GEN_132); // @[LogMagMux.scala 136:11]
  assign _GEN_134 = 9'h78 == logLookUpAddr ? $signed(10'sh9c) : $signed(_GEN_133); // @[LogMagMux.scala 136:11]
  assign _GEN_135 = 9'h79 == logLookUpAddr ? $signed(10'sh9d) : $signed(_GEN_134); // @[LogMagMux.scala 136:11]
  assign _GEN_136 = 9'h7a == logLookUpAddr ? $signed(10'sh9e) : $signed(_GEN_135); // @[LogMagMux.scala 136:11]
  assign _GEN_137 = 9'h7b == logLookUpAddr ? $signed(10'sh9f) : $signed(_GEN_136); // @[LogMagMux.scala 136:11]
  assign _GEN_138 = 9'h7c == logLookUpAddr ? $signed(10'sha0) : $signed(_GEN_137); // @[LogMagMux.scala 136:11]
  assign _GEN_139 = 9'h7d == logLookUpAddr ? $signed(10'sha1) : $signed(_GEN_138); // @[LogMagMux.scala 136:11]
  assign _GEN_140 = 9'h7e == logLookUpAddr ? $signed(10'sha3) : $signed(_GEN_139); // @[LogMagMux.scala 136:11]
  assign _GEN_141 = 9'h7f == logLookUpAddr ? $signed(10'sha4) : $signed(_GEN_140); // @[LogMagMux.scala 136:11]
  assign _GEN_142 = 9'h80 == logLookUpAddr ? $signed(10'sha5) : $signed(_GEN_141); // @[LogMagMux.scala 136:11]
  assign _GEN_143 = 9'h81 == logLookUpAddr ? $signed(10'sha6) : $signed(_GEN_142); // @[LogMagMux.scala 136:11]
  assign _GEN_144 = 9'h82 == logLookUpAddr ? $signed(10'sha7) : $signed(_GEN_143); // @[LogMagMux.scala 136:11]
  assign _GEN_145 = 9'h83 == logLookUpAddr ? $signed(10'sha8) : $signed(_GEN_144); // @[LogMagMux.scala 136:11]
  assign _GEN_146 = 9'h84 == logLookUpAddr ? $signed(10'sha9) : $signed(_GEN_145); // @[LogMagMux.scala 136:11]
  assign _GEN_147 = 9'h85 == logLookUpAddr ? $signed(10'shab) : $signed(_GEN_146); // @[LogMagMux.scala 136:11]
  assign _GEN_148 = 9'h86 == logLookUpAddr ? $signed(10'shac) : $signed(_GEN_147); // @[LogMagMux.scala 136:11]
  assign _GEN_149 = 9'h87 == logLookUpAddr ? $signed(10'shad) : $signed(_GEN_148); // @[LogMagMux.scala 136:11]
  assign _GEN_150 = 9'h88 == logLookUpAddr ? $signed(10'shae) : $signed(_GEN_149); // @[LogMagMux.scala 136:11]
  assign _GEN_151 = 9'h89 == logLookUpAddr ? $signed(10'shaf) : $signed(_GEN_150); // @[LogMagMux.scala 136:11]
  assign _GEN_152 = 9'h8a == logLookUpAddr ? $signed(10'shb0) : $signed(_GEN_151); // @[LogMagMux.scala 136:11]
  assign _GEN_153 = 9'h8b == logLookUpAddr ? $signed(10'shb1) : $signed(_GEN_152); // @[LogMagMux.scala 136:11]
  assign _GEN_154 = 9'h8c == logLookUpAddr ? $signed(10'shb3) : $signed(_GEN_153); // @[LogMagMux.scala 136:11]
  assign _GEN_155 = 9'h8d == logLookUpAddr ? $signed(10'shb4) : $signed(_GEN_154); // @[LogMagMux.scala 136:11]
  assign _GEN_156 = 9'h8e == logLookUpAddr ? $signed(10'shb5) : $signed(_GEN_155); // @[LogMagMux.scala 136:11]
  assign _GEN_157 = 9'h8f == logLookUpAddr ? $signed(10'shb6) : $signed(_GEN_156); // @[LogMagMux.scala 136:11]
  assign _GEN_158 = 9'h90 == logLookUpAddr ? $signed(10'shb7) : $signed(_GEN_157); // @[LogMagMux.scala 136:11]
  assign _GEN_159 = 9'h91 == logLookUpAddr ? $signed(10'shb8) : $signed(_GEN_158); // @[LogMagMux.scala 136:11]
  assign _GEN_160 = 9'h92 == logLookUpAddr ? $signed(10'shb9) : $signed(_GEN_159); // @[LogMagMux.scala 136:11]
  assign _GEN_161 = 9'h93 == logLookUpAddr ? $signed(10'shba) : $signed(_GEN_160); // @[LogMagMux.scala 136:11]
  assign _GEN_162 = 9'h94 == logLookUpAddr ? $signed(10'shbc) : $signed(_GEN_161); // @[LogMagMux.scala 136:11]
  assign _GEN_163 = 9'h95 == logLookUpAddr ? $signed(10'shbd) : $signed(_GEN_162); // @[LogMagMux.scala 136:11]
  assign _GEN_164 = 9'h96 == logLookUpAddr ? $signed(10'shbe) : $signed(_GEN_163); // @[LogMagMux.scala 136:11]
  assign _GEN_165 = 9'h97 == logLookUpAddr ? $signed(10'shbf) : $signed(_GEN_164); // @[LogMagMux.scala 136:11]
  assign _GEN_166 = 9'h98 == logLookUpAddr ? $signed(10'shc0) : $signed(_GEN_165); // @[LogMagMux.scala 136:11]
  assign _GEN_167 = 9'h99 == logLookUpAddr ? $signed(10'shc1) : $signed(_GEN_166); // @[LogMagMux.scala 136:11]
  assign _GEN_168 = 9'h9a == logLookUpAddr ? $signed(10'shc2) : $signed(_GEN_167); // @[LogMagMux.scala 136:11]
  assign _GEN_169 = 9'h9b == logLookUpAddr ? $signed(10'shc3) : $signed(_GEN_168); // @[LogMagMux.scala 136:11]
  assign _GEN_170 = 9'h9c == logLookUpAddr ? $signed(10'shc4) : $signed(_GEN_169); // @[LogMagMux.scala 136:11]
  assign _GEN_171 = 9'h9d == logLookUpAddr ? $signed(10'shc6) : $signed(_GEN_170); // @[LogMagMux.scala 136:11]
  assign _GEN_172 = 9'h9e == logLookUpAddr ? $signed(10'shc7) : $signed(_GEN_171); // @[LogMagMux.scala 136:11]
  assign _GEN_173 = 9'h9f == logLookUpAddr ? $signed(10'shc8) : $signed(_GEN_172); // @[LogMagMux.scala 136:11]
  assign _GEN_174 = 9'ha0 == logLookUpAddr ? $signed(10'shc9) : $signed(_GEN_173); // @[LogMagMux.scala 136:11]
  assign _GEN_175 = 9'ha1 == logLookUpAddr ? $signed(10'shca) : $signed(_GEN_174); // @[LogMagMux.scala 136:11]
  assign _GEN_176 = 9'ha2 == logLookUpAddr ? $signed(10'shcb) : $signed(_GEN_175); // @[LogMagMux.scala 136:11]
  assign _GEN_177 = 9'ha3 == logLookUpAddr ? $signed(10'shcc) : $signed(_GEN_176); // @[LogMagMux.scala 136:11]
  assign _GEN_178 = 9'ha4 == logLookUpAddr ? $signed(10'shcd) : $signed(_GEN_177); // @[LogMagMux.scala 136:11]
  assign _GEN_179 = 9'ha5 == logLookUpAddr ? $signed(10'shce) : $signed(_GEN_178); // @[LogMagMux.scala 136:11]
  assign _GEN_180 = 9'ha6 == logLookUpAddr ? $signed(10'shcf) : $signed(_GEN_179); // @[LogMagMux.scala 136:11]
  assign _GEN_181 = 9'ha7 == logLookUpAddr ? $signed(10'shd1) : $signed(_GEN_180); // @[LogMagMux.scala 136:11]
  assign _GEN_182 = 9'ha8 == logLookUpAddr ? $signed(10'shd2) : $signed(_GEN_181); // @[LogMagMux.scala 136:11]
  assign _GEN_183 = 9'ha9 == logLookUpAddr ? $signed(10'shd3) : $signed(_GEN_182); // @[LogMagMux.scala 136:11]
  assign _GEN_184 = 9'haa == logLookUpAddr ? $signed(10'shd4) : $signed(_GEN_183); // @[LogMagMux.scala 136:11]
  assign _GEN_185 = 9'hab == logLookUpAddr ? $signed(10'shd5) : $signed(_GEN_184); // @[LogMagMux.scala 136:11]
  assign _GEN_186 = 9'hac == logLookUpAddr ? $signed(10'shd6) : $signed(_GEN_185); // @[LogMagMux.scala 136:11]
  assign _GEN_187 = 9'had == logLookUpAddr ? $signed(10'shd7) : $signed(_GEN_186); // @[LogMagMux.scala 136:11]
  assign _GEN_188 = 9'hae == logLookUpAddr ? $signed(10'shd8) : $signed(_GEN_187); // @[LogMagMux.scala 136:11]
  assign _GEN_189 = 9'haf == logLookUpAddr ? $signed(10'shd9) : $signed(_GEN_188); // @[LogMagMux.scala 136:11]
  assign _GEN_190 = 9'hb0 == logLookUpAddr ? $signed(10'shda) : $signed(_GEN_189); // @[LogMagMux.scala 136:11]
  assign _GEN_191 = 9'hb1 == logLookUpAddr ? $signed(10'shdb) : $signed(_GEN_190); // @[LogMagMux.scala 136:11]
  assign _GEN_192 = 9'hb2 == logLookUpAddr ? $signed(10'shdc) : $signed(_GEN_191); // @[LogMagMux.scala 136:11]
  assign _GEN_193 = 9'hb3 == logLookUpAddr ? $signed(10'shdd) : $signed(_GEN_192); // @[LogMagMux.scala 136:11]
  assign _GEN_194 = 9'hb4 == logLookUpAddr ? $signed(10'shdf) : $signed(_GEN_193); // @[LogMagMux.scala 136:11]
  assign _GEN_195 = 9'hb5 == logLookUpAddr ? $signed(10'she0) : $signed(_GEN_194); // @[LogMagMux.scala 136:11]
  assign _GEN_196 = 9'hb6 == logLookUpAddr ? $signed(10'she1) : $signed(_GEN_195); // @[LogMagMux.scala 136:11]
  assign _GEN_197 = 9'hb7 == logLookUpAddr ? $signed(10'she2) : $signed(_GEN_196); // @[LogMagMux.scala 136:11]
  assign _GEN_198 = 9'hb8 == logLookUpAddr ? $signed(10'she3) : $signed(_GEN_197); // @[LogMagMux.scala 136:11]
  assign _GEN_199 = 9'hb9 == logLookUpAddr ? $signed(10'she4) : $signed(_GEN_198); // @[LogMagMux.scala 136:11]
  assign _GEN_200 = 9'hba == logLookUpAddr ? $signed(10'she5) : $signed(_GEN_199); // @[LogMagMux.scala 136:11]
  assign _GEN_201 = 9'hbb == logLookUpAddr ? $signed(10'she6) : $signed(_GEN_200); // @[LogMagMux.scala 136:11]
  assign _GEN_202 = 9'hbc == logLookUpAddr ? $signed(10'she7) : $signed(_GEN_201); // @[LogMagMux.scala 136:11]
  assign _GEN_203 = 9'hbd == logLookUpAddr ? $signed(10'she8) : $signed(_GEN_202); // @[LogMagMux.scala 136:11]
  assign _GEN_204 = 9'hbe == logLookUpAddr ? $signed(10'she9) : $signed(_GEN_203); // @[LogMagMux.scala 136:11]
  assign _GEN_205 = 9'hbf == logLookUpAddr ? $signed(10'shea) : $signed(_GEN_204); // @[LogMagMux.scala 136:11]
  assign _GEN_206 = 9'hc0 == logLookUpAddr ? $signed(10'sheb) : $signed(_GEN_205); // @[LogMagMux.scala 136:11]
  assign _GEN_207 = 9'hc1 == logLookUpAddr ? $signed(10'shec) : $signed(_GEN_206); // @[LogMagMux.scala 136:11]
  assign _GEN_208 = 9'hc2 == logLookUpAddr ? $signed(10'shed) : $signed(_GEN_207); // @[LogMagMux.scala 136:11]
  assign _GEN_209 = 9'hc3 == logLookUpAddr ? $signed(10'shee) : $signed(_GEN_208); // @[LogMagMux.scala 136:11]
  assign _GEN_210 = 9'hc4 == logLookUpAddr ? $signed(10'shef) : $signed(_GEN_209); // @[LogMagMux.scala 136:11]
  assign _GEN_211 = 9'hc5 == logLookUpAddr ? $signed(10'shf0) : $signed(_GEN_210); // @[LogMagMux.scala 136:11]
  assign _GEN_212 = 9'hc6 == logLookUpAddr ? $signed(10'shf1) : $signed(_GEN_211); // @[LogMagMux.scala 136:11]
  assign _GEN_213 = 9'hc7 == logLookUpAddr ? $signed(10'shf3) : $signed(_GEN_212); // @[LogMagMux.scala 136:11]
  assign _GEN_214 = 9'hc8 == logLookUpAddr ? $signed(10'shf4) : $signed(_GEN_213); // @[LogMagMux.scala 136:11]
  assign _GEN_215 = 9'hc9 == logLookUpAddr ? $signed(10'shf5) : $signed(_GEN_214); // @[LogMagMux.scala 136:11]
  assign _GEN_216 = 9'hca == logLookUpAddr ? $signed(10'shf6) : $signed(_GEN_215); // @[LogMagMux.scala 136:11]
  assign _GEN_217 = 9'hcb == logLookUpAddr ? $signed(10'shf7) : $signed(_GEN_216); // @[LogMagMux.scala 136:11]
  assign _GEN_218 = 9'hcc == logLookUpAddr ? $signed(10'shf8) : $signed(_GEN_217); // @[LogMagMux.scala 136:11]
  assign _GEN_219 = 9'hcd == logLookUpAddr ? $signed(10'shf9) : $signed(_GEN_218); // @[LogMagMux.scala 136:11]
  assign _GEN_220 = 9'hce == logLookUpAddr ? $signed(10'shfa) : $signed(_GEN_219); // @[LogMagMux.scala 136:11]
  assign _GEN_221 = 9'hcf == logLookUpAddr ? $signed(10'shfb) : $signed(_GEN_220); // @[LogMagMux.scala 136:11]
  assign _GEN_222 = 9'hd0 == logLookUpAddr ? $signed(10'shfc) : $signed(_GEN_221); // @[LogMagMux.scala 136:11]
  assign _GEN_223 = 9'hd1 == logLookUpAddr ? $signed(10'shfd) : $signed(_GEN_222); // @[LogMagMux.scala 136:11]
  assign _GEN_224 = 9'hd2 == logLookUpAddr ? $signed(10'shfe) : $signed(_GEN_223); // @[LogMagMux.scala 136:11]
  assign _GEN_225 = 9'hd3 == logLookUpAddr ? $signed(10'shff) : $signed(_GEN_224); // @[LogMagMux.scala 136:11]
  assign _GEN_226 = 9'hd4 == logLookUpAddr ? $signed(10'sh100) : $signed(_GEN_225); // @[LogMagMux.scala 136:11]
  assign _GEN_227 = 9'hd5 == logLookUpAddr ? $signed(10'sh101) : $signed(_GEN_226); // @[LogMagMux.scala 136:11]
  assign _GEN_228 = 9'hd6 == logLookUpAddr ? $signed(10'sh102) : $signed(_GEN_227); // @[LogMagMux.scala 136:11]
  assign _GEN_229 = 9'hd7 == logLookUpAddr ? $signed(10'sh103) : $signed(_GEN_228); // @[LogMagMux.scala 136:11]
  assign _GEN_230 = 9'hd8 == logLookUpAddr ? $signed(10'sh104) : $signed(_GEN_229); // @[LogMagMux.scala 136:11]
  assign _GEN_231 = 9'hd9 == logLookUpAddr ? $signed(10'sh105) : $signed(_GEN_230); // @[LogMagMux.scala 136:11]
  assign _GEN_232 = 9'hda == logLookUpAddr ? $signed(10'sh106) : $signed(_GEN_231); // @[LogMagMux.scala 136:11]
  assign _GEN_233 = 9'hdb == logLookUpAddr ? $signed(10'sh107) : $signed(_GEN_232); // @[LogMagMux.scala 136:11]
  assign _GEN_234 = 9'hdc == logLookUpAddr ? $signed(10'sh108) : $signed(_GEN_233); // @[LogMagMux.scala 136:11]
  assign _GEN_235 = 9'hdd == logLookUpAddr ? $signed(10'sh109) : $signed(_GEN_234); // @[LogMagMux.scala 136:11]
  assign _GEN_236 = 9'hde == logLookUpAddr ? $signed(10'sh10a) : $signed(_GEN_235); // @[LogMagMux.scala 136:11]
  assign _GEN_237 = 9'hdf == logLookUpAddr ? $signed(10'sh10b) : $signed(_GEN_236); // @[LogMagMux.scala 136:11]
  assign _GEN_238 = 9'he0 == logLookUpAddr ? $signed(10'sh10c) : $signed(_GEN_237); // @[LogMagMux.scala 136:11]
  assign _GEN_239 = 9'he1 == logLookUpAddr ? $signed(10'sh10d) : $signed(_GEN_238); // @[LogMagMux.scala 136:11]
  assign _GEN_240 = 9'he2 == logLookUpAddr ? $signed(10'sh10e) : $signed(_GEN_239); // @[LogMagMux.scala 136:11]
  assign _GEN_241 = 9'he3 == logLookUpAddr ? $signed(10'sh10f) : $signed(_GEN_240); // @[LogMagMux.scala 136:11]
  assign _GEN_242 = 9'he4 == logLookUpAddr ? $signed(10'sh110) : $signed(_GEN_241); // @[LogMagMux.scala 136:11]
  assign _GEN_243 = 9'he5 == logLookUpAddr ? $signed(10'sh111) : $signed(_GEN_242); // @[LogMagMux.scala 136:11]
  assign _GEN_244 = 9'he6 == logLookUpAddr ? $signed(10'sh112) : $signed(_GEN_243); // @[LogMagMux.scala 136:11]
  assign _GEN_245 = 9'he7 == logLookUpAddr ? $signed(10'sh113) : $signed(_GEN_244); // @[LogMagMux.scala 136:11]
  assign _GEN_246 = 9'he8 == logLookUpAddr ? $signed(10'sh114) : $signed(_GEN_245); // @[LogMagMux.scala 136:11]
  assign _GEN_247 = 9'he9 == logLookUpAddr ? $signed(10'sh115) : $signed(_GEN_246); // @[LogMagMux.scala 136:11]
  assign _GEN_248 = 9'hea == logLookUpAddr ? $signed(10'sh116) : $signed(_GEN_247); // @[LogMagMux.scala 136:11]
  assign _GEN_249 = 9'heb == logLookUpAddr ? $signed(10'sh117) : $signed(_GEN_248); // @[LogMagMux.scala 136:11]
  assign _GEN_250 = 9'hec == logLookUpAddr ? $signed(10'sh118) : $signed(_GEN_249); // @[LogMagMux.scala 136:11]
  assign _GEN_251 = 9'hed == logLookUpAddr ? $signed(10'sh119) : $signed(_GEN_250); // @[LogMagMux.scala 136:11]
  assign _GEN_252 = 9'hee == logLookUpAddr ? $signed(10'sh11a) : $signed(_GEN_251); // @[LogMagMux.scala 136:11]
  assign _GEN_253 = 9'hef == logLookUpAddr ? $signed(10'sh11b) : $signed(_GEN_252); // @[LogMagMux.scala 136:11]
  assign _GEN_254 = 9'hf0 == logLookUpAddr ? $signed(10'sh11c) : $signed(_GEN_253); // @[LogMagMux.scala 136:11]
  assign _GEN_255 = 9'hf1 == logLookUpAddr ? $signed(10'sh11d) : $signed(_GEN_254); // @[LogMagMux.scala 136:11]
  assign _GEN_256 = 9'hf2 == logLookUpAddr ? $signed(10'sh11e) : $signed(_GEN_255); // @[LogMagMux.scala 136:11]
  assign _GEN_257 = 9'hf3 == logLookUpAddr ? $signed(10'sh11f) : $signed(_GEN_256); // @[LogMagMux.scala 136:11]
  assign _GEN_258 = 9'hf4 == logLookUpAddr ? $signed(10'sh120) : $signed(_GEN_257); // @[LogMagMux.scala 136:11]
  assign _GEN_259 = 9'hf5 == logLookUpAddr ? $signed(10'sh121) : $signed(_GEN_258); // @[LogMagMux.scala 136:11]
  assign _GEN_260 = 9'hf6 == logLookUpAddr ? $signed(10'sh122) : $signed(_GEN_259); // @[LogMagMux.scala 136:11]
  assign _GEN_261 = 9'hf7 == logLookUpAddr ? $signed(10'sh123) : $signed(_GEN_260); // @[LogMagMux.scala 136:11]
  assign _GEN_262 = 9'hf8 == logLookUpAddr ? $signed(10'sh124) : $signed(_GEN_261); // @[LogMagMux.scala 136:11]
  assign _GEN_263 = 9'hf9 == logLookUpAddr ? $signed(10'sh125) : $signed(_GEN_262); // @[LogMagMux.scala 136:11]
  assign _GEN_264 = 9'hfa == logLookUpAddr ? $signed(10'sh126) : $signed(_GEN_263); // @[LogMagMux.scala 136:11]
  assign _GEN_265 = 9'hfb == logLookUpAddr ? $signed(10'sh127) : $signed(_GEN_264); // @[LogMagMux.scala 136:11]
  assign _GEN_266 = 9'hfc == logLookUpAddr ? $signed(10'sh128) : $signed(_GEN_265); // @[LogMagMux.scala 136:11]
  assign _GEN_267 = 9'hfd == logLookUpAddr ? $signed(10'sh129) : $signed(_GEN_266); // @[LogMagMux.scala 136:11]
  assign _GEN_268 = 9'hfe == logLookUpAddr ? $signed(10'sh12a) : $signed(_GEN_267); // @[LogMagMux.scala 136:11]
  assign _GEN_269 = 9'hff == logLookUpAddr ? $signed(10'sh12b) : $signed(_GEN_268); // @[LogMagMux.scala 136:11]
  assign _GEN_270 = 9'h100 == logLookUpAddr ? $signed(10'sh12c) : $signed(_GEN_269); // @[LogMagMux.scala 136:11]
  assign _GEN_271 = 9'h101 == logLookUpAddr ? $signed(10'sh12c) : $signed(_GEN_270); // @[LogMagMux.scala 136:11]
  assign _GEN_272 = 9'h102 == logLookUpAddr ? $signed(10'sh12d) : $signed(_GEN_271); // @[LogMagMux.scala 136:11]
  assign _GEN_273 = 9'h103 == logLookUpAddr ? $signed(10'sh12e) : $signed(_GEN_272); // @[LogMagMux.scala 136:11]
  assign _GEN_274 = 9'h104 == logLookUpAddr ? $signed(10'sh12f) : $signed(_GEN_273); // @[LogMagMux.scala 136:11]
  assign _GEN_275 = 9'h105 == logLookUpAddr ? $signed(10'sh130) : $signed(_GEN_274); // @[LogMagMux.scala 136:11]
  assign _GEN_276 = 9'h106 == logLookUpAddr ? $signed(10'sh131) : $signed(_GEN_275); // @[LogMagMux.scala 136:11]
  assign _GEN_277 = 9'h107 == logLookUpAddr ? $signed(10'sh132) : $signed(_GEN_276); // @[LogMagMux.scala 136:11]
  assign _GEN_278 = 9'h108 == logLookUpAddr ? $signed(10'sh133) : $signed(_GEN_277); // @[LogMagMux.scala 136:11]
  assign _GEN_279 = 9'h109 == logLookUpAddr ? $signed(10'sh134) : $signed(_GEN_278); // @[LogMagMux.scala 136:11]
  assign _GEN_280 = 9'h10a == logLookUpAddr ? $signed(10'sh135) : $signed(_GEN_279); // @[LogMagMux.scala 136:11]
  assign _GEN_281 = 9'h10b == logLookUpAddr ? $signed(10'sh136) : $signed(_GEN_280); // @[LogMagMux.scala 136:11]
  assign _GEN_282 = 9'h10c == logLookUpAddr ? $signed(10'sh137) : $signed(_GEN_281); // @[LogMagMux.scala 136:11]
  assign _GEN_283 = 9'h10d == logLookUpAddr ? $signed(10'sh138) : $signed(_GEN_282); // @[LogMagMux.scala 136:11]
  assign _GEN_284 = 9'h10e == logLookUpAddr ? $signed(10'sh139) : $signed(_GEN_283); // @[LogMagMux.scala 136:11]
  assign _GEN_285 = 9'h10f == logLookUpAddr ? $signed(10'sh13a) : $signed(_GEN_284); // @[LogMagMux.scala 136:11]
  assign _GEN_286 = 9'h110 == logLookUpAddr ? $signed(10'sh13b) : $signed(_GEN_285); // @[LogMagMux.scala 136:11]
  assign _GEN_287 = 9'h111 == logLookUpAddr ? $signed(10'sh13c) : $signed(_GEN_286); // @[LogMagMux.scala 136:11]
  assign _GEN_288 = 9'h112 == logLookUpAddr ? $signed(10'sh13d) : $signed(_GEN_287); // @[LogMagMux.scala 136:11]
  assign _GEN_289 = 9'h113 == logLookUpAddr ? $signed(10'sh13e) : $signed(_GEN_288); // @[LogMagMux.scala 136:11]
  assign _GEN_290 = 9'h114 == logLookUpAddr ? $signed(10'sh13e) : $signed(_GEN_289); // @[LogMagMux.scala 136:11]
  assign _GEN_291 = 9'h115 == logLookUpAddr ? $signed(10'sh13f) : $signed(_GEN_290); // @[LogMagMux.scala 136:11]
  assign _GEN_292 = 9'h116 == logLookUpAddr ? $signed(10'sh140) : $signed(_GEN_291); // @[LogMagMux.scala 136:11]
  assign _GEN_293 = 9'h117 == logLookUpAddr ? $signed(10'sh141) : $signed(_GEN_292); // @[LogMagMux.scala 136:11]
  assign _GEN_294 = 9'h118 == logLookUpAddr ? $signed(10'sh142) : $signed(_GEN_293); // @[LogMagMux.scala 136:11]
  assign _GEN_295 = 9'h119 == logLookUpAddr ? $signed(10'sh143) : $signed(_GEN_294); // @[LogMagMux.scala 136:11]
  assign _GEN_296 = 9'h11a == logLookUpAddr ? $signed(10'sh144) : $signed(_GEN_295); // @[LogMagMux.scala 136:11]
  assign _GEN_297 = 9'h11b == logLookUpAddr ? $signed(10'sh145) : $signed(_GEN_296); // @[LogMagMux.scala 136:11]
  assign _GEN_298 = 9'h11c == logLookUpAddr ? $signed(10'sh146) : $signed(_GEN_297); // @[LogMagMux.scala 136:11]
  assign _GEN_299 = 9'h11d == logLookUpAddr ? $signed(10'sh147) : $signed(_GEN_298); // @[LogMagMux.scala 136:11]
  assign _GEN_300 = 9'h11e == logLookUpAddr ? $signed(10'sh148) : $signed(_GEN_299); // @[LogMagMux.scala 136:11]
  assign _GEN_301 = 9'h11f == logLookUpAddr ? $signed(10'sh149) : $signed(_GEN_300); // @[LogMagMux.scala 136:11]
  assign _GEN_302 = 9'h120 == logLookUpAddr ? $signed(10'sh14a) : $signed(_GEN_301); // @[LogMagMux.scala 136:11]
  assign _GEN_303 = 9'h121 == logLookUpAddr ? $signed(10'sh14b) : $signed(_GEN_302); // @[LogMagMux.scala 136:11]
  assign _GEN_304 = 9'h122 == logLookUpAddr ? $signed(10'sh14b) : $signed(_GEN_303); // @[LogMagMux.scala 136:11]
  assign _GEN_305 = 9'h123 == logLookUpAddr ? $signed(10'sh14c) : $signed(_GEN_304); // @[LogMagMux.scala 136:11]
  assign _GEN_306 = 9'h124 == logLookUpAddr ? $signed(10'sh14d) : $signed(_GEN_305); // @[LogMagMux.scala 136:11]
  assign _GEN_307 = 9'h125 == logLookUpAddr ? $signed(10'sh14e) : $signed(_GEN_306); // @[LogMagMux.scala 136:11]
  assign _GEN_308 = 9'h126 == logLookUpAddr ? $signed(10'sh14f) : $signed(_GEN_307); // @[LogMagMux.scala 136:11]
  assign _GEN_309 = 9'h127 == logLookUpAddr ? $signed(10'sh150) : $signed(_GEN_308); // @[LogMagMux.scala 136:11]
  assign _GEN_310 = 9'h128 == logLookUpAddr ? $signed(10'sh151) : $signed(_GEN_309); // @[LogMagMux.scala 136:11]
  assign _GEN_311 = 9'h129 == logLookUpAddr ? $signed(10'sh152) : $signed(_GEN_310); // @[LogMagMux.scala 136:11]
  assign _GEN_312 = 9'h12a == logLookUpAddr ? $signed(10'sh153) : $signed(_GEN_311); // @[LogMagMux.scala 136:11]
  assign _GEN_313 = 9'h12b == logLookUpAddr ? $signed(10'sh154) : $signed(_GEN_312); // @[LogMagMux.scala 136:11]
  assign _GEN_314 = 9'h12c == logLookUpAddr ? $signed(10'sh155) : $signed(_GEN_313); // @[LogMagMux.scala 136:11]
  assign _GEN_315 = 9'h12d == logLookUpAddr ? $signed(10'sh156) : $signed(_GEN_314); // @[LogMagMux.scala 136:11]
  assign _GEN_316 = 9'h12e == logLookUpAddr ? $signed(10'sh156) : $signed(_GEN_315); // @[LogMagMux.scala 136:11]
  assign _GEN_317 = 9'h12f == logLookUpAddr ? $signed(10'sh157) : $signed(_GEN_316); // @[LogMagMux.scala 136:11]
  assign _GEN_318 = 9'h130 == logLookUpAddr ? $signed(10'sh158) : $signed(_GEN_317); // @[LogMagMux.scala 136:11]
  assign _GEN_319 = 9'h131 == logLookUpAddr ? $signed(10'sh159) : $signed(_GEN_318); // @[LogMagMux.scala 136:11]
  assign _GEN_320 = 9'h132 == logLookUpAddr ? $signed(10'sh15a) : $signed(_GEN_319); // @[LogMagMux.scala 136:11]
  assign _GEN_321 = 9'h133 == logLookUpAddr ? $signed(10'sh15b) : $signed(_GEN_320); // @[LogMagMux.scala 136:11]
  assign _GEN_322 = 9'h134 == logLookUpAddr ? $signed(10'sh15c) : $signed(_GEN_321); // @[LogMagMux.scala 136:11]
  assign _GEN_323 = 9'h135 == logLookUpAddr ? $signed(10'sh15d) : $signed(_GEN_322); // @[LogMagMux.scala 136:11]
  assign _GEN_324 = 9'h136 == logLookUpAddr ? $signed(10'sh15e) : $signed(_GEN_323); // @[LogMagMux.scala 136:11]
  assign _GEN_325 = 9'h137 == logLookUpAddr ? $signed(10'sh15f) : $signed(_GEN_324); // @[LogMagMux.scala 136:11]
  assign _GEN_326 = 9'h138 == logLookUpAddr ? $signed(10'sh15f) : $signed(_GEN_325); // @[LogMagMux.scala 136:11]
  assign _GEN_327 = 9'h139 == logLookUpAddr ? $signed(10'sh160) : $signed(_GEN_326); // @[LogMagMux.scala 136:11]
  assign _GEN_328 = 9'h13a == logLookUpAddr ? $signed(10'sh161) : $signed(_GEN_327); // @[LogMagMux.scala 136:11]
  assign _GEN_329 = 9'h13b == logLookUpAddr ? $signed(10'sh162) : $signed(_GEN_328); // @[LogMagMux.scala 136:11]
  assign _GEN_330 = 9'h13c == logLookUpAddr ? $signed(10'sh163) : $signed(_GEN_329); // @[LogMagMux.scala 136:11]
  assign _GEN_331 = 9'h13d == logLookUpAddr ? $signed(10'sh164) : $signed(_GEN_330); // @[LogMagMux.scala 136:11]
  assign _GEN_332 = 9'h13e == logLookUpAddr ? $signed(10'sh165) : $signed(_GEN_331); // @[LogMagMux.scala 136:11]
  assign _GEN_333 = 9'h13f == logLookUpAddr ? $signed(10'sh166) : $signed(_GEN_332); // @[LogMagMux.scala 136:11]
  assign _GEN_334 = 9'h140 == logLookUpAddr ? $signed(10'sh167) : $signed(_GEN_333); // @[LogMagMux.scala 136:11]
  assign _GEN_335 = 9'h141 == logLookUpAddr ? $signed(10'sh168) : $signed(_GEN_334); // @[LogMagMux.scala 136:11]
  assign _GEN_336 = 9'h142 == logLookUpAddr ? $signed(10'sh168) : $signed(_GEN_335); // @[LogMagMux.scala 136:11]
  assign _GEN_337 = 9'h143 == logLookUpAddr ? $signed(10'sh169) : $signed(_GEN_336); // @[LogMagMux.scala 136:11]
  assign _GEN_338 = 9'h144 == logLookUpAddr ? $signed(10'sh16a) : $signed(_GEN_337); // @[LogMagMux.scala 136:11]
  assign _GEN_339 = 9'h145 == logLookUpAddr ? $signed(10'sh16b) : $signed(_GEN_338); // @[LogMagMux.scala 136:11]
  assign _GEN_340 = 9'h146 == logLookUpAddr ? $signed(10'sh16c) : $signed(_GEN_339); // @[LogMagMux.scala 136:11]
  assign _GEN_341 = 9'h147 == logLookUpAddr ? $signed(10'sh16d) : $signed(_GEN_340); // @[LogMagMux.scala 136:11]
  assign _GEN_342 = 9'h148 == logLookUpAddr ? $signed(10'sh16e) : $signed(_GEN_341); // @[LogMagMux.scala 136:11]
  assign _GEN_343 = 9'h149 == logLookUpAddr ? $signed(10'sh16f) : $signed(_GEN_342); // @[LogMagMux.scala 136:11]
  assign _GEN_344 = 9'h14a == logLookUpAddr ? $signed(10'sh16f) : $signed(_GEN_343); // @[LogMagMux.scala 136:11]
  assign _GEN_345 = 9'h14b == logLookUpAddr ? $signed(10'sh170) : $signed(_GEN_344); // @[LogMagMux.scala 136:11]
  assign _GEN_346 = 9'h14c == logLookUpAddr ? $signed(10'sh171) : $signed(_GEN_345); // @[LogMagMux.scala 136:11]
  assign _GEN_347 = 9'h14d == logLookUpAddr ? $signed(10'sh172) : $signed(_GEN_346); // @[LogMagMux.scala 136:11]
  assign _GEN_348 = 9'h14e == logLookUpAddr ? $signed(10'sh173) : $signed(_GEN_347); // @[LogMagMux.scala 136:11]
  assign _GEN_349 = 9'h14f == logLookUpAddr ? $signed(10'sh174) : $signed(_GEN_348); // @[LogMagMux.scala 136:11]
  assign _GEN_350 = 9'h150 == logLookUpAddr ? $signed(10'sh175) : $signed(_GEN_349); // @[LogMagMux.scala 136:11]
  assign _GEN_351 = 9'h151 == logLookUpAddr ? $signed(10'sh176) : $signed(_GEN_350); // @[LogMagMux.scala 136:11]
  assign _GEN_352 = 9'h152 == logLookUpAddr ? $signed(10'sh176) : $signed(_GEN_351); // @[LogMagMux.scala 136:11]
  assign _GEN_353 = 9'h153 == logLookUpAddr ? $signed(10'sh177) : $signed(_GEN_352); // @[LogMagMux.scala 136:11]
  assign _GEN_354 = 9'h154 == logLookUpAddr ? $signed(10'sh178) : $signed(_GEN_353); // @[LogMagMux.scala 136:11]
  assign _GEN_355 = 9'h155 == logLookUpAddr ? $signed(10'sh179) : $signed(_GEN_354); // @[LogMagMux.scala 136:11]
  assign _GEN_356 = 9'h156 == logLookUpAddr ? $signed(10'sh17a) : $signed(_GEN_355); // @[LogMagMux.scala 136:11]
  assign _GEN_357 = 9'h157 == logLookUpAddr ? $signed(10'sh17b) : $signed(_GEN_356); // @[LogMagMux.scala 136:11]
  assign _GEN_358 = 9'h158 == logLookUpAddr ? $signed(10'sh17c) : $signed(_GEN_357); // @[LogMagMux.scala 136:11]
  assign _GEN_359 = 9'h159 == logLookUpAddr ? $signed(10'sh17c) : $signed(_GEN_358); // @[LogMagMux.scala 136:11]
  assign _GEN_360 = 9'h15a == logLookUpAddr ? $signed(10'sh17d) : $signed(_GEN_359); // @[LogMagMux.scala 136:11]
  assign _GEN_361 = 9'h15b == logLookUpAddr ? $signed(10'sh17e) : $signed(_GEN_360); // @[LogMagMux.scala 136:11]
  assign _GEN_362 = 9'h15c == logLookUpAddr ? $signed(10'sh17f) : $signed(_GEN_361); // @[LogMagMux.scala 136:11]
  assign _GEN_363 = 9'h15d == logLookUpAddr ? $signed(10'sh180) : $signed(_GEN_362); // @[LogMagMux.scala 136:11]
  assign _GEN_364 = 9'h15e == logLookUpAddr ? $signed(10'sh181) : $signed(_GEN_363); // @[LogMagMux.scala 136:11]
  assign _GEN_365 = 9'h15f == logLookUpAddr ? $signed(10'sh182) : $signed(_GEN_364); // @[LogMagMux.scala 136:11]
  assign _GEN_366 = 9'h160 == logLookUpAddr ? $signed(10'sh183) : $signed(_GEN_365); // @[LogMagMux.scala 136:11]
  assign _GEN_367 = 9'h161 == logLookUpAddr ? $signed(10'sh183) : $signed(_GEN_366); // @[LogMagMux.scala 136:11]
  assign _GEN_368 = 9'h162 == logLookUpAddr ? $signed(10'sh184) : $signed(_GEN_367); // @[LogMagMux.scala 136:11]
  assign _GEN_369 = 9'h163 == logLookUpAddr ? $signed(10'sh185) : $signed(_GEN_368); // @[LogMagMux.scala 136:11]
  assign _GEN_370 = 9'h164 == logLookUpAddr ? $signed(10'sh186) : $signed(_GEN_369); // @[LogMagMux.scala 136:11]
  assign _GEN_371 = 9'h165 == logLookUpAddr ? $signed(10'sh187) : $signed(_GEN_370); // @[LogMagMux.scala 136:11]
  assign _GEN_372 = 9'h166 == logLookUpAddr ? $signed(10'sh188) : $signed(_GEN_371); // @[LogMagMux.scala 136:11]
  assign _GEN_373 = 9'h167 == logLookUpAddr ? $signed(10'sh188) : $signed(_GEN_372); // @[LogMagMux.scala 136:11]
  assign _GEN_374 = 9'h168 == logLookUpAddr ? $signed(10'sh189) : $signed(_GEN_373); // @[LogMagMux.scala 136:11]
  assign _GEN_375 = 9'h169 == logLookUpAddr ? $signed(10'sh18a) : $signed(_GEN_374); // @[LogMagMux.scala 136:11]
  assign _GEN_376 = 9'h16a == logLookUpAddr ? $signed(10'sh18b) : $signed(_GEN_375); // @[LogMagMux.scala 136:11]
  assign _GEN_377 = 9'h16b == logLookUpAddr ? $signed(10'sh18c) : $signed(_GEN_376); // @[LogMagMux.scala 136:11]
  assign _GEN_378 = 9'h16c == logLookUpAddr ? $signed(10'sh18d) : $signed(_GEN_377); // @[LogMagMux.scala 136:11]
  assign _GEN_379 = 9'h16d == logLookUpAddr ? $signed(10'sh18e) : $signed(_GEN_378); // @[LogMagMux.scala 136:11]
  assign _GEN_380 = 9'h16e == logLookUpAddr ? $signed(10'sh18e) : $signed(_GEN_379); // @[LogMagMux.scala 136:11]
  assign _GEN_381 = 9'h16f == logLookUpAddr ? $signed(10'sh18f) : $signed(_GEN_380); // @[LogMagMux.scala 136:11]
  assign _GEN_382 = 9'h170 == logLookUpAddr ? $signed(10'sh190) : $signed(_GEN_381); // @[LogMagMux.scala 136:11]
  assign _GEN_383 = 9'h171 == logLookUpAddr ? $signed(10'sh191) : $signed(_GEN_382); // @[LogMagMux.scala 136:11]
  assign _GEN_384 = 9'h172 == logLookUpAddr ? $signed(10'sh192) : $signed(_GEN_383); // @[LogMagMux.scala 136:11]
  assign _GEN_385 = 9'h173 == logLookUpAddr ? $signed(10'sh193) : $signed(_GEN_384); // @[LogMagMux.scala 136:11]
  assign _GEN_386 = 9'h174 == logLookUpAddr ? $signed(10'sh193) : $signed(_GEN_385); // @[LogMagMux.scala 136:11]
  assign _GEN_387 = 9'h175 == logLookUpAddr ? $signed(10'sh194) : $signed(_GEN_386); // @[LogMagMux.scala 136:11]
  assign _GEN_388 = 9'h176 == logLookUpAddr ? $signed(10'sh195) : $signed(_GEN_387); // @[LogMagMux.scala 136:11]
  assign _GEN_389 = 9'h177 == logLookUpAddr ? $signed(10'sh196) : $signed(_GEN_388); // @[LogMagMux.scala 136:11]
  assign _GEN_390 = 9'h178 == logLookUpAddr ? $signed(10'sh197) : $signed(_GEN_389); // @[LogMagMux.scala 136:11]
  assign _GEN_391 = 9'h179 == logLookUpAddr ? $signed(10'sh198) : $signed(_GEN_390); // @[LogMagMux.scala 136:11]
  assign _GEN_392 = 9'h17a == logLookUpAddr ? $signed(10'sh198) : $signed(_GEN_391); // @[LogMagMux.scala 136:11]
  assign _GEN_393 = 9'h17b == logLookUpAddr ? $signed(10'sh199) : $signed(_GEN_392); // @[LogMagMux.scala 136:11]
  assign _GEN_394 = 9'h17c == logLookUpAddr ? $signed(10'sh19a) : $signed(_GEN_393); // @[LogMagMux.scala 136:11]
  assign _GEN_395 = 9'h17d == logLookUpAddr ? $signed(10'sh19b) : $signed(_GEN_394); // @[LogMagMux.scala 136:11]
  assign _GEN_396 = 9'h17e == logLookUpAddr ? $signed(10'sh19c) : $signed(_GEN_395); // @[LogMagMux.scala 136:11]
  assign _GEN_397 = 9'h17f == logLookUpAddr ? $signed(10'sh19d) : $signed(_GEN_396); // @[LogMagMux.scala 136:11]
  assign _GEN_398 = 9'h180 == logLookUpAddr ? $signed(10'sh19d) : $signed(_GEN_397); // @[LogMagMux.scala 136:11]
  assign _GEN_399 = 9'h181 == logLookUpAddr ? $signed(10'sh19e) : $signed(_GEN_398); // @[LogMagMux.scala 136:11]
  assign _GEN_400 = 9'h182 == logLookUpAddr ? $signed(10'sh19f) : $signed(_GEN_399); // @[LogMagMux.scala 136:11]
  assign _GEN_401 = 9'h183 == logLookUpAddr ? $signed(10'sh1a0) : $signed(_GEN_400); // @[LogMagMux.scala 136:11]
  assign _GEN_402 = 9'h184 == logLookUpAddr ? $signed(10'sh1a1) : $signed(_GEN_401); // @[LogMagMux.scala 136:11]
  assign _GEN_403 = 9'h185 == logLookUpAddr ? $signed(10'sh1a1) : $signed(_GEN_402); // @[LogMagMux.scala 136:11]
  assign _GEN_404 = 9'h186 == logLookUpAddr ? $signed(10'sh1a2) : $signed(_GEN_403); // @[LogMagMux.scala 136:11]
  assign _GEN_405 = 9'h187 == logLookUpAddr ? $signed(10'sh1a3) : $signed(_GEN_404); // @[LogMagMux.scala 136:11]
  assign _GEN_406 = 9'h188 == logLookUpAddr ? $signed(10'sh1a4) : $signed(_GEN_405); // @[LogMagMux.scala 136:11]
  assign _GEN_407 = 9'h189 == logLookUpAddr ? $signed(10'sh1a5) : $signed(_GEN_406); // @[LogMagMux.scala 136:11]
  assign _GEN_408 = 9'h18a == logLookUpAddr ? $signed(10'sh1a6) : $signed(_GEN_407); // @[LogMagMux.scala 136:11]
  assign _GEN_409 = 9'h18b == logLookUpAddr ? $signed(10'sh1a6) : $signed(_GEN_408); // @[LogMagMux.scala 136:11]
  assign _GEN_410 = 9'h18c == logLookUpAddr ? $signed(10'sh1a7) : $signed(_GEN_409); // @[LogMagMux.scala 136:11]
  assign _GEN_411 = 9'h18d == logLookUpAddr ? $signed(10'sh1a8) : $signed(_GEN_410); // @[LogMagMux.scala 136:11]
  assign _GEN_412 = 9'h18e == logLookUpAddr ? $signed(10'sh1a9) : $signed(_GEN_411); // @[LogMagMux.scala 136:11]
  assign _GEN_413 = 9'h18f == logLookUpAddr ? $signed(10'sh1aa) : $signed(_GEN_412); // @[LogMagMux.scala 136:11]
  assign _GEN_414 = 9'h190 == logLookUpAddr ? $signed(10'sh1aa) : $signed(_GEN_413); // @[LogMagMux.scala 136:11]
  assign _GEN_415 = 9'h191 == logLookUpAddr ? $signed(10'sh1ab) : $signed(_GEN_414); // @[LogMagMux.scala 136:11]
  assign _GEN_416 = 9'h192 == logLookUpAddr ? $signed(10'sh1ac) : $signed(_GEN_415); // @[LogMagMux.scala 136:11]
  assign _GEN_417 = 9'h193 == logLookUpAddr ? $signed(10'sh1ad) : $signed(_GEN_416); // @[LogMagMux.scala 136:11]
  assign _GEN_418 = 9'h194 == logLookUpAddr ? $signed(10'sh1ae) : $signed(_GEN_417); // @[LogMagMux.scala 136:11]
  assign _GEN_419 = 9'h195 == logLookUpAddr ? $signed(10'sh1ae) : $signed(_GEN_418); // @[LogMagMux.scala 136:11]
  assign _GEN_420 = 9'h196 == logLookUpAddr ? $signed(10'sh1af) : $signed(_GEN_419); // @[LogMagMux.scala 136:11]
  assign _GEN_421 = 9'h197 == logLookUpAddr ? $signed(10'sh1b0) : $signed(_GEN_420); // @[LogMagMux.scala 136:11]
  assign _GEN_422 = 9'h198 == logLookUpAddr ? $signed(10'sh1b1) : $signed(_GEN_421); // @[LogMagMux.scala 136:11]
  assign _GEN_423 = 9'h199 == logLookUpAddr ? $signed(10'sh1b2) : $signed(_GEN_422); // @[LogMagMux.scala 136:11]
  assign _GEN_424 = 9'h19a == logLookUpAddr ? $signed(10'sh1b2) : $signed(_GEN_423); // @[LogMagMux.scala 136:11]
  assign _GEN_425 = 9'h19b == logLookUpAddr ? $signed(10'sh1b3) : $signed(_GEN_424); // @[LogMagMux.scala 136:11]
  assign _GEN_426 = 9'h19c == logLookUpAddr ? $signed(10'sh1b4) : $signed(_GEN_425); // @[LogMagMux.scala 136:11]
  assign _GEN_427 = 9'h19d == logLookUpAddr ? $signed(10'sh1b5) : $signed(_GEN_426); // @[LogMagMux.scala 136:11]
  assign _GEN_428 = 9'h19e == logLookUpAddr ? $signed(10'sh1b6) : $signed(_GEN_427); // @[LogMagMux.scala 136:11]
  assign _GEN_429 = 9'h19f == logLookUpAddr ? $signed(10'sh1b6) : $signed(_GEN_428); // @[LogMagMux.scala 136:11]
  assign _GEN_430 = 9'h1a0 == logLookUpAddr ? $signed(10'sh1b7) : $signed(_GEN_429); // @[LogMagMux.scala 136:11]
  assign _GEN_431 = 9'h1a1 == logLookUpAddr ? $signed(10'sh1b8) : $signed(_GEN_430); // @[LogMagMux.scala 136:11]
  assign _GEN_432 = 9'h1a2 == logLookUpAddr ? $signed(10'sh1b9) : $signed(_GEN_431); // @[LogMagMux.scala 136:11]
  assign _GEN_433 = 9'h1a3 == logLookUpAddr ? $signed(10'sh1ba) : $signed(_GEN_432); // @[LogMagMux.scala 136:11]
  assign _GEN_434 = 9'h1a4 == logLookUpAddr ? $signed(10'sh1ba) : $signed(_GEN_433); // @[LogMagMux.scala 136:11]
  assign _GEN_435 = 9'h1a5 == logLookUpAddr ? $signed(10'sh1bb) : $signed(_GEN_434); // @[LogMagMux.scala 136:11]
  assign _GEN_436 = 9'h1a6 == logLookUpAddr ? $signed(10'sh1bc) : $signed(_GEN_435); // @[LogMagMux.scala 136:11]
  assign _GEN_437 = 9'h1a7 == logLookUpAddr ? $signed(10'sh1bd) : $signed(_GEN_436); // @[LogMagMux.scala 136:11]
  assign _GEN_438 = 9'h1a8 == logLookUpAddr ? $signed(10'sh1be) : $signed(_GEN_437); // @[LogMagMux.scala 136:11]
  assign _GEN_439 = 9'h1a9 == logLookUpAddr ? $signed(10'sh1be) : $signed(_GEN_438); // @[LogMagMux.scala 136:11]
  assign _GEN_440 = 9'h1aa == logLookUpAddr ? $signed(10'sh1bf) : $signed(_GEN_439); // @[LogMagMux.scala 136:11]
  assign _GEN_441 = 9'h1ab == logLookUpAddr ? $signed(10'sh1c0) : $signed(_GEN_440); // @[LogMagMux.scala 136:11]
  assign _GEN_442 = 9'h1ac == logLookUpAddr ? $signed(10'sh1c1) : $signed(_GEN_441); // @[LogMagMux.scala 136:11]
  assign _GEN_443 = 9'h1ad == logLookUpAddr ? $signed(10'sh1c2) : $signed(_GEN_442); // @[LogMagMux.scala 136:11]
  assign _GEN_444 = 9'h1ae == logLookUpAddr ? $signed(10'sh1c2) : $signed(_GEN_443); // @[LogMagMux.scala 136:11]
  assign _GEN_445 = 9'h1af == logLookUpAddr ? $signed(10'sh1c3) : $signed(_GEN_444); // @[LogMagMux.scala 136:11]
  assign _GEN_446 = 9'h1b0 == logLookUpAddr ? $signed(10'sh1c4) : $signed(_GEN_445); // @[LogMagMux.scala 136:11]
  assign _GEN_447 = 9'h1b1 == logLookUpAddr ? $signed(10'sh1c5) : $signed(_GEN_446); // @[LogMagMux.scala 136:11]
  assign _GEN_448 = 9'h1b2 == logLookUpAddr ? $signed(10'sh1c5) : $signed(_GEN_447); // @[LogMagMux.scala 136:11]
  assign _GEN_449 = 9'h1b3 == logLookUpAddr ? $signed(10'sh1c6) : $signed(_GEN_448); // @[LogMagMux.scala 136:11]
  assign _GEN_450 = 9'h1b4 == logLookUpAddr ? $signed(10'sh1c7) : $signed(_GEN_449); // @[LogMagMux.scala 136:11]
  assign _GEN_451 = 9'h1b5 == logLookUpAddr ? $signed(10'sh1c8) : $signed(_GEN_450); // @[LogMagMux.scala 136:11]
  assign _GEN_452 = 9'h1b6 == logLookUpAddr ? $signed(10'sh1c9) : $signed(_GEN_451); // @[LogMagMux.scala 136:11]
  assign _GEN_453 = 9'h1b7 == logLookUpAddr ? $signed(10'sh1c9) : $signed(_GEN_452); // @[LogMagMux.scala 136:11]
  assign _GEN_454 = 9'h1b8 == logLookUpAddr ? $signed(10'sh1ca) : $signed(_GEN_453); // @[LogMagMux.scala 136:11]
  assign _GEN_455 = 9'h1b9 == logLookUpAddr ? $signed(10'sh1cb) : $signed(_GEN_454); // @[LogMagMux.scala 136:11]
  assign _GEN_456 = 9'h1ba == logLookUpAddr ? $signed(10'sh1cc) : $signed(_GEN_455); // @[LogMagMux.scala 136:11]
  assign _GEN_457 = 9'h1bb == logLookUpAddr ? $signed(10'sh1cc) : $signed(_GEN_456); // @[LogMagMux.scala 136:11]
  assign _GEN_458 = 9'h1bc == logLookUpAddr ? $signed(10'sh1cd) : $signed(_GEN_457); // @[LogMagMux.scala 136:11]
  assign _GEN_459 = 9'h1bd == logLookUpAddr ? $signed(10'sh1ce) : $signed(_GEN_458); // @[LogMagMux.scala 136:11]
  assign _GEN_460 = 9'h1be == logLookUpAddr ? $signed(10'sh1cf) : $signed(_GEN_459); // @[LogMagMux.scala 136:11]
  assign _GEN_461 = 9'h1bf == logLookUpAddr ? $signed(10'sh1d0) : $signed(_GEN_460); // @[LogMagMux.scala 136:11]
  assign _GEN_462 = 9'h1c0 == logLookUpAddr ? $signed(10'sh1d0) : $signed(_GEN_461); // @[LogMagMux.scala 136:11]
  assign _GEN_463 = 9'h1c1 == logLookUpAddr ? $signed(10'sh1d1) : $signed(_GEN_462); // @[LogMagMux.scala 136:11]
  assign _GEN_464 = 9'h1c2 == logLookUpAddr ? $signed(10'sh1d2) : $signed(_GEN_463); // @[LogMagMux.scala 136:11]
  assign _GEN_465 = 9'h1c3 == logLookUpAddr ? $signed(10'sh1d3) : $signed(_GEN_464); // @[LogMagMux.scala 136:11]
  assign _GEN_466 = 9'h1c4 == logLookUpAddr ? $signed(10'sh1d3) : $signed(_GEN_465); // @[LogMagMux.scala 136:11]
  assign _GEN_467 = 9'h1c5 == logLookUpAddr ? $signed(10'sh1d4) : $signed(_GEN_466); // @[LogMagMux.scala 136:11]
  assign _GEN_468 = 9'h1c6 == logLookUpAddr ? $signed(10'sh1d5) : $signed(_GEN_467); // @[LogMagMux.scala 136:11]
  assign _GEN_469 = 9'h1c7 == logLookUpAddr ? $signed(10'sh1d6) : $signed(_GEN_468); // @[LogMagMux.scala 136:11]
  assign _GEN_470 = 9'h1c8 == logLookUpAddr ? $signed(10'sh1d6) : $signed(_GEN_469); // @[LogMagMux.scala 136:11]
  assign _GEN_471 = 9'h1c9 == logLookUpAddr ? $signed(10'sh1d7) : $signed(_GEN_470); // @[LogMagMux.scala 136:11]
  assign _GEN_472 = 9'h1ca == logLookUpAddr ? $signed(10'sh1d8) : $signed(_GEN_471); // @[LogMagMux.scala 136:11]
  assign _GEN_473 = 9'h1cb == logLookUpAddr ? $signed(10'sh1d9) : $signed(_GEN_472); // @[LogMagMux.scala 136:11]
  assign _GEN_474 = 9'h1cc == logLookUpAddr ? $signed(10'sh1da) : $signed(_GEN_473); // @[LogMagMux.scala 136:11]
  assign _GEN_475 = 9'h1cd == logLookUpAddr ? $signed(10'sh1da) : $signed(_GEN_474); // @[LogMagMux.scala 136:11]
  assign _GEN_476 = 9'h1ce == logLookUpAddr ? $signed(10'sh1db) : $signed(_GEN_475); // @[LogMagMux.scala 136:11]
  assign _GEN_477 = 9'h1cf == logLookUpAddr ? $signed(10'sh1dc) : $signed(_GEN_476); // @[LogMagMux.scala 136:11]
  assign _GEN_478 = 9'h1d0 == logLookUpAddr ? $signed(10'sh1dd) : $signed(_GEN_477); // @[LogMagMux.scala 136:11]
  assign _GEN_479 = 9'h1d1 == logLookUpAddr ? $signed(10'sh1dd) : $signed(_GEN_478); // @[LogMagMux.scala 136:11]
  assign _GEN_480 = 9'h1d2 == logLookUpAddr ? $signed(10'sh1de) : $signed(_GEN_479); // @[LogMagMux.scala 136:11]
  assign _GEN_481 = 9'h1d3 == logLookUpAddr ? $signed(10'sh1df) : $signed(_GEN_480); // @[LogMagMux.scala 136:11]
  assign _GEN_482 = 9'h1d4 == logLookUpAddr ? $signed(10'sh1e0) : $signed(_GEN_481); // @[LogMagMux.scala 136:11]
  assign _GEN_483 = 9'h1d5 == logLookUpAddr ? $signed(10'sh1e0) : $signed(_GEN_482); // @[LogMagMux.scala 136:11]
  assign _GEN_484 = 9'h1d6 == logLookUpAddr ? $signed(10'sh1e1) : $signed(_GEN_483); // @[LogMagMux.scala 136:11]
  assign _GEN_485 = 9'h1d7 == logLookUpAddr ? $signed(10'sh1e2) : $signed(_GEN_484); // @[LogMagMux.scala 136:11]
  assign _GEN_486 = 9'h1d8 == logLookUpAddr ? $signed(10'sh1e3) : $signed(_GEN_485); // @[LogMagMux.scala 136:11]
  assign _GEN_487 = 9'h1d9 == logLookUpAddr ? $signed(10'sh1e3) : $signed(_GEN_486); // @[LogMagMux.scala 136:11]
  assign _GEN_488 = 9'h1da == logLookUpAddr ? $signed(10'sh1e4) : $signed(_GEN_487); // @[LogMagMux.scala 136:11]
  assign _GEN_489 = 9'h1db == logLookUpAddr ? $signed(10'sh1e5) : $signed(_GEN_488); // @[LogMagMux.scala 136:11]
  assign _GEN_490 = 9'h1dc == logLookUpAddr ? $signed(10'sh1e6) : $signed(_GEN_489); // @[LogMagMux.scala 136:11]
  assign _GEN_491 = 9'h1dd == logLookUpAddr ? $signed(10'sh1e6) : $signed(_GEN_490); // @[LogMagMux.scala 136:11]
  assign _GEN_492 = 9'h1de == logLookUpAddr ? $signed(10'sh1e7) : $signed(_GEN_491); // @[LogMagMux.scala 136:11]
  assign _GEN_493 = 9'h1df == logLookUpAddr ? $signed(10'sh1e8) : $signed(_GEN_492); // @[LogMagMux.scala 136:11]
  assign _GEN_494 = 9'h1e0 == logLookUpAddr ? $signed(10'sh1e9) : $signed(_GEN_493); // @[LogMagMux.scala 136:11]
  assign _GEN_495 = 9'h1e1 == logLookUpAddr ? $signed(10'sh1e9) : $signed(_GEN_494); // @[LogMagMux.scala 136:11]
  assign _GEN_496 = 9'h1e2 == logLookUpAddr ? $signed(10'sh1ea) : $signed(_GEN_495); // @[LogMagMux.scala 136:11]
  assign _GEN_497 = 9'h1e3 == logLookUpAddr ? $signed(10'sh1eb) : $signed(_GEN_496); // @[LogMagMux.scala 136:11]
  assign _GEN_498 = 9'h1e4 == logLookUpAddr ? $signed(10'sh1ec) : $signed(_GEN_497); // @[LogMagMux.scala 136:11]
  assign _GEN_499 = 9'h1e5 == logLookUpAddr ? $signed(10'sh1ec) : $signed(_GEN_498); // @[LogMagMux.scala 136:11]
  assign _GEN_500 = 9'h1e6 == logLookUpAddr ? $signed(10'sh1ed) : $signed(_GEN_499); // @[LogMagMux.scala 136:11]
  assign _GEN_501 = 9'h1e7 == logLookUpAddr ? $signed(10'sh1ee) : $signed(_GEN_500); // @[LogMagMux.scala 136:11]
  assign _GEN_502 = 9'h1e8 == logLookUpAddr ? $signed(10'sh1ee) : $signed(_GEN_501); // @[LogMagMux.scala 136:11]
  assign _GEN_503 = 9'h1e9 == logLookUpAddr ? $signed(10'sh1ef) : $signed(_GEN_502); // @[LogMagMux.scala 136:11]
  assign _GEN_504 = 9'h1ea == logLookUpAddr ? $signed(10'sh1f0) : $signed(_GEN_503); // @[LogMagMux.scala 136:11]
  assign _GEN_505 = 9'h1eb == logLookUpAddr ? $signed(10'sh1f1) : $signed(_GEN_504); // @[LogMagMux.scala 136:11]
  assign _GEN_506 = 9'h1ec == logLookUpAddr ? $signed(10'sh1f1) : $signed(_GEN_505); // @[LogMagMux.scala 136:11]
  assign _GEN_507 = 9'h1ed == logLookUpAddr ? $signed(10'sh1f2) : $signed(_GEN_506); // @[LogMagMux.scala 136:11]
  assign _GEN_508 = 9'h1ee == logLookUpAddr ? $signed(10'sh1f3) : $signed(_GEN_507); // @[LogMagMux.scala 136:11]
  assign _GEN_509 = 9'h1ef == logLookUpAddr ? $signed(10'sh1f4) : $signed(_GEN_508); // @[LogMagMux.scala 136:11]
  assign _GEN_510 = 9'h1f0 == logLookUpAddr ? $signed(10'sh1f4) : $signed(_GEN_509); // @[LogMagMux.scala 136:11]
  assign _GEN_511 = 9'h1f1 == logLookUpAddr ? $signed(10'sh1f5) : $signed(_GEN_510); // @[LogMagMux.scala 136:11]
  assign _GEN_512 = 9'h1f2 == logLookUpAddr ? $signed(10'sh1f6) : $signed(_GEN_511); // @[LogMagMux.scala 136:11]
  assign _GEN_513 = 9'h1f3 == logLookUpAddr ? $signed(10'sh1f7) : $signed(_GEN_512); // @[LogMagMux.scala 136:11]
  assign _GEN_514 = 9'h1f4 == logLookUpAddr ? $signed(10'sh1f7) : $signed(_GEN_513); // @[LogMagMux.scala 136:11]
  assign _GEN_515 = 9'h1f5 == logLookUpAddr ? $signed(10'sh1f8) : $signed(_GEN_514); // @[LogMagMux.scala 136:11]
  assign _GEN_516 = 9'h1f6 == logLookUpAddr ? $signed(10'sh1f9) : $signed(_GEN_515); // @[LogMagMux.scala 136:11]
  assign _GEN_517 = 9'h1f7 == logLookUpAddr ? $signed(10'sh1f9) : $signed(_GEN_516); // @[LogMagMux.scala 136:11]
  assign _GEN_518 = 9'h1f8 == logLookUpAddr ? $signed(10'sh1fa) : $signed(_GEN_517); // @[LogMagMux.scala 136:11]
  assign _GEN_519 = 9'h1f9 == logLookUpAddr ? $signed(10'sh1fb) : $signed(_GEN_518); // @[LogMagMux.scala 136:11]
  assign _GEN_520 = 9'h1fa == logLookUpAddr ? $signed(10'sh1fc) : $signed(_GEN_519); // @[LogMagMux.scala 136:11]
  assign _GEN_521 = 9'h1fb == logLookUpAddr ? $signed(10'sh1fc) : $signed(_GEN_520); // @[LogMagMux.scala 136:11]
  assign _GEN_522 = 9'h1fc == logLookUpAddr ? $signed(10'sh1fd) : $signed(_GEN_521); // @[LogMagMux.scala 136:11]
  assign _GEN_523 = 9'h1fd == logLookUpAddr ? $signed(10'sh1fe) : $signed(_GEN_522); // @[LogMagMux.scala 136:11]
  assign _GEN_524 = 9'h1fe == logLookUpAddr ? $signed(10'sh1ff) : $signed(_GEN_523); // @[LogMagMux.scala 136:11]
  assign logFrac = 9'h1ff == logLookUpAddr ? $signed(10'sh1ff) : $signed(_GEN_524); // @[LogMagMux.scala 136:11]
  assign _GEN_564 = {$signed(_T_601), 9'h0}; // @[LogMagMux.scala 141:91]
  assign _GEN_565 = {{4{logFrac[9]}},logFrac}; // @[LogMagMux.scala 141:91]
  assign _T_604 = $signed(_GEN_564) + $signed(_GEN_565); // @[LogMagMux.scala 141:91]
  assign log2MagOut_imag = {{2{_T_604[13]}},_T_604}; // @[LogMagMux.scala 160:38]
  assign _T_630 = 2'h3 == _T_617; // @[Mux.scala 68:19]
  assign _T_633_real = _T_630 ? $signed(16'sh0) : $signed(io_in_bits_real); // @[Mux.scala 68:16]
  assign _T_633_imag = _T_630 ? $signed(log2MagOut_imag) : $signed(io_in_bits_imag); // @[Mux.scala 68:16]
  assign _T_634 = 2'h2 == _T_617; // @[Mux.scala 68:19]
  assign _T_637_real = _T_634 ? $signed(16'sh0) : $signed(_T_633_real); // @[Mux.scala 68:16]
  assign jplMagOut_imag = jplMag[15:0]; // @[LogMagMux.scala 151:23 LogMagMux.scala 154:18]
  assign _T_637_imag = _T_634 ? $signed(jplMagOut_imag) : $signed(_T_633_imag); // @[Mux.scala 68:16]
  assign _T_638 = 2'h1 == _T_617; // @[Mux.scala 68:19]
  assign _T_641_real = _T_638 ? $signed(16'sh0) : $signed(_T_637_real); // @[Mux.scala 68:16]
  assign _GEN_567 = _T_31[33:1]; // @[LogMagMux.scala 95:20 LogMagMux.scala 105:10]
  assign magSqr = _GEN_567[15:0]; // @[LogMagMux.scala 95:20 LogMagMux.scala 105:10]
  assign _T_641_imag = _T_638 ? $signed(magSqr) : $signed(_T_637_imag); // @[Mux.scala 68:16]
  assign _T_642 = 2'h0 == _T_617; // @[Mux.scala 68:19]
  assign output_mux_real = _T_642 ? $signed(_T_629_real) : $signed(_T_641_real); // @[Mux.scala 68:16]
  assign output_mux_imag = _T_642 ? $signed(_T_629_imag) : $signed(_T_641_imag); // @[Mux.scala 68:16]
  assign _T_645 = io_in_ready & io_in_valid; // @[Decoupled.scala 40:37]
  assign _T_656 = _T_653 + 3'h1; // @[LogMagMux.scala 193:22]
  assign _T_657 = _T_653 == 3'h3; // @[LogMagMux.scala 196:18]
  assign _T_659 = _T_657 & _T_645; // @[LogMagMux.scala 196:39]
  assign _GEN_544 = _T_659 | initialInDone; // @[LogMagMux.scala 196:56]
  assign _T_667 = ~initialInDone; // @[Skid.scala 29:30]
  assign _T_668 = io_out_ready | _T_667; // @[Skid.scala 29:27]
  assign skidInData_ready = _T_668; // @[LogMagMux.scala 205:24 Skid.scala 29:14]
  assign skidInData_valid = io_in_valid; // @[LogMagMux.scala 205:24 LogMagMux.scala 207:20]
  assign _T_662 = skidInData_ready & skidInData_valid; // @[Decoupled.scala 40:37]
  assign _T_677 = _T_668 & io_in_valid; // @[Decoupled.scala 40:37]
  assign skidInData_bits_real = output_mux_real; // @[LogMagMux.scala 205:24 LogMagMux.scala 206:19]
  assign skidInData_bits_imag = output_mux_imag; // @[LogMagMux.scala 205:24 LogMagMux.scala 206:19]
  assign io_in_ready = skidInData_ready; // @[LogMagMux.scala 210:15]
  assign io_out_valid = Queue_io_deq_valid; // @[Skid.scala 31:15]
  assign io_out_bits_real = Queue_io_deq_bits_real; // @[Skid.scala 32:14]
  assign io_out_bits_imag = Queue_io_deq_bits_imag; // @[Skid.scala 32:14]
  assign io_lastOut = Queue_1_io_deq_bits; // @[LogMagMux.scala 220:20]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = _T_666; // @[Skid.scala 25:24]
  assign Queue_io_enq_bits_real = output_mux_real; // @[LogMagMux.scala 211:52]
  assign Queue_io_enq_bits_imag = output_mux_imag; // @[LogMagMux.scala 211:52]
  assign Queue_io_deq_ready = io_out_ready; // @[Skid.scala 30:24]
  assign Queue_1_clock = clock;
  assign Queue_1_reset = reset;
  assign Queue_1_io_enq_valid = _T_681; // @[Skid.scala 25:24]
  assign Queue_1_io_enq_bits = _T_676; // @[LogMagMux.scala 219:59]
  assign Queue_1_io_deq_ready = io_out_ready; // @[Skid.scala 30:24]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_16 = _RAND_0[16:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  jplMagOp1 = _RAND_1[16:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  tmpOp2 = _RAND_2[16:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_20 = _RAND_3[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  jplMagOp2 = _RAND_4[17:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_23 = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_26 = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {2{`RANDOM}};
  _T_29 = _RAND_7[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {2{`RANDOM}};
  _T_30 = _RAND_8[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {2{`RANDOM}};
  _T_31 = _RAND_9[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_33 = _RAND_10[17:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  jplMag = _RAND_11[17:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  noLeadOne = _RAND_12[17:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  shiftNum = _RAND_13[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_601 = _RAND_14[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_614 = _RAND_15[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_615 = _RAND_16[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_616 = _RAND_17[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_617 = _RAND_18[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_620_real = _RAND_19[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_620_imag = _RAND_20[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_623_real = _RAND_21[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_623_imag = _RAND_22[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_626_real = _RAND_23[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_626_imag = _RAND_24[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_629_real = _RAND_25[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_629_imag = _RAND_26[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  initialInDone = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_653 = _RAND_28[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_663 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_664 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T_665 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _T_666 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _T_673 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _T_674 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _T_675 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _T_676 = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _T_678 = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _T_679 = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _T_680 = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _T_681 = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_16 <= $signed(u) + $signed(_GEN_559);
    jplMagOp1 <= _T_16;
    tmpOp2 <= $signed(u) - $signed(_GEN_560);
    _T_20 <= v[15:1];
    jplMagOp2 <= $signed(tmpOp2) + $signed(_GEN_561);
    _T_23 <= $signed(absInReal) * $signed(absInReal);
    _T_26 <= $signed(absInImag) * $signed(absInImag);
    _T_29 <= $signed(_T_24) + $signed(_T_27);
    _T_30 <= _T_29;
    _T_31 <= _T_30;
    if (_T_32) begin
      _T_33 <= {{1{jplMagOp1[16]}},jplMagOp1};
    end else begin
      _T_33 <= jplMagOp2;
    end
    jplMag <= _T_33;
    noLeadOne <= _T_589 - _T_590[17:0];
    shiftNum <= _T_596 - 5'h1;
    _T_601 <= logUInt - 5'h0;
    _T_614 <= io_sel;
    _T_615 <= _T_614;
    _T_616 <= _T_615;
    _T_617 <= _T_616;
    _T_620_real <= io_in_bits_real;
    _T_620_imag <= io_in_bits_imag;
    _T_623_real <= _T_620_real;
    _T_623_imag <= _T_620_imag;
    _T_626_real <= _T_623_real;
    _T_626_imag <= _T_623_imag;
    _T_629_real <= _T_626_real;
    _T_629_imag <= _T_626_imag;
    if (reset) begin
      initialInDone <= 1'h0;
    end else if (io_lastOut) begin
      initialInDone <= 1'h0;
    end else begin
      initialInDone <= _GEN_544;
    end
    if (reset) begin
      _T_653 <= 3'h0;
    end else if (io_lastOut) begin
      _T_653 <= 3'h0;
    end else if (_T_645) begin
      _T_653 <= _T_656;
    end
    if (reset) begin
      _T_663 <= 1'h0;
    end else begin
      _T_663 <= _T_662;
    end
    if (reset) begin
      _T_664 <= 1'h0;
    end else begin
      _T_664 <= _T_663;
    end
    if (reset) begin
      _T_665 <= 1'h0;
    end else begin
      _T_665 <= _T_664;
    end
    if (reset) begin
      _T_666 <= 1'h0;
    end else begin
      _T_666 <= _T_665;
    end
    _T_673 <= io_lastIn & _T_645;
    _T_674 <= _T_673;
    _T_675 <= _T_674;
    _T_676 <= _T_675;
    if (reset) begin
      _T_678 <= 1'h0;
    end else begin
      _T_678 <= _T_677;
    end
    if (reset) begin
      _T_679 <= 1'h0;
    end else begin
      _T_679 <= _T_678;
    end
    if (reset) begin
      _T_680 <= 1'h0;
    end else begin
      _T_680 <= _T_679;
    end
    if (reset) begin
      _T_681 <= 1'h0;
    end else begin
      _T_681 <= _T_680;
    end
  end
endmodule
module AXI4LogMagMuxBlock(
  input         clock,
  input         reset,
  output        auto_mem_in_aw_ready,
  input         auto_mem_in_aw_valid,
  input         auto_mem_in_aw_bits_id,
  input  [29:0] auto_mem_in_aw_bits_addr,
  output        auto_mem_in_w_ready,
  input         auto_mem_in_w_valid,
  input  [31:0] auto_mem_in_w_bits_data,
  input  [3:0]  auto_mem_in_w_bits_strb,
  input         auto_mem_in_b_ready,
  output        auto_mem_in_b_valid,
  output        auto_mem_in_b_bits_id,
  output        auto_mem_in_ar_ready,
  input         auto_mem_in_ar_valid,
  input         auto_mem_in_ar_bits_id,
  input  [29:0] auto_mem_in_ar_bits_addr,
  input  [2:0]  auto_mem_in_ar_bits_size,
  input         auto_mem_in_r_ready,
  output        auto_mem_in_r_valid,
  output        auto_mem_in_r_bits_id,
  output [31:0] auto_mem_in_r_bits_data,
  output        auto_stream_in_ready,
  input         auto_stream_in_valid,
  input  [31:0] auto_stream_in_bits_data,
  input         auto_stream_in_bits_last,
  input         auto_stream_out_ready,
  output        auto_stream_out_valid,
  output [31:0] auto_stream_out_bits_data,
  output        auto_stream_out_bits_last
);
  wire  logMagMux_clock; // @[LogMagMuxDspBlock.scala 27:27]
  wire  logMagMux_reset; // @[LogMagMuxDspBlock.scala 27:27]
  wire  logMagMux_io_in_ready; // @[LogMagMuxDspBlock.scala 27:27]
  wire  logMagMux_io_in_valid; // @[LogMagMuxDspBlock.scala 27:27]
  wire [15:0] logMagMux_io_in_bits_real; // @[LogMagMuxDspBlock.scala 27:27]
  wire [15:0] logMagMux_io_in_bits_imag; // @[LogMagMuxDspBlock.scala 27:27]
  wire  logMagMux_io_lastIn; // @[LogMagMuxDspBlock.scala 27:27]
  wire  logMagMux_io_out_ready; // @[LogMagMuxDspBlock.scala 27:27]
  wire  logMagMux_io_out_valid; // @[LogMagMuxDspBlock.scala 27:27]
  wire [15:0] logMagMux_io_out_bits_real; // @[LogMagMuxDspBlock.scala 27:27]
  wire [15:0] logMagMux_io_out_bits_imag; // @[LogMagMuxDspBlock.scala 27:27]
  wire [1:0] logMagMux_io_sel; // @[LogMagMuxDspBlock.scala 27:27]
  wire  logMagMux_io_lastOut; // @[LogMagMuxDspBlock.scala 27:27]
  wire  Queue_clock; // @[Decoupled.scala 287:21]
  wire  Queue_reset; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_read; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_enq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_extra; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_read; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_deq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_extra; // @[Decoupled.scala 287:21]
  reg [1:0] selReg; // @[LogMagMuxDspBlock.scala 29:33]
  reg [31:0] _RAND_0;
  wire  _T_2; // @[RegisterRouter.scala 40:39]
  wire  _T_3; // @[RegisterRouter.scala 40:26]
  wire  _T_4; // @[RegisterRouter.scala 42:29]
  wire  _T_47_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 290:17]
  wire [29:0] _T_11; // @[RegisterRouter.scala 48:19]
  wire  _T_53; // @[RegisterRouter.scala 59:16]
  wire  _T_5; // @[RegisterRouter.scala 42:26]
  wire [1:0] _T_14; // @[OneHot.scala 65:12]
  wire [1:0] _T_16; // @[Misc.scala 200:81]
  wire  _T_17; // @[Misc.scala 204:21]
  wire  _T_20; // @[Misc.scala 209:20]
  wire  _T_22; // @[Misc.scala 213:38]
  wire  _T_23; // @[Misc.scala 213:29]
  wire  _T_25; // @[Misc.scala 213:38]
  wire  _T_26; // @[Misc.scala 213:29]
  wire  _T_29; // @[Misc.scala 209:20]
  wire  _T_30; // @[Misc.scala 212:27]
  wire  _T_31; // @[Misc.scala 213:38]
  wire  _T_32; // @[Misc.scala 213:29]
  wire  _T_33; // @[Misc.scala 212:27]
  wire  _T_34; // @[Misc.scala 213:38]
  wire  _T_35; // @[Misc.scala 213:29]
  wire  _T_36; // @[Misc.scala 212:27]
  wire  _T_37; // @[Misc.scala 213:38]
  wire  _T_38; // @[Misc.scala 213:29]
  wire  _T_39; // @[Misc.scala 212:27]
  wire  _T_40; // @[Misc.scala 213:38]
  wire  _T_41; // @[Misc.scala 213:29]
  wire [3:0] _T_44; // @[Cat.scala 29:58]
  wire [3:0] _T_46; // @[RegisterRouter.scala 54:25]
  wire [7:0] _T_63; // @[Bitwise.scala 72:12]
  wire [7:0] _T_65; // @[Bitwise.scala 72:12]
  wire [7:0] _T_67; // @[Bitwise.scala 72:12]
  wire [7:0] _T_69; // @[Bitwise.scala 72:12]
  wire [31:0] _T_72; // @[Cat.scala 29:58]
  wire  _T_91; // @[RegisterRouter.scala 59:16]
  wire  _T_117; // @[RegisterRouter.scala 59:16]
  wire  _T_129; // @[RegisterRouter.scala 59:16]
  wire  _T_132; // @[RegisterRouter.scala 59:16]
  wire  _T_98; // @[RegisterRouter.scala 59:16]
  wire [1:0] _T_171; // @[RegisterRouter.scala 59:16]
  wire  _T_172_bits_read; // @[Decoupled.scala 308:19 Decoupled.scala 309:14]
  wire  _T_172_valid; // @[Decoupled.scala 308:19 Decoupled.scala 310:15]
  wire  _T_175; // @[RegisterRouter.scala 65:29]
  LogMagMux logMagMux ( // @[LogMagMuxDspBlock.scala 27:27]
    .clock(logMagMux_clock),
    .reset(logMagMux_reset),
    .io_in_ready(logMagMux_io_in_ready),
    .io_in_valid(logMagMux_io_in_valid),
    .io_in_bits_real(logMagMux_io_in_bits_real),
    .io_in_bits_imag(logMagMux_io_in_bits_imag),
    .io_lastIn(logMagMux_io_lastIn),
    .io_out_ready(logMagMux_io_out_ready),
    .io_out_valid(logMagMux_io_out_valid),
    .io_out_bits_real(logMagMux_io_out_bits_real),
    .io_out_bits_imag(logMagMux_io_out_bits_imag),
    .io_sel(logMagMux_io_sel),
    .io_lastOut(logMagMux_io_lastOut)
  );
  Queue Queue ( // @[Decoupled.scala 287:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_read(Queue_io_enq_bits_read),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_extra(Queue_io_enq_bits_extra),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_read(Queue_io_deq_bits_read),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_extra(Queue_io_deq_bits_extra)
  );
  assign _T_2 = auto_mem_in_aw_valid & auto_mem_in_w_valid; // @[RegisterRouter.scala 40:39]
  assign _T_3 = auto_mem_in_ar_valid | _T_2; // @[RegisterRouter.scala 40:26]
  assign _T_4 = ~auto_mem_in_ar_valid; // @[RegisterRouter.scala 42:29]
  assign _T_47_ready = Queue_io_enq_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 290:17]
  assign _T_11 = auto_mem_in_ar_valid ? auto_mem_in_ar_bits_addr : auto_mem_in_aw_bits_addr; // @[RegisterRouter.scala 48:19]
  assign _T_53 = _T_11[7:2] == 6'h0; // @[RegisterRouter.scala 59:16]
  assign _T_5 = _T_47_ready & _T_4; // @[RegisterRouter.scala 42:26]
  assign _T_14 = 2'h1 << auto_mem_in_ar_bits_size[0]; // @[OneHot.scala 65:12]
  assign _T_16 = _T_14 | 2'h1; // @[Misc.scala 200:81]
  assign _T_17 = auto_mem_in_ar_bits_size >= 3'h2; // @[Misc.scala 204:21]
  assign _T_20 = ~auto_mem_in_ar_bits_addr[1]; // @[Misc.scala 209:20]
  assign _T_22 = _T_16[1] & _T_20; // @[Misc.scala 213:38]
  assign _T_23 = _T_17 | _T_22; // @[Misc.scala 213:29]
  assign _T_25 = _T_16[1] & auto_mem_in_ar_bits_addr[1]; // @[Misc.scala 213:38]
  assign _T_26 = _T_17 | _T_25; // @[Misc.scala 213:29]
  assign _T_29 = ~auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 209:20]
  assign _T_30 = _T_20 & _T_29; // @[Misc.scala 212:27]
  assign _T_31 = _T_16[0] & _T_30; // @[Misc.scala 213:38]
  assign _T_32 = _T_23 | _T_31; // @[Misc.scala 213:29]
  assign _T_33 = _T_20 & auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  assign _T_34 = _T_16[0] & _T_33; // @[Misc.scala 213:38]
  assign _T_35 = _T_23 | _T_34; // @[Misc.scala 213:29]
  assign _T_36 = auto_mem_in_ar_bits_addr[1] & _T_29; // @[Misc.scala 212:27]
  assign _T_37 = _T_16[0] & _T_36; // @[Misc.scala 213:38]
  assign _T_38 = _T_26 | _T_37; // @[Misc.scala 213:29]
  assign _T_39 = auto_mem_in_ar_bits_addr[1] & auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  assign _T_40 = _T_16[0] & _T_39; // @[Misc.scala 213:38]
  assign _T_41 = _T_26 | _T_40; // @[Misc.scala 213:29]
  assign _T_44 = {_T_41,_T_38,_T_35,_T_32}; // @[Cat.scala 29:58]
  assign _T_46 = auto_mem_in_ar_valid ? _T_44 : auto_mem_in_w_bits_strb; // @[RegisterRouter.scala 54:25]
  assign _T_63 = _T_46[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_65 = _T_46[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_67 = _T_46[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_69 = _T_46[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_72 = {_T_69,_T_67,_T_65,_T_63}; // @[Cat.scala 29:58]
  assign _T_91 = _T_72[1:0] == 2'h3; // @[RegisterRouter.scala 59:16]
  assign _T_117 = _T_3 & _T_47_ready; // @[RegisterRouter.scala 59:16]
  assign _T_129 = _T_117 & _T_4; // @[RegisterRouter.scala 59:16]
  assign _T_132 = _T_129 & _T_53; // @[RegisterRouter.scala 59:16]
  assign _T_98 = _T_132 & _T_91; // @[RegisterRouter.scala 59:16]
  assign _T_171 = _T_53 ? selReg : 2'h0; // @[RegisterRouter.scala 59:16]
  assign _T_172_bits_read = Queue_io_deq_bits_read; // @[Decoupled.scala 308:19 Decoupled.scala 309:14]
  assign _T_172_valid = Queue_io_deq_valid; // @[Decoupled.scala 308:19 Decoupled.scala 310:15]
  assign _T_175 = ~_T_172_bits_read; // @[RegisterRouter.scala 65:29]
  assign auto_mem_in_aw_ready = _T_5 & auto_mem_in_w_valid; // @[LazyModule.scala 173:31]
  assign auto_mem_in_w_ready = _T_5 & auto_mem_in_aw_valid; // @[LazyModule.scala 173:31]
  assign auto_mem_in_b_valid = _T_172_valid & _T_175; // @[LazyModule.scala 173:31]
  assign auto_mem_in_b_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_mem_in_ar_ready = Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_valid = _T_172_valid & _T_172_bits_read; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 173:31]
  assign auto_stream_in_ready = logMagMux_io_in_ready; // @[LazyModule.scala 173:31]
  assign auto_stream_out_valid = logMagMux_io_out_valid; // @[LazyModule.scala 173:49]
  assign auto_stream_out_bits_data = {logMagMux_io_out_bits_real,logMagMux_io_out_bits_imag}; // @[LazyModule.scala 173:49]
  assign auto_stream_out_bits_last = logMagMux_io_lastOut; // @[LazyModule.scala 173:49]
  assign logMagMux_clock = clock;
  assign logMagMux_reset = reset;
  assign logMagMux_io_in_valid = auto_stream_in_valid; // @[LogMagMuxDspBlock.scala 40:30]
  assign logMagMux_io_in_bits_real = auto_stream_in_bits_data[31:16]; // @[LogMagMuxDspBlock.scala 41:30]
  assign logMagMux_io_in_bits_imag = auto_stream_in_bits_data[15:0]; // @[LogMagMuxDspBlock.scala 41:30]
  assign logMagMux_io_lastIn = auto_stream_in_bits_last; // @[LogMagMuxDspBlock.scala 44:31]
  assign logMagMux_io_out_ready = auto_stream_out_ready; // @[LogMagMuxDspBlock.scala 49:28]
  assign logMagMux_io_sel = selReg; // @[LogMagMuxDspBlock.scala 35:22]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_mem_in_ar_valid | _T_2; // @[Decoupled.scala 288:22]
  assign Queue_io_enq_bits_read = auto_mem_in_ar_valid; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_data = {{30'd0}, _T_171}; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_extra = auto_mem_in_ar_valid ? auto_mem_in_ar_bits_id : auto_mem_in_aw_bits_id; // @[Decoupled.scala 289:21]
  assign Queue_io_deq_ready = _T_172_bits_read ? auto_mem_in_r_ready : auto_mem_in_b_ready; // @[Decoupled.scala 311:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  selReg = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      selReg <= 2'h0;
    end else if (_T_98) begin
      selReg <= auto_mem_in_w_bits_data[1:0];
    end
  end
endmodule
module AXI4Splitter_4(
  input         clock,
  input         reset,
  output        auto_mem_in_aw_ready,
  input         auto_mem_in_aw_valid,
  input         auto_mem_in_aw_bits_id,
  input  [29:0] auto_mem_in_aw_bits_addr,
  output        auto_mem_in_w_ready,
  input         auto_mem_in_w_valid,
  input  [31:0] auto_mem_in_w_bits_data,
  input  [3:0]  auto_mem_in_w_bits_strb,
  input         auto_mem_in_b_ready,
  output        auto_mem_in_b_valid,
  output        auto_mem_in_b_bits_id,
  output        auto_mem_in_ar_ready,
  input         auto_mem_in_ar_valid,
  input         auto_mem_in_ar_bits_id,
  input  [29:0] auto_mem_in_ar_bits_addr,
  input  [2:0]  auto_mem_in_ar_bits_size,
  input         auto_mem_in_r_ready,
  output        auto_mem_in_r_valid,
  output        auto_mem_in_r_bits_id,
  output [31:0] auto_mem_in_r_bits_data,
  output        auto_stream_in_ready,
  input         auto_stream_in_valid,
  input  [31:0] auto_stream_in_bits_data,
  input         auto_stream_in_bits_last,
  input         auto_stream_out_1_ready,
  output        auto_stream_out_1_valid,
  output [31:0] auto_stream_out_1_bits_data,
  output        auto_stream_out_1_bits_last,
  input         auto_stream_out_0_ready,
  output        auto_stream_out_0_valid,
  output [31:0] auto_stream_out_0_bits_data,
  output        auto_stream_out_0_bits_last
);
  wire  Queue_clock; // @[Decoupled.scala 287:21]
  wire  Queue_reset; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_read; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_enq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_extra; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_read; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_deq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_extra; // @[Decoupled.scala 287:21]
  reg [31:0] ctrlReg; // @[Splitter.scala 27:26]
  reg [31:0] _RAND_0;
  reg [31:0] maskReg; // @[Splitter.scala 28:26]
  reg [31:0] _RAND_1;
  wire  _T_4; // @[RegisterRouter.scala 40:39]
  wire  _T_5; // @[RegisterRouter.scala 40:26]
  wire  _T_6; // @[RegisterRouter.scala 42:29]
  wire  _T_49_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 290:17]
  wire [29:0] _T_13; // @[RegisterRouter.scala 48:19]
  wire [1:0] _T_53; // @[RegisterRouter.scala 59:16]
  wire  _T_55; // @[RegisterRouter.scala 59:16]
  wire  _T_7; // @[RegisterRouter.scala 42:26]
  wire [1:0] _T_16; // @[OneHot.scala 65:12]
  wire [1:0] _T_18; // @[Misc.scala 200:81]
  wire  _T_19; // @[Misc.scala 204:21]
  wire  _T_22; // @[Misc.scala 209:20]
  wire  _T_24; // @[Misc.scala 213:38]
  wire  _T_25; // @[Misc.scala 213:29]
  wire  _T_27; // @[Misc.scala 213:38]
  wire  _T_28; // @[Misc.scala 213:29]
  wire  _T_31; // @[Misc.scala 209:20]
  wire  _T_32; // @[Misc.scala 212:27]
  wire  _T_33; // @[Misc.scala 213:38]
  wire  _T_34; // @[Misc.scala 213:29]
  wire  _T_35; // @[Misc.scala 212:27]
  wire  _T_36; // @[Misc.scala 213:38]
  wire  _T_37; // @[Misc.scala 213:29]
  wire  _T_38; // @[Misc.scala 212:27]
  wire  _T_39; // @[Misc.scala 213:38]
  wire  _T_40; // @[Misc.scala 213:29]
  wire  _T_41; // @[Misc.scala 212:27]
  wire  _T_42; // @[Misc.scala 213:38]
  wire  _T_43; // @[Misc.scala 213:29]
  wire [3:0] _T_46; // @[Cat.scala 29:58]
  wire [3:0] _T_48; // @[RegisterRouter.scala 54:25]
  wire [7:0] _T_67; // @[Bitwise.scala 72:12]
  wire [7:0] _T_69; // @[Bitwise.scala 72:12]
  wire [7:0] _T_71; // @[Bitwise.scala 72:12]
  wire [7:0] _T_73; // @[Bitwise.scala 72:12]
  wire [31:0] _T_76; // @[Cat.scala 29:58]
  wire  _T_95; // @[RegisterRouter.scala 59:16]
  wire  _T_148; // @[RegisterRouter.scala 59:16]
  wire [1:0] _T_142; // @[OneHot.scala 58:35]
  wire  _T_165; // @[RegisterRouter.scala 59:16]
  wire  _T_172; // @[RegisterRouter.scala 59:16]
  wire  _T_173; // @[RegisterRouter.scala 59:16]
  wire  _T_102; // @[RegisterRouter.scala 59:16]
  wire  _T_167; // @[RegisterRouter.scala 59:16]
  wire  _T_168; // @[RegisterRouter.scala 59:16]
  wire  _T_125; // @[RegisterRouter.scala 59:16]
  wire  _GEN_11; // @[MuxLiteral.scala 48:10]
  wire [31:0] _GEN_13; // @[MuxLiteral.scala 48:10]
  wire  _T_223_bits_read; // @[Decoupled.scala 308:19 Decoupled.scala 309:14]
  wire  _T_223_valid; // @[Decoupled.scala 308:19 Decoupled.scala 310:15]
  wire  _T_226; // @[RegisterRouter.scala 65:29]
  wire  readyOR; // @[Splitter.scala 45:34]
  wire  readyAND; // @[Splitter.scala 46:34]
  wire  _T_229; // @[Splitter.scala 49:19]
  wire  _T_230; // @[Splitter.scala 52:24]
  wire  _GEN_14; // @[Splitter.scala 52:33]
  wire  _T_233; // @[Splitter.scala 62:34]
  wire  _T_237; // @[Splitter.scala 62:34]
  Queue Queue ( // @[Decoupled.scala 287:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_read(Queue_io_enq_bits_read),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_extra(Queue_io_enq_bits_extra),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_read(Queue_io_deq_bits_read),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_extra(Queue_io_deq_bits_extra)
  );
  assign _T_4 = auto_mem_in_aw_valid & auto_mem_in_w_valid; // @[RegisterRouter.scala 40:39]
  assign _T_5 = auto_mem_in_ar_valid | _T_4; // @[RegisterRouter.scala 40:26]
  assign _T_6 = ~auto_mem_in_ar_valid; // @[RegisterRouter.scala 42:29]
  assign _T_49_ready = Queue_io_enq_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 290:17]
  assign _T_13 = auto_mem_in_ar_valid ? auto_mem_in_ar_bits_addr : auto_mem_in_aw_bits_addr; // @[RegisterRouter.scala 48:19]
  assign _T_53 = _T_13[3:2] & 2'h2; // @[RegisterRouter.scala 59:16]
  assign _T_55 = _T_53 == 2'h0; // @[RegisterRouter.scala 59:16]
  assign _T_7 = _T_49_ready & _T_6; // @[RegisterRouter.scala 42:26]
  assign _T_16 = 2'h1 << auto_mem_in_ar_bits_size[0]; // @[OneHot.scala 65:12]
  assign _T_18 = _T_16 | 2'h1; // @[Misc.scala 200:81]
  assign _T_19 = auto_mem_in_ar_bits_size >= 3'h2; // @[Misc.scala 204:21]
  assign _T_22 = ~auto_mem_in_ar_bits_addr[1]; // @[Misc.scala 209:20]
  assign _T_24 = _T_18[1] & _T_22; // @[Misc.scala 213:38]
  assign _T_25 = _T_19 | _T_24; // @[Misc.scala 213:29]
  assign _T_27 = _T_18[1] & auto_mem_in_ar_bits_addr[1]; // @[Misc.scala 213:38]
  assign _T_28 = _T_19 | _T_27; // @[Misc.scala 213:29]
  assign _T_31 = ~auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 209:20]
  assign _T_32 = _T_22 & _T_31; // @[Misc.scala 212:27]
  assign _T_33 = _T_18[0] & _T_32; // @[Misc.scala 213:38]
  assign _T_34 = _T_25 | _T_33; // @[Misc.scala 213:29]
  assign _T_35 = _T_22 & auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  assign _T_36 = _T_18[0] & _T_35; // @[Misc.scala 213:38]
  assign _T_37 = _T_25 | _T_36; // @[Misc.scala 213:29]
  assign _T_38 = auto_mem_in_ar_bits_addr[1] & _T_31; // @[Misc.scala 212:27]
  assign _T_39 = _T_18[0] & _T_38; // @[Misc.scala 213:38]
  assign _T_40 = _T_28 | _T_39; // @[Misc.scala 213:29]
  assign _T_41 = auto_mem_in_ar_bits_addr[1] & auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  assign _T_42 = _T_18[0] & _T_41; // @[Misc.scala 213:38]
  assign _T_43 = _T_28 | _T_42; // @[Misc.scala 213:29]
  assign _T_46 = {_T_43,_T_40,_T_37,_T_34}; // @[Cat.scala 29:58]
  assign _T_48 = auto_mem_in_ar_valid ? _T_46 : auto_mem_in_w_bits_strb; // @[RegisterRouter.scala 54:25]
  assign _T_67 = _T_48[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_69 = _T_48[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_71 = _T_48[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_73 = _T_48[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_76 = {_T_73,_T_71,_T_69,_T_67}; // @[Cat.scala 29:58]
  assign _T_95 = _T_76 == 32'hffffffff; // @[RegisterRouter.scala 59:16]
  assign _T_148 = _T_5 & _T_49_ready; // @[RegisterRouter.scala 59:16]
  assign _T_142 = 2'h1 << _T_13[2]; // @[OneHot.scala 58:35]
  assign _T_165 = _T_148 & _T_6; // @[RegisterRouter.scala 59:16]
  assign _T_172 = _T_165 & _T_142[1]; // @[RegisterRouter.scala 59:16]
  assign _T_173 = _T_172 & _T_55; // @[RegisterRouter.scala 59:16]
  assign _T_102 = _T_173 & _T_95; // @[RegisterRouter.scala 59:16]
  assign _T_167 = _T_165 & _T_142[0]; // @[RegisterRouter.scala 59:16]
  assign _T_168 = _T_167 & _T_55; // @[RegisterRouter.scala 59:16]
  assign _T_125 = _T_168 & _T_95; // @[RegisterRouter.scala 59:16]
  assign _GEN_11 = _T_13[2] ? _T_55 : _T_55; // @[MuxLiteral.scala 48:10]
  assign _GEN_13 = _T_13[2] ? maskReg : ctrlReg; // @[MuxLiteral.scala 48:10]
  assign _T_223_bits_read = Queue_io_deq_bits_read; // @[Decoupled.scala 308:19 Decoupled.scala 309:14]
  assign _T_223_valid = Queue_io_deq_valid; // @[Decoupled.scala 308:19 Decoupled.scala 310:15]
  assign _T_226 = ~_T_223_bits_read; // @[RegisterRouter.scala 65:29]
  assign readyOR = auto_stream_out_0_ready | auto_stream_out_1_ready; // @[Splitter.scala 45:34]
  assign readyAND = auto_stream_out_0_ready & auto_stream_out_1_ready; // @[Splitter.scala 46:34]
  assign _T_229 = ctrlReg == 32'h0; // @[Splitter.scala 49:19]
  assign _T_230 = ctrlReg == 32'h1; // @[Splitter.scala 52:24]
  assign _GEN_14 = _T_230 & readyOR; // @[Splitter.scala 52:33]
  assign _T_233 = ~maskReg[0]; // @[Splitter.scala 62:34]
  assign _T_237 = ~maskReg[1]; // @[Splitter.scala 62:34]
  assign auto_mem_in_aw_ready = _T_7 & auto_mem_in_w_valid; // @[LazyModule.scala 173:31]
  assign auto_mem_in_w_ready = _T_7 & auto_mem_in_aw_valid; // @[LazyModule.scala 173:31]
  assign auto_mem_in_b_valid = _T_223_valid & _T_226; // @[LazyModule.scala 173:31]
  assign auto_mem_in_b_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_mem_in_ar_ready = Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_valid = _T_223_valid & _T_223_bits_read; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 173:31]
  assign auto_stream_in_ready = _T_229 ? readyAND : _GEN_14; // @[LazyModule.scala 173:31]
  assign auto_stream_out_1_valid = auto_stream_in_valid & _T_237; // @[LazyModule.scala 173:49]
  assign auto_stream_out_1_bits_data = auto_stream_in_bits_data; // @[LazyModule.scala 173:49]
  assign auto_stream_out_1_bits_last = auto_stream_in_bits_last; // @[LazyModule.scala 173:49]
  assign auto_stream_out_0_valid = auto_stream_in_valid & _T_233; // @[LazyModule.scala 173:49]
  assign auto_stream_out_0_bits_data = auto_stream_in_bits_data; // @[LazyModule.scala 173:49]
  assign auto_stream_out_0_bits_last = auto_stream_in_bits_last; // @[LazyModule.scala 173:49]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_mem_in_ar_valid | _T_4; // @[Decoupled.scala 288:22]
  assign Queue_io_enq_bits_read = auto_mem_in_ar_valid; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_data = _GEN_11 ? _GEN_13 : 32'h0; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_extra = auto_mem_in_ar_valid ? auto_mem_in_ar_bits_id : auto_mem_in_aw_bits_id; // @[Decoupled.scala 289:21]
  assign Queue_io_deq_ready = _T_223_bits_read ? auto_mem_in_r_ready : auto_mem_in_b_ready; // @[Decoupled.scala 311:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ctrlReg = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  maskReg = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      ctrlReg <= 32'h0;
    end else if (_T_125) begin
      ctrlReg <= auto_mem_in_w_bits_data;
    end
    if (reset) begin
      maskReg <= 32'h0;
    end else if (_T_102) begin
      maskReg <= auto_mem_in_w_bits_data;
    end
  end
endmodule
module AXI4StreamMux_6(
  input         clock,
  input         reset,
  output        auto_register_in_aw_ready,
  input         auto_register_in_aw_valid,
  input         auto_register_in_aw_bits_id,
  input  [29:0] auto_register_in_aw_bits_addr,
  output        auto_register_in_w_ready,
  input         auto_register_in_w_valid,
  input  [31:0] auto_register_in_w_bits_data,
  input  [3:0]  auto_register_in_w_bits_strb,
  input         auto_register_in_b_ready,
  output        auto_register_in_b_valid,
  output        auto_register_in_b_bits_id,
  output        auto_register_in_ar_ready,
  input         auto_register_in_ar_valid,
  input         auto_register_in_ar_bits_id,
  input  [29:0] auto_register_in_ar_bits_addr,
  input  [2:0]  auto_register_in_ar_bits_size,
  input         auto_register_in_r_ready,
  output        auto_register_in_r_valid,
  output        auto_register_in_r_bits_id,
  output [31:0] auto_register_in_r_bits_data,
  output        auto_stream_in_2_ready,
  input         auto_stream_in_2_valid,
  input  [31:0] auto_stream_in_2_bits_data,
  input         auto_stream_in_2_bits_last,
  output        auto_stream_in_1_ready,
  input         auto_stream_in_1_valid,
  input  [31:0] auto_stream_in_1_bits_data,
  input         auto_stream_in_1_bits_last,
  output        auto_stream_in_0_ready,
  input         auto_stream_in_0_valid,
  input  [31:0] auto_stream_in_0_bits_data,
  input         auto_stream_in_0_bits_last,
  input         auto_stream_out_0_ready,
  output        auto_stream_out_0_valid,
  output [31:0] auto_stream_out_0_bits_data,
  output        auto_stream_out_0_bits_last
);
  wire  Queue_clock; // @[Decoupled.scala 287:21]
  wire  Queue_reset; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_read; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_enq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_extra; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_read; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_deq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_extra; // @[Decoupled.scala 287:21]
  reg [2:0] sels_0; // @[Mux.scala 32:23]
  reg [31:0] _RAND_0;
  reg [2:0] sels_1; // @[Mux.scala 32:23]
  reg [31:0] _RAND_1;
  wire  _T_3; // @[Mux.scala 45:28]
  wire  _GEN_7; // @[Mux.scala 45:41]
  wire  _GEN_8; // @[Mux.scala 45:41]
  wire  _T_4; // @[Mux.scala 45:28]
  wire  _GEN_12; // @[Mux.scala 45:41]
  wire [31:0] _GEN_15; // @[Mux.scala 45:41]
  wire  _GEN_16; // @[Mux.scala 45:41]
  wire  _GEN_17; // @[Mux.scala 45:41]
  wire  _T_5; // @[Mux.scala 45:28]
  wire  _GEN_21; // @[Mux.scala 45:41]
  wire [31:0] _GEN_24; // @[Mux.scala 45:41]
  wire  _GEN_25; // @[Mux.scala 45:41]
  wire  _GEN_26; // @[Mux.scala 45:41]
  wire  _T_6; // @[Mux.scala 45:28]
  wire  _GEN_30; // @[Mux.scala 45:41]
  wire [31:0] _GEN_33; // @[Mux.scala 45:41]
  wire  _GEN_34; // @[Mux.scala 45:41]
  wire  _T_7; // @[Mux.scala 45:28]
  wire  _T_8; // @[Mux.scala 40:46]
  wire [2:0] _T_10; // @[Mux.scala 41:29]
  wire  _T_11; // @[Mux.scala 45:28]
  wire  _T_12; // @[Mux.scala 45:28]
  wire  _T_13; // @[Mux.scala 45:28]
  wire  _T_17; // @[RegisterRouter.scala 40:39]
  wire  _T_18; // @[RegisterRouter.scala 40:26]
  wire  _T_19; // @[RegisterRouter.scala 42:29]
  wire  _T_62_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 290:17]
  wire [29:0] _T_26; // @[RegisterRouter.scala 48:19]
  wire [1:0] _T_66; // @[RegisterRouter.scala 59:16]
  wire  _T_68; // @[RegisterRouter.scala 59:16]
  wire  _T_20; // @[RegisterRouter.scala 42:26]
  wire [1:0] _T_29; // @[OneHot.scala 65:12]
  wire [1:0] _T_31; // @[Misc.scala 200:81]
  wire  _T_32; // @[Misc.scala 204:21]
  wire  _T_35; // @[Misc.scala 209:20]
  wire  _T_37; // @[Misc.scala 213:38]
  wire  _T_38; // @[Misc.scala 213:29]
  wire  _T_40; // @[Misc.scala 213:38]
  wire  _T_41; // @[Misc.scala 213:29]
  wire  _T_44; // @[Misc.scala 209:20]
  wire  _T_45; // @[Misc.scala 212:27]
  wire  _T_46; // @[Misc.scala 213:38]
  wire  _T_47; // @[Misc.scala 213:29]
  wire  _T_48; // @[Misc.scala 212:27]
  wire  _T_49; // @[Misc.scala 213:38]
  wire  _T_50; // @[Misc.scala 213:29]
  wire  _T_51; // @[Misc.scala 212:27]
  wire  _T_52; // @[Misc.scala 213:38]
  wire  _T_53; // @[Misc.scala 213:29]
  wire  _T_54; // @[Misc.scala 212:27]
  wire  _T_55; // @[Misc.scala 213:38]
  wire  _T_56; // @[Misc.scala 213:29]
  wire [3:0] _T_59; // @[Cat.scala 29:58]
  wire [3:0] _T_61; // @[RegisterRouter.scala 54:25]
  wire [7:0] _T_80; // @[Bitwise.scala 72:12]
  wire [7:0] _T_82; // @[Bitwise.scala 72:12]
  wire [7:0] _T_84; // @[Bitwise.scala 72:12]
  wire [7:0] _T_86; // @[Bitwise.scala 72:12]
  wire [31:0] _T_89; // @[Cat.scala 29:58]
  wire  _T_108; // @[RegisterRouter.scala 59:16]
  wire  _T_161; // @[RegisterRouter.scala 59:16]
  wire [1:0] _T_155; // @[OneHot.scala 58:35]
  wire  _T_178; // @[RegisterRouter.scala 59:16]
  wire  _T_185; // @[RegisterRouter.scala 59:16]
  wire  _T_186; // @[RegisterRouter.scala 59:16]
  wire  _T_115; // @[RegisterRouter.scala 59:16]
  wire  _T_180; // @[RegisterRouter.scala 59:16]
  wire  _T_181; // @[RegisterRouter.scala 59:16]
  wire  _T_138; // @[RegisterRouter.scala 59:16]
  wire  _GEN_101; // @[MuxLiteral.scala 48:10]
  wire [2:0] _GEN_103; // @[MuxLiteral.scala 48:10]
  wire [2:0] _T_235; // @[RegisterRouter.scala 59:16]
  wire  _T_236_bits_read; // @[Decoupled.scala 308:19 Decoupled.scala 309:14]
  wire  _T_236_valid; // @[Decoupled.scala 308:19 Decoupled.scala 310:15]
  wire  _T_239; // @[RegisterRouter.scala 65:29]
  Queue Queue ( // @[Decoupled.scala 287:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_read(Queue_io_enq_bits_read),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_extra(Queue_io_enq_bits_extra),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_read(Queue_io_deq_bits_read),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_extra(Queue_io_deq_bits_extra)
  );
  assign _T_3 = sels_0 == 3'h0; // @[Mux.scala 45:28]
  assign _GEN_7 = _T_3 & auto_stream_in_0_valid; // @[Mux.scala 45:41]
  assign _GEN_8 = _T_3 & auto_stream_out_0_ready; // @[Mux.scala 45:41]
  assign _T_4 = sels_0 == 3'h1; // @[Mux.scala 45:28]
  assign _GEN_12 = _T_4 ? auto_stream_in_1_bits_last : auto_stream_in_0_bits_last; // @[Mux.scala 45:41]
  assign _GEN_15 = _T_4 ? auto_stream_in_1_bits_data : auto_stream_in_0_bits_data; // @[Mux.scala 45:41]
  assign _GEN_16 = _T_4 ? auto_stream_in_1_valid : _GEN_7; // @[Mux.scala 45:41]
  assign _GEN_17 = _T_4 & auto_stream_out_0_ready; // @[Mux.scala 45:41]
  assign _T_5 = sels_0 == 3'h2; // @[Mux.scala 45:28]
  assign _GEN_21 = _T_5 ? auto_stream_in_2_bits_last : _GEN_12; // @[Mux.scala 45:41]
  assign _GEN_24 = _T_5 ? auto_stream_in_2_bits_data : _GEN_15; // @[Mux.scala 45:41]
  assign _GEN_25 = _T_5 ? auto_stream_in_2_valid : _GEN_16; // @[Mux.scala 45:41]
  assign _GEN_26 = _T_5 & auto_stream_out_0_ready; // @[Mux.scala 45:41]
  assign _T_6 = sels_0 == 3'h3; // @[Mux.scala 45:28]
  assign _GEN_30 = _T_6 ? 1'h0 : _GEN_21; // @[Mux.scala 45:41]
  assign _GEN_33 = _T_6 ? 32'hffffffff : _GEN_24; // @[Mux.scala 45:41]
  assign _GEN_34 = _T_6 | _GEN_25; // @[Mux.scala 45:41]
  assign _T_7 = sels_0 == 3'h4; // @[Mux.scala 45:28]
  assign _T_8 = sels_0 == sels_1; // @[Mux.scala 40:46]
  assign _T_10 = _T_8 ? 3'h5 : sels_1; // @[Mux.scala 41:29]
  assign _T_11 = _T_10 == 3'h0; // @[Mux.scala 45:28]
  assign _T_12 = _T_10 == 3'h1; // @[Mux.scala 45:28]
  assign _T_13 = _T_10 == 3'h2; // @[Mux.scala 45:28]
  assign _T_17 = auto_register_in_aw_valid & auto_register_in_w_valid; // @[RegisterRouter.scala 40:39]
  assign _T_18 = auto_register_in_ar_valid | _T_17; // @[RegisterRouter.scala 40:26]
  assign _T_19 = ~auto_register_in_ar_valid; // @[RegisterRouter.scala 42:29]
  assign _T_62_ready = Queue_io_enq_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 290:17]
  assign _T_26 = auto_register_in_ar_valid ? auto_register_in_ar_bits_addr : auto_register_in_aw_bits_addr; // @[RegisterRouter.scala 48:19]
  assign _T_66 = _T_26[3:2] & 2'h2; // @[RegisterRouter.scala 59:16]
  assign _T_68 = _T_66 == 2'h0; // @[RegisterRouter.scala 59:16]
  assign _T_20 = _T_62_ready & _T_19; // @[RegisterRouter.scala 42:26]
  assign _T_29 = 2'h1 << auto_register_in_ar_bits_size[0]; // @[OneHot.scala 65:12]
  assign _T_31 = _T_29 | 2'h1; // @[Misc.scala 200:81]
  assign _T_32 = auto_register_in_ar_bits_size >= 3'h2; // @[Misc.scala 204:21]
  assign _T_35 = ~auto_register_in_ar_bits_addr[1]; // @[Misc.scala 209:20]
  assign _T_37 = _T_31[1] & _T_35; // @[Misc.scala 213:38]
  assign _T_38 = _T_32 | _T_37; // @[Misc.scala 213:29]
  assign _T_40 = _T_31[1] & auto_register_in_ar_bits_addr[1]; // @[Misc.scala 213:38]
  assign _T_41 = _T_32 | _T_40; // @[Misc.scala 213:29]
  assign _T_44 = ~auto_register_in_ar_bits_addr[0]; // @[Misc.scala 209:20]
  assign _T_45 = _T_35 & _T_44; // @[Misc.scala 212:27]
  assign _T_46 = _T_31[0] & _T_45; // @[Misc.scala 213:38]
  assign _T_47 = _T_38 | _T_46; // @[Misc.scala 213:29]
  assign _T_48 = _T_35 & auto_register_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  assign _T_49 = _T_31[0] & _T_48; // @[Misc.scala 213:38]
  assign _T_50 = _T_38 | _T_49; // @[Misc.scala 213:29]
  assign _T_51 = auto_register_in_ar_bits_addr[1] & _T_44; // @[Misc.scala 212:27]
  assign _T_52 = _T_31[0] & _T_51; // @[Misc.scala 213:38]
  assign _T_53 = _T_41 | _T_52; // @[Misc.scala 213:29]
  assign _T_54 = auto_register_in_ar_bits_addr[1] & auto_register_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  assign _T_55 = _T_31[0] & _T_54; // @[Misc.scala 213:38]
  assign _T_56 = _T_41 | _T_55; // @[Misc.scala 213:29]
  assign _T_59 = {_T_56,_T_53,_T_50,_T_47}; // @[Cat.scala 29:58]
  assign _T_61 = auto_register_in_ar_valid ? _T_59 : auto_register_in_w_bits_strb; // @[RegisterRouter.scala 54:25]
  assign _T_80 = _T_61[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_82 = _T_61[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_84 = _T_61[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_86 = _T_61[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_89 = {_T_86,_T_84,_T_82,_T_80}; // @[Cat.scala 29:58]
  assign _T_108 = _T_89[2:0] == 3'h7; // @[RegisterRouter.scala 59:16]
  assign _T_161 = _T_18 & _T_62_ready; // @[RegisterRouter.scala 59:16]
  assign _T_155 = 2'h1 << _T_26[2]; // @[OneHot.scala 58:35]
  assign _T_178 = _T_161 & _T_19; // @[RegisterRouter.scala 59:16]
  assign _T_185 = _T_178 & _T_155[1]; // @[RegisterRouter.scala 59:16]
  assign _T_186 = _T_185 & _T_68; // @[RegisterRouter.scala 59:16]
  assign _T_115 = _T_186 & _T_108; // @[RegisterRouter.scala 59:16]
  assign _T_180 = _T_178 & _T_155[0]; // @[RegisterRouter.scala 59:16]
  assign _T_181 = _T_180 & _T_68; // @[RegisterRouter.scala 59:16]
  assign _T_138 = _T_181 & _T_108; // @[RegisterRouter.scala 59:16]
  assign _GEN_101 = _T_26[2] ? _T_68 : _T_68; // @[MuxLiteral.scala 48:10]
  assign _GEN_103 = _T_26[2] ? sels_1 : sels_0; // @[MuxLiteral.scala 48:10]
  assign _T_235 = _GEN_101 ? _GEN_103 : 3'h0; // @[RegisterRouter.scala 59:16]
  assign _T_236_bits_read = Queue_io_deq_bits_read; // @[Decoupled.scala 308:19 Decoupled.scala 309:14]
  assign _T_236_valid = Queue_io_deq_valid; // @[Decoupled.scala 308:19 Decoupled.scala 310:15]
  assign _T_239 = ~_T_236_bits_read; // @[RegisterRouter.scala 65:29]
  assign auto_register_in_aw_ready = _T_20 & auto_register_in_w_valid; // @[LazyModule.scala 173:31]
  assign auto_register_in_w_ready = _T_20 & auto_register_in_aw_valid; // @[LazyModule.scala 173:31]
  assign auto_register_in_b_valid = _T_236_valid & _T_239; // @[LazyModule.scala 173:31]
  assign auto_register_in_b_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_register_in_ar_ready = Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_register_in_r_valid = _T_236_valid & _T_236_bits_read; // @[LazyModule.scala 173:31]
  assign auto_register_in_r_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_register_in_r_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 173:31]
  assign auto_stream_in_2_ready = _T_13 | _GEN_26; // @[LazyModule.scala 173:31]
  assign auto_stream_in_1_ready = _T_12 | _GEN_17; // @[LazyModule.scala 173:31]
  assign auto_stream_in_0_ready = _T_11 | _GEN_8; // @[LazyModule.scala 173:31]
  assign auto_stream_out_0_valid = _T_7 | _GEN_34; // @[LazyModule.scala 173:49]
  assign auto_stream_out_0_bits_data = _T_7 ? 32'h0 : _GEN_33; // @[LazyModule.scala 173:49]
  assign auto_stream_out_0_bits_last = _T_7 ? 1'h0 : _GEN_30; // @[LazyModule.scala 173:49]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_register_in_ar_valid | _T_17; // @[Decoupled.scala 288:22]
  assign Queue_io_enq_bits_read = auto_register_in_ar_valid; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_data = {{29'd0}, _T_235}; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_extra = auto_register_in_ar_valid ? auto_register_in_ar_bits_id : auto_register_in_aw_bits_id; // @[Decoupled.scala 289:21]
  assign Queue_io_deq_ready = _T_236_bits_read ? auto_register_in_r_ready : auto_register_in_b_ready; // @[Decoupled.scala 311:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  sels_0 = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  sels_1 = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      sels_0 <= 3'h5;
    end else if (_T_138) begin
      sels_0 <= auto_register_in_w_bits_data[2:0];
    end
    if (reset) begin
      sels_1 <= 3'h5;
    end else if (_T_115) begin
      sels_1 <= auto_register_in_w_bits_data[2:0];
    end
  end
endmodule
module AXI4StreamMux_7(
  input         clock,
  input         reset,
  output        auto_register_in_aw_ready,
  input         auto_register_in_aw_valid,
  input         auto_register_in_aw_bits_id,
  input  [29:0] auto_register_in_aw_bits_addr,
  output        auto_register_in_w_ready,
  input         auto_register_in_w_valid,
  input  [31:0] auto_register_in_w_bits_data,
  input  [3:0]  auto_register_in_w_bits_strb,
  input         auto_register_in_b_ready,
  output        auto_register_in_b_valid,
  output        auto_register_in_b_bits_id,
  output        auto_register_in_ar_ready,
  input         auto_register_in_ar_valid,
  input         auto_register_in_ar_bits_id,
  input  [29:0] auto_register_in_ar_bits_addr,
  input  [2:0]  auto_register_in_ar_bits_size,
  input         auto_register_in_r_ready,
  output        auto_register_in_r_valid,
  output        auto_register_in_r_bits_id,
  output [31:0] auto_register_in_r_bits_data,
  output        auto_stream_in_ready,
  input         auto_stream_in_valid,
  input  [31:0] auto_stream_in_bits_data,
  input         auto_stream_in_bits_last,
  input         auto_stream_out_1_ready,
  output        auto_stream_out_1_valid,
  output [31:0] auto_stream_out_1_bits_data,
  output        auto_stream_out_1_bits_last
);
  wire  Queue_clock; // @[Decoupled.scala 287:21]
  wire  Queue_reset; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_read; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_enq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_extra; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_read; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_deq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_extra; // @[Decoupled.scala 287:21]
  reg  sels_0; // @[Mux.scala 32:23]
  reg [31:0] _RAND_0;
  reg  sels_1; // @[Mux.scala 32:23]
  reg [31:0] _RAND_1;
  wire  _T_3; // @[Mux.scala 45:28]
  wire  _T_4; // @[Mux.scala 40:46]
  wire  _T_6; // @[Mux.scala 41:29]
  wire  _T_7; // @[Mux.scala 45:28]
  wire  _T_9; // @[RegisterRouter.scala 40:39]
  wire  _T_10; // @[RegisterRouter.scala 40:26]
  wire  _T_11; // @[RegisterRouter.scala 42:29]
  wire  _T_54_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 290:17]
  wire [29:0] _T_18; // @[RegisterRouter.scala 48:19]
  wire [1:0] _T_58; // @[RegisterRouter.scala 59:16]
  wire  _T_60; // @[RegisterRouter.scala 59:16]
  wire  _T_12; // @[RegisterRouter.scala 42:26]
  wire [1:0] _T_21; // @[OneHot.scala 65:12]
  wire [1:0] _T_23; // @[Misc.scala 200:81]
  wire  _T_24; // @[Misc.scala 204:21]
  wire  _T_27; // @[Misc.scala 209:20]
  wire  _T_29; // @[Misc.scala 213:38]
  wire  _T_30; // @[Misc.scala 213:29]
  wire  _T_32; // @[Misc.scala 213:38]
  wire  _T_33; // @[Misc.scala 213:29]
  wire  _T_36; // @[Misc.scala 209:20]
  wire  _T_37; // @[Misc.scala 212:27]
  wire  _T_38; // @[Misc.scala 213:38]
  wire  _T_39; // @[Misc.scala 213:29]
  wire  _T_40; // @[Misc.scala 212:27]
  wire  _T_41; // @[Misc.scala 213:38]
  wire  _T_42; // @[Misc.scala 213:29]
  wire  _T_43; // @[Misc.scala 212:27]
  wire  _T_44; // @[Misc.scala 213:38]
  wire  _T_45; // @[Misc.scala 213:29]
  wire  _T_46; // @[Misc.scala 212:27]
  wire  _T_47; // @[Misc.scala 213:38]
  wire  _T_48; // @[Misc.scala 213:29]
  wire [3:0] _T_51; // @[Cat.scala 29:58]
  wire [3:0] _T_53; // @[RegisterRouter.scala 54:25]
  wire [7:0] _T_72; // @[Bitwise.scala 72:12]
  wire [7:0] _T_74; // @[Bitwise.scala 72:12]
  wire [7:0] _T_76; // @[Bitwise.scala 72:12]
  wire [7:0] _T_78; // @[Bitwise.scala 72:12]
  wire [31:0] _T_81; // @[Cat.scala 29:58]
  wire  _T_153; // @[RegisterRouter.scala 59:16]
  wire [1:0] _T_147; // @[OneHot.scala 58:35]
  wire  _T_170; // @[RegisterRouter.scala 59:16]
  wire  _T_177; // @[RegisterRouter.scala 59:16]
  wire  _T_178; // @[RegisterRouter.scala 59:16]
  wire  _T_107; // @[RegisterRouter.scala 59:16]
  wire  _GEN_18; // @[RegField.scala 134:88]
  wire  _T_172; // @[RegisterRouter.scala 59:16]
  wire  _T_173; // @[RegisterRouter.scala 59:16]
  wire  _T_130; // @[RegisterRouter.scala 59:16]
  wire  _GEN_19; // @[RegField.scala 134:88]
  wire  _GEN_29; // @[MuxLiteral.scala 48:10]
  wire  _GEN_31; // @[MuxLiteral.scala 48:10]
  wire  _T_227; // @[RegisterRouter.scala 59:16]
  wire  _T_228_bits_read; // @[Decoupled.scala 308:19 Decoupled.scala 309:14]
  wire  _T_228_valid; // @[Decoupled.scala 308:19 Decoupled.scala 310:15]
  wire  _T_231; // @[RegisterRouter.scala 65:29]
  Queue Queue ( // @[Decoupled.scala 287:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_read(Queue_io_enq_bits_read),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_extra(Queue_io_enq_bits_extra),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_read(Queue_io_deq_bits_read),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_extra(Queue_io_deq_bits_extra)
  );
  assign _T_3 = ~sels_0; // @[Mux.scala 45:28]
  assign _T_4 = sels_0 == sels_1; // @[Mux.scala 40:46]
  assign _T_6 = _T_4 | sels_1; // @[Mux.scala 41:29]
  assign _T_7 = ~_T_6; // @[Mux.scala 45:28]
  assign _T_9 = auto_register_in_aw_valid & auto_register_in_w_valid; // @[RegisterRouter.scala 40:39]
  assign _T_10 = auto_register_in_ar_valid | _T_9; // @[RegisterRouter.scala 40:26]
  assign _T_11 = ~auto_register_in_ar_valid; // @[RegisterRouter.scala 42:29]
  assign _T_54_ready = Queue_io_enq_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 290:17]
  assign _T_18 = auto_register_in_ar_valid ? auto_register_in_ar_bits_addr : auto_register_in_aw_bits_addr; // @[RegisterRouter.scala 48:19]
  assign _T_58 = _T_18[3:2] & 2'h2; // @[RegisterRouter.scala 59:16]
  assign _T_60 = _T_58 == 2'h0; // @[RegisterRouter.scala 59:16]
  assign _T_12 = _T_54_ready & _T_11; // @[RegisterRouter.scala 42:26]
  assign _T_21 = 2'h1 << auto_register_in_ar_bits_size[0]; // @[OneHot.scala 65:12]
  assign _T_23 = _T_21 | 2'h1; // @[Misc.scala 200:81]
  assign _T_24 = auto_register_in_ar_bits_size >= 3'h2; // @[Misc.scala 204:21]
  assign _T_27 = ~auto_register_in_ar_bits_addr[1]; // @[Misc.scala 209:20]
  assign _T_29 = _T_23[1] & _T_27; // @[Misc.scala 213:38]
  assign _T_30 = _T_24 | _T_29; // @[Misc.scala 213:29]
  assign _T_32 = _T_23[1] & auto_register_in_ar_bits_addr[1]; // @[Misc.scala 213:38]
  assign _T_33 = _T_24 | _T_32; // @[Misc.scala 213:29]
  assign _T_36 = ~auto_register_in_ar_bits_addr[0]; // @[Misc.scala 209:20]
  assign _T_37 = _T_27 & _T_36; // @[Misc.scala 212:27]
  assign _T_38 = _T_23[0] & _T_37; // @[Misc.scala 213:38]
  assign _T_39 = _T_30 | _T_38; // @[Misc.scala 213:29]
  assign _T_40 = _T_27 & auto_register_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  assign _T_41 = _T_23[0] & _T_40; // @[Misc.scala 213:38]
  assign _T_42 = _T_30 | _T_41; // @[Misc.scala 213:29]
  assign _T_43 = auto_register_in_ar_bits_addr[1] & _T_36; // @[Misc.scala 212:27]
  assign _T_44 = _T_23[0] & _T_43; // @[Misc.scala 213:38]
  assign _T_45 = _T_33 | _T_44; // @[Misc.scala 213:29]
  assign _T_46 = auto_register_in_ar_bits_addr[1] & auto_register_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  assign _T_47 = _T_23[0] & _T_46; // @[Misc.scala 213:38]
  assign _T_48 = _T_33 | _T_47; // @[Misc.scala 213:29]
  assign _T_51 = {_T_48,_T_45,_T_42,_T_39}; // @[Cat.scala 29:58]
  assign _T_53 = auto_register_in_ar_valid ? _T_51 : auto_register_in_w_bits_strb; // @[RegisterRouter.scala 54:25]
  assign _T_72 = _T_53[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_74 = _T_53[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_76 = _T_53[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_78 = _T_53[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_81 = {_T_78,_T_76,_T_74,_T_72}; // @[Cat.scala 29:58]
  assign _T_153 = _T_10 & _T_54_ready; // @[RegisterRouter.scala 59:16]
  assign _T_147 = 2'h1 << _T_18[2]; // @[OneHot.scala 58:35]
  assign _T_170 = _T_153 & _T_11; // @[RegisterRouter.scala 59:16]
  assign _T_177 = _T_170 & _T_147[1]; // @[RegisterRouter.scala 59:16]
  assign _T_178 = _T_177 & _T_60; // @[RegisterRouter.scala 59:16]
  assign _T_107 = _T_178 & _T_81[0]; // @[RegisterRouter.scala 59:16]
  assign _GEN_18 = _T_107 ? auto_register_in_w_bits_data[0] : sels_1; // @[RegField.scala 134:88]
  assign _T_172 = _T_170 & _T_147[0]; // @[RegisterRouter.scala 59:16]
  assign _T_173 = _T_172 & _T_60; // @[RegisterRouter.scala 59:16]
  assign _T_130 = _T_173 & _T_81[0]; // @[RegisterRouter.scala 59:16]
  assign _GEN_19 = _T_130 ? auto_register_in_w_bits_data[0] : sels_0; // @[RegField.scala 134:88]
  assign _GEN_29 = _T_18[2] ? _T_60 : _T_60; // @[MuxLiteral.scala 48:10]
  assign _GEN_31 = _T_18[2] ? sels_1 : sels_0; // @[MuxLiteral.scala 48:10]
  assign _T_227 = _GEN_29 & _GEN_31; // @[RegisterRouter.scala 59:16]
  assign _T_228_bits_read = Queue_io_deq_bits_read; // @[Decoupled.scala 308:19 Decoupled.scala 309:14]
  assign _T_228_valid = Queue_io_deq_valid; // @[Decoupled.scala 308:19 Decoupled.scala 310:15]
  assign _T_231 = ~_T_228_bits_read; // @[RegisterRouter.scala 65:29]
  assign auto_register_in_aw_ready = _T_12 & auto_register_in_w_valid; // @[LazyModule.scala 173:31]
  assign auto_register_in_w_ready = _T_12 & auto_register_in_aw_valid; // @[LazyModule.scala 173:31]
  assign auto_register_in_b_valid = _T_228_valid & _T_231; // @[LazyModule.scala 173:31]
  assign auto_register_in_b_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_register_in_ar_ready = Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_register_in_r_valid = _T_228_valid & _T_228_bits_read; // @[LazyModule.scala 173:31]
  assign auto_register_in_r_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_register_in_r_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 173:31]
  assign auto_stream_in_ready = _T_7 ? auto_stream_out_1_ready : _T_3; // @[LazyModule.scala 173:31]
  assign auto_stream_out_1_valid = _T_7 & auto_stream_in_valid; // @[LazyModule.scala 173:49]
  assign auto_stream_out_1_bits_data = auto_stream_in_bits_data; // @[LazyModule.scala 173:49]
  assign auto_stream_out_1_bits_last = auto_stream_in_bits_last; // @[LazyModule.scala 173:49]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_register_in_ar_valid | _T_9; // @[Decoupled.scala 288:22]
  assign Queue_io_enq_bits_read = auto_register_in_ar_valid; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_data = {{31'd0}, _T_227}; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_extra = auto_register_in_ar_valid ? auto_register_in_ar_bits_id : auto_register_in_aw_bits_id; // @[Decoupled.scala 289:21]
  assign Queue_io_deq_ready = _T_228_bits_read ? auto_register_in_r_ready : auto_register_in_b_ready; // @[Decoupled.scala 311:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  sels_0 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  sels_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    sels_0 <= reset | _GEN_19;
    sels_1 <= reset | _GEN_18;
  end
endmodule
module Accumulator(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [15:0] io_in_bits,
  input         io_lastIn,
  input  [6:0]  io_accDepthReg,
  input  [16:0] io_accWindowsReg,
  input         io_out_ready,
  output        io_out_valid,
  output [15:0] io_out_bits,
  output        io_lastOut
);
  reg [31:0] mem [0:63]; // @[Accumulator.scala 35:24]
  reg [31:0] _RAND_0;
  wire [31:0] mem__T_175_data; // @[Accumulator.scala 35:24]
  wire [5:0] mem__T_175_addr; // @[Accumulator.scala 35:24]
  wire [31:0] mem__T_221_data; // @[Accumulator.scala 35:24]
  wire [5:0] mem__T_221_addr; // @[Accumulator.scala 35:24]
  wire  mem__T_221_mask; // @[Accumulator.scala 35:24]
  wire  mem__T_221_en; // @[Accumulator.scala 35:24]
  reg  mem__T_175_en_pipe_0;
  reg [31:0] _RAND_1;
  reg [5:0] mem__T_175_addr_pipe_0;
  reg [31:0] _RAND_2;
  wire  readEn; // @[Decoupled.scala 40:37]
  reg  writeEn; // @[Accumulator.scala 38:24]
  reg [31:0] _RAND_3;
  reg [15:0] inDelayed; // @[Accumulator.scala 39:26]
  reg [31:0] _RAND_4;
  reg [15:0] cntWindows; // @[Accumulator.scala 40:27]
  reg [31:0] _RAND_5;
  reg [5:0] cntLoad; // @[Accumulator.scala 41:24]
  reg [31:0] _RAND_6;
  reg [5:0] cntAcc; // @[Accumulator.scala 42:23]
  reg [31:0] _RAND_7;
  reg [2:0] state; // @[Accumulator.scala 50:22]
  reg [31:0] _RAND_8;
  reg [2:0] statePrev; // @[Accumulator.scala 51:26]
  reg [31:0] _RAND_9;
  reg  last; // @[Accumulator.scala 53:21]
  reg [31:0] _RAND_10;
  wire  _T_3; // @[Conditional.scala 37:30]
  wire  _T_7; // @[Conditional.scala 37:30]
  wire [6:0] _T_9; // @[Accumulator.scala 66:40]
  wire [6:0] _GEN_34; // @[Accumulator.scala 66:20]
  wire  _T_10; // @[Accumulator.scala 66:20]
  wire  _T_12; // @[Accumulator.scala 66:47]
  wire  _T_13; // @[Accumulator.scala 66:63]
  wire  _T_21; // @[Conditional.scala 37:30]
  wire  _T_23; // @[Accumulator.scala 75:26]
  wire  _T_24; // @[Accumulator.scala 77:15]
  wire  _GEN_3; // @[Accumulator.scala 77:30]
  wire [16:0] _T_26; // @[Accumulator.scala 81:51]
  wire [16:0] _GEN_36; // @[Accumulator.scala 81:29]
  wire  _T_27; // @[Accumulator.scala 81:29]
  wire  _T_29; // @[Accumulator.scala 81:58]
  wire  _T_33; // @[Accumulator.scala 81:72]
  wire  _T_36; // @[Conditional.scala 37:30]
  wire [6:0] _GEN_38; // @[Accumulator.scala 90:26]
  wire  _T_41; // @[Accumulator.scala 90:26]
  wire  _T_42; // @[Decoupled.scala 40:37]
  wire  _T_43; // @[Accumulator.scala 90:53]
  wire  _T_46; // @[Accumulator.scala 90:80]
  wire  _T_47; // @[Accumulator.scala 90:70]
  wire  _T_54; // @[Accumulator.scala 93:70]
  wire  _T_58; // @[Accumulator.scala 93:86]
  wire  _T_61; // @[Conditional.scala 37:30]
  wire  _T_62; // @[Accumulator.scala 105:30]
  wire  _T_63; // @[Accumulator.scala 105:65]
  wire  loadingStates; // @[Accumulator.scala 105:55]
  wire  _T_64; // @[Accumulator.scala 106:34]
  wire  storingInitStates; // @[Accumulator.scala 106:56]
  wire  _T_66; // @[Accumulator.scala 107:26]
  wire  _T_67; // @[Accumulator.scala 107:62]
  wire  _T_68; // @[Accumulator.scala 107:49]
  wire  _T_69; // @[Accumulator.scala 107:98]
  wire  _T_71; // @[Accumulator.scala 107:122]
  wire  _T_72; // @[Accumulator.scala 107:84]
  wire  _T_75; // @[Accumulator.scala 107:191]
  wire  isTransit; // @[Accumulator.scala 107:153]
  wire  isOnlyOneFrame; // @[Accumulator.scala 108:47]
  reg  doNotScale; // @[Accumulator.scala 109:27]
  reg [31:0] _RAND_11;
  wire  _T_78; // @[Accumulator.scala 110:38]
  wire  isPrevStoreAndAcc; // @[Accumulator.scala 110:62]
  wire  _GEN_19; // @[Accumulator.scala 116:24]
  wire  _T_88; // @[Accumulator.scala 119:15]
  wire  _T_89; // @[Accumulator.scala 123:28]
  wire  _T_90; // @[Accumulator.scala 123:45]
  wire  _T_91; // @[Accumulator.scala 123:42]
  wire  _T_92; // @[Accumulator.scala 123:64]
  wire [31:0] readVal; // @[Accumulator.scala 43:21 Accumulator.scala 172:11]
  wire [31:0] _GEN_44; // @[FixedPointTypeClass.scala 20:58]
  wire [31:0] _T_95; // @[FixedPointTypeClass.scala 20:58]
  wire [31:0] _GEN_21; // @[Accumulator.scala 123:83]
  wire [5:0] _T_98; // @[Accumulator.scala 130:22]
  wire  _T_99; // @[Accumulator.scala 133:23]
  wire [5:0] _T_101; // @[Accumulator.scala 134:24]
  wire [15:0] _T_111; // @[Accumulator.scala 142:30]
  wire  _T_115; // @[Accumulator.scala 145:49]
  wire  bools_0; // @[Accumulator.scala 159:39]
  wire  bools_1; // @[Accumulator.scala 159:39]
  wire  bools_2; // @[Accumulator.scala 159:39]
  wire  bools_3; // @[Accumulator.scala 159:39]
  wire  bools_4; // @[Accumulator.scala 159:39]
  wire  bools_5; // @[Accumulator.scala 159:39]
  wire  _T_116; // @[Accumulator.scala 160:46]
  wire [5:0] loadAddressBeforeBitReverse; // @[Accumulator.scala 160:40]
  wire [1:0] _T_123; // @[Cat.scala 29:58]
  wire [2:0] _T_130; // @[Cat.scala 29:58]
  wire [3:0] _T_140; // @[Cat.scala 29:58]
  wire [4:0] _T_153; // @[Cat.scala 29:58]
  wire [5:0] _T_169; // @[Cat.scala 29:58]
  wire [5:0] _T_170; // @[Mux.scala 87:16]
  wire [5:0] _T_171; // @[Mux.scala 87:16]
  wire [5:0] _T_172; // @[Mux.scala 87:16]
  wire [5:0] _T_173; // @[Mux.scala 87:16]
  wire [5:0] _T_174; // @[Mux.scala 87:16]
  wire [5:0] loadAddress; // @[Mux.scala 87:16]
  wire [5:0] readAddress; // @[Accumulator.scala 167:24]
  wire  _T_181; // @[CircuitMath.scala 37:22]
  wire  _T_184; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_188; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_189; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_193; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_194; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_195; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_196; // @[Cat.scala 29:58]
  wire  _T_199; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_203; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_204; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_208; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_209; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_210; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_211; // @[Cat.scala 29:58]
  wire [2:0] _T_212; // @[CircuitMath.scala 38:21]
  wire [3:0] _T_213; // @[Cat.scala 29:58]
  wire [3:0] _T_214; // @[CircuitMath.scala 38:21]
  wire [4:0] _T_215; // @[Cat.scala 29:58]
  wire [31:0] _T_216; // @[FixedPointTypeClass.scala 118:51]
  wire [31:0] _T_217; // @[Accumulator.scala 178:17]
  reg [5:0] _T_218; // @[Accumulator.scala 184:22]
  reg [31:0] _RAND_12;
  wire [31:0] writeVal; // @[Accumulator.scala 44:22 Accumulator.scala 124:14 Accumulator.scala 127:14]
  reg  _T_222; // @[Accumulator.scala 187:26]
  reg [31:0] _RAND_13;
  wire  _T_223; // @[Accumulator.scala 187:51]
  reg [5:0] _T_225; // @[Accumulator.scala 188:27]
  reg [31:0] _RAND_14;
  wire [6:0] _GEN_47; // @[Accumulator.scala 188:57]
  wire  _T_228; // @[Accumulator.scala 188:57]
  wire  _T_230; // @[Accumulator.scala 188:84]
  assign mem__T_175_addr = mem__T_175_addr_pipe_0;
  assign mem__T_175_data = mem[mem__T_175_addr]; // @[Accumulator.scala 35:24]
  assign mem__T_221_data = writeVal;
  assign mem__T_221_addr = _T_218;
  assign mem__T_221_mask = 1'h1;
  assign mem__T_221_en = writeEn;
  assign readEn = io_in_ready & io_in_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = 3'h0 == state; // @[Conditional.scala 37:30]
  assign _T_7 = 3'h1 == state; // @[Conditional.scala 37:30]
  assign _T_9 = io_accDepthReg - 7'h1; // @[Accumulator.scala 66:40]
  assign _GEN_34 = {{1'd0}, cntAcc}; // @[Accumulator.scala 66:20]
  assign _T_10 = _GEN_34 == _T_9; // @[Accumulator.scala 66:20]
  assign _T_12 = _T_10 & readEn; // @[Accumulator.scala 66:47]
  assign _T_13 = _T_12 & io_lastIn; // @[Accumulator.scala 66:63]
  assign _T_21 = 3'h2 == state; // @[Conditional.scala 37:30]
  assign _T_23 = readEn & io_lastIn; // @[Accumulator.scala 75:26]
  assign _T_24 = ~io_out_ready; // @[Accumulator.scala 77:15]
  assign _GEN_3 = _T_24 | last; // @[Accumulator.scala 77:30]
  assign _T_26 = io_accWindowsReg - 17'h1; // @[Accumulator.scala 81:51]
  assign _GEN_36 = {{1'd0}, cntWindows}; // @[Accumulator.scala 81:29]
  assign _T_27 = _GEN_36 == _T_26; // @[Accumulator.scala 81:29]
  assign _T_29 = _T_27 & readEn; // @[Accumulator.scala 81:58]
  assign _T_33 = _T_29 & _T_10; // @[Accumulator.scala 81:72]
  assign _T_36 = 3'h3 == state; // @[Conditional.scala 37:30]
  assign _GEN_38 = {{1'd0}, cntLoad}; // @[Accumulator.scala 90:26]
  assign _T_41 = _GEN_38 == _T_9; // @[Accumulator.scala 90:26]
  assign _T_42 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  assign _T_43 = _T_41 & _T_42; // @[Accumulator.scala 90:53]
  assign _T_46 = _GEN_34 < _T_9; // @[Accumulator.scala 90:80]
  assign _T_47 = _T_43 & _T_46; // @[Accumulator.scala 90:70]
  assign _T_54 = _T_43 & readEn; // @[Accumulator.scala 93:70]
  assign _T_58 = _T_54 & _T_10; // @[Accumulator.scala 93:86]
  assign _T_61 = 3'h4 == state; // @[Conditional.scala 37:30]
  assign _T_62 = state == 3'h3; // @[Accumulator.scala 105:30]
  assign _T_63 = state == 3'h4; // @[Accumulator.scala 105:65]
  assign loadingStates = _T_62 | _T_63; // @[Accumulator.scala 105:55]
  assign _T_64 = state == 3'h1; // @[Accumulator.scala 106:34]
  assign storingInitStates = _T_64 | _T_62; // @[Accumulator.scala 106:56]
  assign _T_66 = state == 3'h2; // @[Accumulator.scala 107:26]
  assign _T_67 = statePrev == 3'h1; // @[Accumulator.scala 107:62]
  assign _T_68 = _T_66 & _T_67; // @[Accumulator.scala 107:49]
  assign _T_69 = statePrev == 3'h3; // @[Accumulator.scala 107:98]
  assign _T_71 = _T_69 & _T_64; // @[Accumulator.scala 107:122]
  assign _T_72 = _T_68 | _T_71; // @[Accumulator.scala 107:84]
  assign _T_75 = _T_69 & _T_66; // @[Accumulator.scala 107:191]
  assign isTransit = _T_72 | _T_75; // @[Accumulator.scala 107:153]
  assign isOnlyOneFrame = _T_63 & _T_67; // @[Accumulator.scala 108:47]
  assign _T_78 = statePrev == 3'h2; // @[Accumulator.scala 110:38]
  assign isPrevStoreAndAcc = _T_78 & _T_62; // @[Accumulator.scala 110:62]
  assign _GEN_19 = isOnlyOneFrame | doNotScale; // @[Accumulator.scala 116:24]
  assign _T_88 = state == 3'h0; // @[Accumulator.scala 119:15]
  assign _T_89 = storingInitStates | isTransit; // @[Accumulator.scala 123:28]
  assign _T_90 = ~isPrevStoreAndAcc; // @[Accumulator.scala 123:45]
  assign _T_91 = _T_89 & _T_90; // @[Accumulator.scala 123:42]
  assign _T_92 = _T_91 | isOnlyOneFrame; // @[Accumulator.scala 123:64]
  assign readVal = mem__T_175_data; // @[Accumulator.scala 43:21 Accumulator.scala 172:11]
  assign _GEN_44 = {{16{inDelayed[15]}},inDelayed}; // @[FixedPointTypeClass.scala 20:58]
  assign _T_95 = $signed(_GEN_44) + $signed(readVal); // @[FixedPointTypeClass.scala 20:58]
  assign _GEN_21 = _T_92 ? $signed({{16{inDelayed[15]}},inDelayed}) : $signed(_T_95); // @[Accumulator.scala 123:83]
  assign _T_98 = cntAcc + 6'h1; // @[Accumulator.scala 130:22]
  assign _T_99 = loadingStates & io_out_ready; // @[Accumulator.scala 133:23]
  assign _T_101 = cntLoad + 6'h1; // @[Accumulator.scala 134:24]
  assign _T_111 = cntWindows + 16'h1; // @[Accumulator.scala 142:30]
  assign _T_115 = _T_27 & _T_12; // @[Accumulator.scala 145:49]
  assign bools_0 = 7'h2 == io_accDepthReg; // @[Accumulator.scala 159:39]
  assign bools_1 = 7'h4 == io_accDepthReg; // @[Accumulator.scala 159:39]
  assign bools_2 = 7'h8 == io_accDepthReg; // @[Accumulator.scala 159:39]
  assign bools_3 = 7'h10 == io_accDepthReg; // @[Accumulator.scala 159:39]
  assign bools_4 = 7'h20 == io_accDepthReg; // @[Accumulator.scala 159:39]
  assign bools_5 = 7'h40 == io_accDepthReg; // @[Accumulator.scala 159:39]
  assign _T_116 = last & io_out_ready; // @[Accumulator.scala 160:46]
  assign loadAddressBeforeBitReverse = _T_116 ? _T_101 : cntLoad; // @[Accumulator.scala 160:40]
  assign _T_123 = {loadAddressBeforeBitReverse[0],loadAddressBeforeBitReverse[1]}; // @[Cat.scala 29:58]
  assign _T_130 = {loadAddressBeforeBitReverse[0],loadAddressBeforeBitReverse[1],loadAddressBeforeBitReverse[2]}; // @[Cat.scala 29:58]
  assign _T_140 = {loadAddressBeforeBitReverse[0],loadAddressBeforeBitReverse[1],loadAddressBeforeBitReverse[2],loadAddressBeforeBitReverse[3]}; // @[Cat.scala 29:58]
  assign _T_153 = {loadAddressBeforeBitReverse[0],loadAddressBeforeBitReverse[1],loadAddressBeforeBitReverse[2],loadAddressBeforeBitReverse[3],loadAddressBeforeBitReverse[4]}; // @[Cat.scala 29:58]
  assign _T_169 = {loadAddressBeforeBitReverse[0],loadAddressBeforeBitReverse[1],loadAddressBeforeBitReverse[2],loadAddressBeforeBitReverse[3],loadAddressBeforeBitReverse[4],loadAddressBeforeBitReverse[5]}; // @[Cat.scala 29:58]
  assign _T_170 = bools_5 ? _T_169 : 6'h0; // @[Mux.scala 87:16]
  assign _T_171 = bools_4 ? {{1'd0}, _T_153} : _T_170; // @[Mux.scala 87:16]
  assign _T_172 = bools_3 ? {{2'd0}, _T_140} : _T_171; // @[Mux.scala 87:16]
  assign _T_173 = bools_2 ? {{3'd0}, _T_130} : _T_172; // @[Mux.scala 87:16]
  assign _T_174 = bools_1 ? {{4'd0}, _T_123} : _T_173; // @[Mux.scala 87:16]
  assign loadAddress = bools_0 ? {{5'd0}, loadAddressBeforeBitReverse[0]} : _T_174; // @[Mux.scala 87:16]
  assign readAddress = loadingStates ? loadAddress : cntAcc; // @[Accumulator.scala 167:24]
  assign _T_181 = io_accWindowsReg[15:8] != 8'h0; // @[CircuitMath.scala 37:22]
  assign _T_184 = io_accWindowsReg[15:12] != 4'h0; // @[CircuitMath.scala 37:22]
  assign _T_188 = io_accWindowsReg[14] ? 2'h2 : {{1'd0}, io_accWindowsReg[13]}; // @[CircuitMath.scala 32:10]
  assign _T_189 = io_accWindowsReg[15] ? 2'h3 : _T_188; // @[CircuitMath.scala 32:10]
  assign _T_193 = io_accWindowsReg[10] ? 2'h2 : {{1'd0}, io_accWindowsReg[9]}; // @[CircuitMath.scala 32:10]
  assign _T_194 = io_accWindowsReg[11] ? 2'h3 : _T_193; // @[CircuitMath.scala 32:10]
  assign _T_195 = _T_184 ? _T_189 : _T_194; // @[CircuitMath.scala 38:21]
  assign _T_196 = {_T_184,_T_195}; // @[Cat.scala 29:58]
  assign _T_199 = io_accWindowsReg[7:4] != 4'h0; // @[CircuitMath.scala 37:22]
  assign _T_203 = io_accWindowsReg[6] ? 2'h2 : {{1'd0}, io_accWindowsReg[5]}; // @[CircuitMath.scala 32:10]
  assign _T_204 = io_accWindowsReg[7] ? 2'h3 : _T_203; // @[CircuitMath.scala 32:10]
  assign _T_208 = io_accWindowsReg[2] ? 2'h2 : {{1'd0}, io_accWindowsReg[1]}; // @[CircuitMath.scala 32:10]
  assign _T_209 = io_accWindowsReg[3] ? 2'h3 : _T_208; // @[CircuitMath.scala 32:10]
  assign _T_210 = _T_199 ? _T_204 : _T_209; // @[CircuitMath.scala 38:21]
  assign _T_211 = {_T_199,_T_210}; // @[Cat.scala 29:58]
  assign _T_212 = _T_181 ? _T_196 : _T_211; // @[CircuitMath.scala 38:21]
  assign _T_213 = {_T_181,_T_212}; // @[Cat.scala 29:58]
  assign _T_214 = io_accWindowsReg[16] ? 4'h0 : _T_213; // @[CircuitMath.scala 38:21]
  assign _T_215 = {io_accWindowsReg[16],_T_214}; // @[Cat.scala 29:58]
  assign _T_216 = $signed(readVal) >>> _T_215; // @[FixedPointTypeClass.scala 118:51]
  assign _T_217 = doNotScale ? $signed(readVal) : $signed(_T_216); // @[Accumulator.scala 178:17]
  assign writeVal = _GEN_21; // @[Accumulator.scala 44:22 Accumulator.scala 124:14 Accumulator.scala 127:14]
  assign _T_223 = state != 3'h0; // @[Accumulator.scala 187:51]
  assign _GEN_47 = {{1'd0}, _T_225}; // @[Accumulator.scala 188:57]
  assign _T_228 = _GEN_47 == _T_9; // @[Accumulator.scala 188:57]
  assign _T_230 = _T_228 & _T_42; // @[Accumulator.scala 188:84]
  assign io_in_ready = ~loadingStates; // @[Accumulator.scala 196:18]
  assign io_out_valid = _T_222 & _T_223; // @[Accumulator.scala 187:16]
  assign io_out_bits = _T_217[15:0]; // @[Accumulator.scala 190:16]
  assign io_lastOut = _T_230 & _T_63; // @[Accumulator.scala 188:16]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    mem[initvar] = _RAND_0[31:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  mem__T_175_en_pipe_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  mem__T_175_addr_pipe_0 = _RAND_2[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  writeEn = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  inDelayed = _RAND_4[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  cntWindows = _RAND_5[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  cntLoad = _RAND_6[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  cntAcc = _RAND_7[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  state = _RAND_8[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  statePrev = _RAND_9[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  last = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  doNotScale = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_218 = _RAND_12[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_222 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_225 = _RAND_14[5:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(mem__T_221_en & mem__T_221_mask) begin
      mem[mem__T_221_addr] <= mem__T_221_data; // @[Accumulator.scala 35:24]
    end
    mem__T_175_en_pipe_0 <= 1'h1;
    if (loadingStates) begin
      if (bools_0) begin
        mem__T_175_addr_pipe_0 <= {{5'd0}, loadAddressBeforeBitReverse[0]};
      end else if (bools_1) begin
        mem__T_175_addr_pipe_0 <= {{4'd0}, _T_123};
      end else if (bools_2) begin
        mem__T_175_addr_pipe_0 <= {{3'd0}, _T_130};
      end else if (bools_3) begin
        mem__T_175_addr_pipe_0 <= {{2'd0}, _T_140};
      end else if (bools_4) begin
        mem__T_175_addr_pipe_0 <= {{1'd0}, _T_153};
      end else if (bools_5) begin
        mem__T_175_addr_pipe_0 <= _T_169;
      end else begin
        mem__T_175_addr_pipe_0 <= 6'h0;
      end
    end else begin
      mem__T_175_addr_pipe_0 <= cntAcc;
    end
    if (reset) begin
      writeEn <= 1'h0;
    end else begin
      writeEn <= readEn;
    end
    inDelayed <= io_in_bits;
    if (reset) begin
      cntWindows <= 16'h0;
    end else if (_T_115) begin
      cntWindows <= 16'h0;
    end else if (_T_12) begin
      cntWindows <= _T_111;
    end
    if (reset) begin
      cntLoad <= 6'h0;
    end else if (_T_43) begin
      cntLoad <= 6'h0;
    end else if (_T_99) begin
      cntLoad <= _T_101;
    end else if (_T_99) begin
      cntLoad <= _T_101;
    end
    if (reset) begin
      cntAcc <= 6'h0;
    end else if (_T_12) begin
      cntAcc <= 6'h0;
    end else if (readEn) begin
      cntAcc <= _T_98;
    end
    if (reset) begin
      state <= 3'h0;
    end else if (_T_3) begin
      if (readEn) begin
        state <= 3'h1;
      end
    end else if (_T_7) begin
      if (_T_13) begin
        state <= 3'h4;
      end else if (_T_12) begin
        state <= 3'h2;
      end
    end else if (_T_21) begin
      if (_T_23) begin
        state <= 3'h4;
      end else if (_T_33) begin
        state <= 3'h3;
      end
    end else if (_T_36) begin
      if (_T_23) begin
        state <= 3'h4;
      end else if (_T_47) begin
        state <= 3'h1;
      end else if (_T_58) begin
        state <= 3'h2;
      end
    end else if (_T_61) begin
      if (io_lastOut) begin
        state <= 3'h0;
      end
    end
    if (reset) begin
      statePrev <= 3'h0;
    end else begin
      statePrev <= state;
    end
    if (reset) begin
      last <= 1'h0;
    end else if (_T_3) begin
      last <= 1'h0;
    end else if (!(_T_7)) begin
      if (_T_21) begin
        if (_T_23) begin
          last <= _GEN_3;
        end
      end
    end
    if (reset) begin
      doNotScale <= 1'h0;
    end else if (_T_88) begin
      doNotScale <= 1'h0;
    end else begin
      doNotScale <= _GEN_19;
    end
    _T_218 <= cntAcc;
    _T_222 <= _T_62 | _T_63;
    if (_T_116) begin
      _T_225 <= _T_101;
    end else begin
      _T_225 <= cntLoad;
    end
  end
endmodule
module AXI4AccumulatorBlock(
  input         clock,
  input         reset,
  output        auto_mem_in_aw_ready,
  input         auto_mem_in_aw_valid,
  input         auto_mem_in_aw_bits_id,
  input  [29:0] auto_mem_in_aw_bits_addr,
  output        auto_mem_in_w_ready,
  input         auto_mem_in_w_valid,
  input  [31:0] auto_mem_in_w_bits_data,
  input  [3:0]  auto_mem_in_w_bits_strb,
  input         auto_mem_in_b_ready,
  output        auto_mem_in_b_valid,
  output        auto_mem_in_b_bits_id,
  output        auto_mem_in_ar_ready,
  input         auto_mem_in_ar_valid,
  input         auto_mem_in_ar_bits_id,
  input  [29:0] auto_mem_in_ar_bits_addr,
  input  [2:0]  auto_mem_in_ar_bits_size,
  input         auto_mem_in_r_ready,
  output        auto_mem_in_r_valid,
  output        auto_mem_in_r_bits_id,
  output [31:0] auto_mem_in_r_bits_data,
  input         auto_master_out_ready,
  output        auto_master_out_valid,
  output [15:0] auto_master_out_bits_data,
  output        auto_master_out_bits_last,
  output        auto_slave_in_ready,
  input         auto_slave_in_valid,
  input  [31:0] auto_slave_in_bits_data,
  input         auto_slave_in_bits_last
);
  wire  acc_clock; // @[AccDspBlock.scala 39:21]
  wire  acc_reset; // @[AccDspBlock.scala 39:21]
  wire  acc_io_in_ready; // @[AccDspBlock.scala 39:21]
  wire  acc_io_in_valid; // @[AccDspBlock.scala 39:21]
  wire [15:0] acc_io_in_bits; // @[AccDspBlock.scala 39:21]
  wire  acc_io_lastIn; // @[AccDspBlock.scala 39:21]
  wire [6:0] acc_io_accDepthReg; // @[AccDspBlock.scala 39:21]
  wire [16:0] acc_io_accWindowsReg; // @[AccDspBlock.scala 39:21]
  wire  acc_io_out_ready; // @[AccDspBlock.scala 39:21]
  wire  acc_io_out_valid; // @[AccDspBlock.scala 39:21]
  wire [15:0] acc_io_out_bits; // @[AccDspBlock.scala 39:21]
  wire  acc_io_lastOut; // @[AccDspBlock.scala 39:21]
  wire  Queue_clock; // @[Decoupled.scala 287:21]
  wire  Queue_reset; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_read; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_enq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_extra; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_read; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_deq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_extra; // @[Decoupled.scala 287:21]
  reg [6:0] accDepth; // @[AccDspBlock.scala 42:34]
  reg [31:0] _RAND_0;
  reg [16:0] numWin; // @[AccDspBlock.scala 43:34]
  reg [31:0] _RAND_1;
  wire  _T_2; // @[RegisterRouter.scala 40:39]
  wire  _T_3; // @[RegisterRouter.scala 40:26]
  wire  _T_4; // @[RegisterRouter.scala 42:29]
  wire  _T_47_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 290:17]
  wire [29:0] _T_11; // @[RegisterRouter.scala 48:19]
  wire [1:0] _T_51; // @[RegisterRouter.scala 59:16]
  wire  _T_53; // @[RegisterRouter.scala 59:16]
  wire  _T_5; // @[RegisterRouter.scala 42:26]
  wire [1:0] _T_14; // @[OneHot.scala 65:12]
  wire [1:0] _T_16; // @[Misc.scala 200:81]
  wire  _T_17; // @[Misc.scala 204:21]
  wire  _T_20; // @[Misc.scala 209:20]
  wire  _T_22; // @[Misc.scala 213:38]
  wire  _T_23; // @[Misc.scala 213:29]
  wire  _T_25; // @[Misc.scala 213:38]
  wire  _T_26; // @[Misc.scala 213:29]
  wire  _T_29; // @[Misc.scala 209:20]
  wire  _T_30; // @[Misc.scala 212:27]
  wire  _T_31; // @[Misc.scala 213:38]
  wire  _T_32; // @[Misc.scala 213:29]
  wire  _T_33; // @[Misc.scala 212:27]
  wire  _T_34; // @[Misc.scala 213:38]
  wire  _T_35; // @[Misc.scala 213:29]
  wire  _T_36; // @[Misc.scala 212:27]
  wire  _T_37; // @[Misc.scala 213:38]
  wire  _T_38; // @[Misc.scala 213:29]
  wire  _T_39; // @[Misc.scala 212:27]
  wire  _T_40; // @[Misc.scala 213:38]
  wire  _T_41; // @[Misc.scala 213:29]
  wire [3:0] _T_44; // @[Cat.scala 29:58]
  wire [3:0] _T_46; // @[RegisterRouter.scala 54:25]
  wire [7:0] _T_65; // @[Bitwise.scala 72:12]
  wire [7:0] _T_67; // @[Bitwise.scala 72:12]
  wire [7:0] _T_69; // @[Bitwise.scala 72:12]
  wire [7:0] _T_71; // @[Bitwise.scala 72:12]
  wire [31:0] _T_74; // @[Cat.scala 29:58]
  wire  _T_93; // @[RegisterRouter.scala 59:16]
  wire  _T_146; // @[RegisterRouter.scala 59:16]
  wire [1:0] _T_140; // @[OneHot.scala 58:35]
  wire  _T_163; // @[RegisterRouter.scala 59:16]
  wire  _T_170; // @[RegisterRouter.scala 59:16]
  wire  _T_171; // @[RegisterRouter.scala 59:16]
  wire  _T_100; // @[RegisterRouter.scala 59:16]
  wire  _T_116; // @[RegisterRouter.scala 59:16]
  wire  _T_165; // @[RegisterRouter.scala 59:16]
  wire  _T_166; // @[RegisterRouter.scala 59:16]
  wire  _T_123; // @[RegisterRouter.scala 59:16]
  wire  _GEN_11; // @[MuxLiteral.scala 48:10]
  wire [16:0] _T_218_0; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [16:0] _GEN_13; // @[MuxLiteral.scala 48:10]
  wire [16:0] _T_220; // @[RegisterRouter.scala 59:16]
  wire  _T_221_bits_read; // @[Decoupled.scala 308:19 Decoupled.scala 309:14]
  wire  _T_221_valid; // @[Decoupled.scala 308:19 Decoupled.scala 310:15]
  wire  _T_224; // @[RegisterRouter.scala 65:29]
  wire [31:0] _T_228; // @[AccDspBlock.scala 63:48]
  Accumulator acc ( // @[AccDspBlock.scala 39:21]
    .clock(acc_clock),
    .reset(acc_reset),
    .io_in_ready(acc_io_in_ready),
    .io_in_valid(acc_io_in_valid),
    .io_in_bits(acc_io_in_bits),
    .io_lastIn(acc_io_lastIn),
    .io_accDepthReg(acc_io_accDepthReg),
    .io_accWindowsReg(acc_io_accWindowsReg),
    .io_out_ready(acc_io_out_ready),
    .io_out_valid(acc_io_out_valid),
    .io_out_bits(acc_io_out_bits),
    .io_lastOut(acc_io_lastOut)
  );
  Queue Queue ( // @[Decoupled.scala 287:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_read(Queue_io_enq_bits_read),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_extra(Queue_io_enq_bits_extra),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_read(Queue_io_deq_bits_read),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_extra(Queue_io_deq_bits_extra)
  );
  assign _T_2 = auto_mem_in_aw_valid & auto_mem_in_w_valid; // @[RegisterRouter.scala 40:39]
  assign _T_3 = auto_mem_in_ar_valid | _T_2; // @[RegisterRouter.scala 40:26]
  assign _T_4 = ~auto_mem_in_ar_valid; // @[RegisterRouter.scala 42:29]
  assign _T_47_ready = Queue_io_enq_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 290:17]
  assign _T_11 = auto_mem_in_ar_valid ? auto_mem_in_ar_bits_addr : auto_mem_in_aw_bits_addr; // @[RegisterRouter.scala 48:19]
  assign _T_51 = _T_11[3:2] & 2'h2; // @[RegisterRouter.scala 59:16]
  assign _T_53 = _T_51 == 2'h0; // @[RegisterRouter.scala 59:16]
  assign _T_5 = _T_47_ready & _T_4; // @[RegisterRouter.scala 42:26]
  assign _T_14 = 2'h1 << auto_mem_in_ar_bits_size[0]; // @[OneHot.scala 65:12]
  assign _T_16 = _T_14 | 2'h1; // @[Misc.scala 200:81]
  assign _T_17 = auto_mem_in_ar_bits_size >= 3'h2; // @[Misc.scala 204:21]
  assign _T_20 = ~auto_mem_in_ar_bits_addr[1]; // @[Misc.scala 209:20]
  assign _T_22 = _T_16[1] & _T_20; // @[Misc.scala 213:38]
  assign _T_23 = _T_17 | _T_22; // @[Misc.scala 213:29]
  assign _T_25 = _T_16[1] & auto_mem_in_ar_bits_addr[1]; // @[Misc.scala 213:38]
  assign _T_26 = _T_17 | _T_25; // @[Misc.scala 213:29]
  assign _T_29 = ~auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 209:20]
  assign _T_30 = _T_20 & _T_29; // @[Misc.scala 212:27]
  assign _T_31 = _T_16[0] & _T_30; // @[Misc.scala 213:38]
  assign _T_32 = _T_23 | _T_31; // @[Misc.scala 213:29]
  assign _T_33 = _T_20 & auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  assign _T_34 = _T_16[0] & _T_33; // @[Misc.scala 213:38]
  assign _T_35 = _T_23 | _T_34; // @[Misc.scala 213:29]
  assign _T_36 = auto_mem_in_ar_bits_addr[1] & _T_29; // @[Misc.scala 212:27]
  assign _T_37 = _T_16[0] & _T_36; // @[Misc.scala 213:38]
  assign _T_38 = _T_26 | _T_37; // @[Misc.scala 213:29]
  assign _T_39 = auto_mem_in_ar_bits_addr[1] & auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  assign _T_40 = _T_16[0] & _T_39; // @[Misc.scala 213:38]
  assign _T_41 = _T_26 | _T_40; // @[Misc.scala 213:29]
  assign _T_44 = {_T_41,_T_38,_T_35,_T_32}; // @[Cat.scala 29:58]
  assign _T_46 = auto_mem_in_ar_valid ? _T_44 : auto_mem_in_w_bits_strb; // @[RegisterRouter.scala 54:25]
  assign _T_65 = _T_46[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_67 = _T_46[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_69 = _T_46[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_71 = _T_46[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_74 = {_T_71,_T_69,_T_67,_T_65}; // @[Cat.scala 29:58]
  assign _T_93 = _T_74[16:0] == 17'h1ffff; // @[RegisterRouter.scala 59:16]
  assign _T_146 = _T_3 & _T_47_ready; // @[RegisterRouter.scala 59:16]
  assign _T_140 = 2'h1 << _T_11[2]; // @[OneHot.scala 58:35]
  assign _T_163 = _T_146 & _T_4; // @[RegisterRouter.scala 59:16]
  assign _T_170 = _T_163 & _T_140[1]; // @[RegisterRouter.scala 59:16]
  assign _T_171 = _T_170 & _T_53; // @[RegisterRouter.scala 59:16]
  assign _T_100 = _T_171 & _T_93; // @[RegisterRouter.scala 59:16]
  assign _T_116 = _T_74[6:0] == 7'h7f; // @[RegisterRouter.scala 59:16]
  assign _T_165 = _T_163 & _T_140[0]; // @[RegisterRouter.scala 59:16]
  assign _T_166 = _T_165 & _T_53; // @[RegisterRouter.scala 59:16]
  assign _T_123 = _T_166 & _T_116; // @[RegisterRouter.scala 59:16]
  assign _GEN_11 = _T_11[2] ? _T_53 : _T_53; // @[MuxLiteral.scala 48:10]
  assign _T_218_0 = {{10'd0}, accDepth}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  assign _GEN_13 = _T_11[2] ? numWin : _T_218_0; // @[MuxLiteral.scala 48:10]
  assign _T_220 = _GEN_11 ? _GEN_13 : 17'h0; // @[RegisterRouter.scala 59:16]
  assign _T_221_bits_read = Queue_io_deq_bits_read; // @[Decoupled.scala 308:19 Decoupled.scala 309:14]
  assign _T_221_valid = Queue_io_deq_valid; // @[Decoupled.scala 308:19 Decoupled.scala 310:15]
  assign _T_224 = ~_T_221_bits_read; // @[RegisterRouter.scala 65:29]
  assign _T_228 = auto_slave_in_bits_data; // @[AccDspBlock.scala 63:48]
  assign auto_mem_in_aw_ready = _T_5 & auto_mem_in_w_valid; // @[LazyModule.scala 173:31]
  assign auto_mem_in_w_ready = _T_5 & auto_mem_in_aw_valid; // @[LazyModule.scala 173:31]
  assign auto_mem_in_b_valid = _T_221_valid & _T_224; // @[LazyModule.scala 173:31]
  assign auto_mem_in_b_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_mem_in_ar_ready = Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_valid = _T_221_valid & _T_221_bits_read; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 173:31]
  assign auto_master_out_valid = acc_io_out_valid; // @[LazyModule.scala 173:49]
  assign auto_master_out_bits_data = acc_io_out_bits; // @[LazyModule.scala 173:49]
  assign auto_master_out_bits_last = acc_io_lastOut; // @[LazyModule.scala 173:49]
  assign auto_slave_in_ready = acc_io_in_ready; // @[LazyModule.scala 173:31]
  assign acc_clock = clock;
  assign acc_reset = reset;
  assign acc_io_in_valid = auto_slave_in_valid; // @[AccDspBlock.scala 61:24]
  assign acc_io_in_bits = _T_228[15:0]; // @[AccDspBlock.scala 63:24]
  assign acc_io_lastIn = auto_slave_in_bits_last; // @[AccDspBlock.scala 66:24]
  assign acc_io_accDepthReg = accDepth; // @[AccDspBlock.scala 45:26]
  assign acc_io_accWindowsReg = numWin; // @[AccDspBlock.scala 46:26]
  assign acc_io_out_ready = auto_master_out_ready; // @[AccDspBlock.scala 70:22]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_mem_in_ar_valid | _T_2; // @[Decoupled.scala 288:22]
  assign Queue_io_enq_bits_read = auto_mem_in_ar_valid; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_data = {{15'd0}, _T_220}; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_extra = auto_mem_in_ar_valid ? auto_mem_in_ar_bits_id : auto_mem_in_aw_bits_id; // @[Decoupled.scala 289:21]
  assign Queue_io_deq_ready = _T_221_bits_read ? auto_mem_in_r_ready : auto_mem_in_b_ready; // @[Decoupled.scala 311:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  accDepth = _RAND_0[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  numWin = _RAND_1[16:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      accDepth <= 7'h40;
    end else if (_T_123) begin
      accDepth <= auto_mem_in_w_bits_data[6:0];
    end
    if (reset) begin
      numWin <= 17'h10000;
    end else if (_T_100) begin
      numWin <= auto_mem_in_w_bits_data[16:0];
    end
  end
endmodule
module Queue_22(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [15:0] io_enq_bits_data,
  input         io_enq_bits_last,
  input         io_deq_ready,
  output        io_deq_valid,
  output [15:0] io_deq_bits_data,
  output        io_deq_bits_last
);
  reg [15:0] _T_data [0:63]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_0;
  wire [15:0] _T_data__T_18_data; // @[Decoupled.scala 209:24]
  wire [5:0] _T_data__T_18_addr; // @[Decoupled.scala 209:24]
  wire [15:0] _T_data__T_10_data; // @[Decoupled.scala 209:24]
  wire [5:0] _T_data__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T_data__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T_data__T_10_en; // @[Decoupled.scala 209:24]
  reg  _T_last [0:63]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_1;
  wire  _T_last__T_18_data; // @[Decoupled.scala 209:24]
  wire [5:0] _T_last__T_18_addr; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_data; // @[Decoupled.scala 209:24]
  wire [5:0] _T_last__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_en; // @[Decoupled.scala 209:24]
  reg [5:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_2;
  reg [5:0] value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_3;
  reg  _T_1; // @[Decoupled.scala 212:35]
  reg [31:0] _RAND_4;
  wire  _T_2; // @[Decoupled.scala 214:41]
  wire  _T_3; // @[Decoupled.scala 215:36]
  wire  _T_4; // @[Decoupled.scala 215:33]
  wire  _T_5; // @[Decoupled.scala 216:32]
  wire  _T_6; // @[Decoupled.scala 40:37]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire [5:0] _T_12; // @[Counter.scala 39:22]
  wire [5:0] _T_14; // @[Counter.scala 39:22]
  wire  _T_15; // @[Decoupled.scala 227:16]
  assign _T_data__T_18_addr = value_1;
  assign _T_data__T_18_data = _T_data[_T_data__T_18_addr]; // @[Decoupled.scala 209:24]
  assign _T_data__T_10_data = io_enq_bits_data;
  assign _T_data__T_10_addr = value;
  assign _T_data__T_10_mask = 1'h1;
  assign _T_data__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_last__T_18_addr = value_1;
  assign _T_last__T_18_data = _T_last[_T_last__T_18_addr]; // @[Decoupled.scala 209:24]
  assign _T_last__T_10_data = io_enq_bits_last;
  assign _T_last__T_10_addr = value;
  assign _T_last__T_10_mask = 1'h1;
  assign _T_last__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_2 = value == value_1; // @[Decoupled.scala 214:41]
  assign _T_3 = ~_T_1; // @[Decoupled.scala 215:36]
  assign _T_4 = _T_2 & _T_3; // @[Decoupled.scala 215:33]
  assign _T_5 = _T_2 & _T_1; // @[Decoupled.scala 216:32]
  assign _T_6 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  assign _T_8 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  assign _T_12 = value + 6'h1; // @[Counter.scala 39:22]
  assign _T_14 = value_1 + 6'h1; // @[Counter.scala 39:22]
  assign _T_15 = _T_6 != _T_8; // @[Decoupled.scala 227:16]
  assign io_enq_ready = ~_T_5; // @[Decoupled.scala 232:16]
  assign io_deq_valid = ~_T_4; // @[Decoupled.scala 231:16]
  assign io_deq_bits_data = _T_data__T_18_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_last = _T_last__T_18_data; // @[Decoupled.scala 233:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    _T_data[initvar] = _RAND_0[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    _T_last[initvar] = _RAND_1[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  value = _RAND_2[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  value_1 = _RAND_3[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T_data__T_10_en & _T_data__T_10_mask) begin
      _T_data[_T_data__T_10_addr] <= _T_data__T_10_data; // @[Decoupled.scala 209:24]
    end
    if(_T_last__T_10_en & _T_last__T_10_mask) begin
      _T_last[_T_last__T_10_addr] <= _T_last__T_10_data; // @[Decoupled.scala 209:24]
    end
    if (reset) begin
      value <= 6'h0;
    end else if (_T_6) begin
      value <= _T_12;
    end
    if (reset) begin
      value_1 <= 6'h0;
    end else if (_T_8) begin
      value_1 <= _T_14;
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else if (_T_15) begin
      _T_1 <= _T_6;
    end
  end
endmodule
module Queue_23(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input         io_enq_bits_read,
  input  [9:0]  io_enq_bits_index,
  input  [31:0] io_enq_bits_data,
  input  [3:0]  io_enq_bits_mask,
  input         io_enq_bits_extra,
  input         io_deq_ready,
  output        io_deq_valid,
  output        io_deq_bits_read,
  output [9:0]  io_deq_bits_index,
  output [31:0] io_deq_bits_data,
  output [3:0]  io_deq_bits_mask,
  output        io_deq_bits_extra
);
  reg  _T_read [0:3]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_0;
  wire  _T_read__T_18_data; // @[Decoupled.scala 209:24]
  wire [1:0] _T_read__T_18_addr; // @[Decoupled.scala 209:24]
  wire  _T_read__T_10_data; // @[Decoupled.scala 209:24]
  wire [1:0] _T_read__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T_read__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T_read__T_10_en; // @[Decoupled.scala 209:24]
  reg [9:0] _T_index [0:3]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_1;
  wire [9:0] _T_index__T_18_data; // @[Decoupled.scala 209:24]
  wire [1:0] _T_index__T_18_addr; // @[Decoupled.scala 209:24]
  wire [9:0] _T_index__T_10_data; // @[Decoupled.scala 209:24]
  wire [1:0] _T_index__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T_index__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T_index__T_10_en; // @[Decoupled.scala 209:24]
  reg [31:0] _T_data [0:3]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_2;
  wire [31:0] _T_data__T_18_data; // @[Decoupled.scala 209:24]
  wire [1:0] _T_data__T_18_addr; // @[Decoupled.scala 209:24]
  wire [31:0] _T_data__T_10_data; // @[Decoupled.scala 209:24]
  wire [1:0] _T_data__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T_data__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T_data__T_10_en; // @[Decoupled.scala 209:24]
  reg [3:0] _T_mask [0:3]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_3;
  wire [3:0] _T_mask__T_18_data; // @[Decoupled.scala 209:24]
  wire [1:0] _T_mask__T_18_addr; // @[Decoupled.scala 209:24]
  wire [3:0] _T_mask__T_10_data; // @[Decoupled.scala 209:24]
  wire [1:0] _T_mask__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T_mask__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T_mask__T_10_en; // @[Decoupled.scala 209:24]
  reg  _T_extra [0:3]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_4;
  wire  _T_extra__T_18_data; // @[Decoupled.scala 209:24]
  wire [1:0] _T_extra__T_18_addr; // @[Decoupled.scala 209:24]
  wire  _T_extra__T_10_data; // @[Decoupled.scala 209:24]
  wire [1:0] _T_extra__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T_extra__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T_extra__T_10_en; // @[Decoupled.scala 209:24]
  reg [1:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  reg [1:0] value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_6;
  reg  _T_1; // @[Decoupled.scala 212:35]
  reg [31:0] _RAND_7;
  wire  _T_2; // @[Decoupled.scala 214:41]
  wire  _T_3; // @[Decoupled.scala 215:36]
  wire  _T_4; // @[Decoupled.scala 215:33]
  wire  _T_5; // @[Decoupled.scala 216:32]
  wire  _T_6; // @[Decoupled.scala 40:37]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire [1:0] _T_12; // @[Counter.scala 39:22]
  wire [1:0] _T_14; // @[Counter.scala 39:22]
  wire  _T_15; // @[Decoupled.scala 227:16]
  assign _T_read__T_18_addr = value_1;
  assign _T_read__T_18_data = _T_read[_T_read__T_18_addr]; // @[Decoupled.scala 209:24]
  assign _T_read__T_10_data = io_enq_bits_read;
  assign _T_read__T_10_addr = value;
  assign _T_read__T_10_mask = 1'h1;
  assign _T_read__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_index__T_18_addr = value_1;
  assign _T_index__T_18_data = _T_index[_T_index__T_18_addr]; // @[Decoupled.scala 209:24]
  assign _T_index__T_10_data = io_enq_bits_index;
  assign _T_index__T_10_addr = value;
  assign _T_index__T_10_mask = 1'h1;
  assign _T_index__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_data__T_18_addr = value_1;
  assign _T_data__T_18_data = _T_data[_T_data__T_18_addr]; // @[Decoupled.scala 209:24]
  assign _T_data__T_10_data = io_enq_bits_data;
  assign _T_data__T_10_addr = value;
  assign _T_data__T_10_mask = 1'h1;
  assign _T_data__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_mask__T_18_addr = value_1;
  assign _T_mask__T_18_data = _T_mask[_T_mask__T_18_addr]; // @[Decoupled.scala 209:24]
  assign _T_mask__T_10_data = io_enq_bits_mask;
  assign _T_mask__T_10_addr = value;
  assign _T_mask__T_10_mask = 1'h1;
  assign _T_mask__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_extra__T_18_addr = value_1;
  assign _T_extra__T_18_data = _T_extra[_T_extra__T_18_addr]; // @[Decoupled.scala 209:24]
  assign _T_extra__T_10_data = io_enq_bits_extra;
  assign _T_extra__T_10_addr = value;
  assign _T_extra__T_10_mask = 1'h1;
  assign _T_extra__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_2 = value == value_1; // @[Decoupled.scala 214:41]
  assign _T_3 = ~_T_1; // @[Decoupled.scala 215:36]
  assign _T_4 = _T_2 & _T_3; // @[Decoupled.scala 215:33]
  assign _T_5 = _T_2 & _T_1; // @[Decoupled.scala 216:32]
  assign _T_6 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  assign _T_8 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  assign _T_12 = value + 2'h1; // @[Counter.scala 39:22]
  assign _T_14 = value_1 + 2'h1; // @[Counter.scala 39:22]
  assign _T_15 = _T_6 != _T_8; // @[Decoupled.scala 227:16]
  assign io_enq_ready = ~_T_5; // @[Decoupled.scala 232:16]
  assign io_deq_valid = ~_T_4; // @[Decoupled.scala 231:16]
  assign io_deq_bits_read = _T_read__T_18_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_index = _T_index__T_18_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_data = _T_data__T_18_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_mask = _T_mask__T_18_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_extra = _T_extra__T_18_data; // @[Decoupled.scala 233:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    _T_read[initvar] = _RAND_0[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    _T_index[initvar] = _RAND_1[9:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    _T_data[initvar] = _RAND_2[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    _T_mask[initvar] = _RAND_3[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_4 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    _T_extra[initvar] = _RAND_4[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  value_1 = _RAND_6[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_1 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T_read__T_10_en & _T_read__T_10_mask) begin
      _T_read[_T_read__T_10_addr] <= _T_read__T_10_data; // @[Decoupled.scala 209:24]
    end
    if(_T_index__T_10_en & _T_index__T_10_mask) begin
      _T_index[_T_index__T_10_addr] <= _T_index__T_10_data; // @[Decoupled.scala 209:24]
    end
    if(_T_data__T_10_en & _T_data__T_10_mask) begin
      _T_data[_T_data__T_10_addr] <= _T_data__T_10_data; // @[Decoupled.scala 209:24]
    end
    if(_T_mask__T_10_en & _T_mask__T_10_mask) begin
      _T_mask[_T_mask__T_10_addr] <= _T_mask__T_10_data; // @[Decoupled.scala 209:24]
    end
    if(_T_extra__T_10_en & _T_extra__T_10_mask) begin
      _T_extra[_T_extra__T_10_addr] <= _T_extra__T_10_data; // @[Decoupled.scala 209:24]
    end
    if (reset) begin
      value <= 2'h0;
    end else if (_T_6) begin
      value <= _T_12;
    end
    if (reset) begin
      value_1 <= 2'h0;
    end else if (_T_8) begin
      value_1 <= _T_14;
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else if (_T_15) begin
      _T_1 <= _T_6;
    end
  end
endmodule
module AXI4DspQueueBlock(
  input         clock,
  input         reset,
  output        auto_stream_in_ready,
  input         auto_stream_in_valid,
  input  [15:0] auto_stream_in_bits_data,
  input         auto_stream_in_bits_last,
  input         auto_stream_out_ready,
  output        auto_stream_out_valid,
  output [15:0] auto_stream_out_bits_data,
  output        auto_stream_out_bits_last,
  output        auto_in_aw_ready,
  input         auto_in_aw_valid,
  input         auto_in_aw_bits_id,
  input  [29:0] auto_in_aw_bits_addr,
  output        auto_in_w_ready,
  input         auto_in_w_valid,
  input  [31:0] auto_in_w_bits_data,
  input  [3:0]  auto_in_w_bits_strb,
  input         auto_in_b_ready,
  output        auto_in_b_valid,
  output        auto_in_b_bits_id,
  output        auto_in_ar_ready,
  input         auto_in_ar_valid,
  input         auto_in_ar_bits_id,
  input  [29:0] auto_in_ar_bits_addr,
  input  [2:0]  auto_in_ar_bits_size,
  input         auto_in_r_ready,
  output        auto_in_r_valid,
  output        auto_in_r_bits_id,
  output [31:0] auto_in_r_bits_data
);
  wire  queuedStream_clock; // @[Decoupled.scala 287:21]
  wire  queuedStream_reset; // @[Decoupled.scala 287:21]
  wire  queuedStream_io_enq_ready; // @[Decoupled.scala 287:21]
  wire  queuedStream_io_enq_valid; // @[Decoupled.scala 287:21]
  wire [15:0] queuedStream_io_enq_bits_data; // @[Decoupled.scala 287:21]
  wire  queuedStream_io_enq_bits_last; // @[Decoupled.scala 287:21]
  wire  queuedStream_io_deq_ready; // @[Decoupled.scala 287:21]
  wire  queuedStream_io_deq_valid; // @[Decoupled.scala 287:21]
  wire [15:0] queuedStream_io_deq_bits_data; // @[Decoupled.scala 287:21]
  wire  queuedStream_io_deq_bits_last; // @[Decoupled.scala 287:21]
  wire  Queue_clock; // @[Decoupled.scala 287:21]
  wire  Queue_reset; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_read; // @[Decoupled.scala 287:21]
  wire [9:0] Queue_io_enq_bits_index; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_enq_bits_data; // @[Decoupled.scala 287:21]
  wire [3:0] Queue_io_enq_bits_mask; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_extra; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_read; // @[Decoupled.scala 287:21]
  wire [9:0] Queue_io_deq_bits_index; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_deq_bits_data; // @[Decoupled.scala 287:21]
  wire [3:0] Queue_io_deq_bits_mask; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_extra; // @[Decoupled.scala 287:21]
  wire  Queue_1_clock; // @[Decoupled.scala 287:21]
  wire  Queue_1_reset; // @[Decoupled.scala 287:21]
  wire  Queue_1_io_enq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_1_io_enq_valid; // @[Decoupled.scala 287:21]
  wire  Queue_1_io_enq_bits_read; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_1_io_enq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_1_io_enq_bits_extra; // @[Decoupled.scala 287:21]
  wire  Queue_1_io_deq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_1_io_deq_valid; // @[Decoupled.scala 287:21]
  wire  Queue_1_io_deq_bits_read; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_1_io_deq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_1_io_deq_bits_extra; // @[Decoupled.scala 287:21]
  wire  _T_53_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 290:17]
  wire  _T_154; // @[RegisterRouter.scala 59:16]
  wire  _T_155; // @[RegisterRouter.scala 59:16]
  wire  _T_156; // @[RegisterRouter.scala 59:16]
  wire [9:0] _T_57; // @[RegisterRouter.scala 59:16]
  wire  _T_59; // @[RegisterRouter.scala 59:16]
  wire  _T_159; // @[RegisterRouter.scala 59:16]
  wire [7:0] _T_90; // @[Bitwise.scala 72:12]
  wire [7:0] _T_88; // @[Bitwise.scala 72:12]
  wire [7:0] _T_86; // @[Bitwise.scala 72:12]
  wire [7:0] _T_84; // @[Bitwise.scala 72:12]
  wire [31:0] _T_93; // @[Cat.scala 29:58]
  wire  _T_101; // @[RegisterRouter.scala 59:16]
  wire  _T_105; // @[RegisterRouter.scala 59:16]
  wire [31:0] _T_106; // @[RegisterRouter.scala 59:16]
  wire [31:0] queueThreshold; // @[RegField.scala 134:88]
  wire  _T_8; // @[RegisterRouter.scala 40:39]
  wire  _T_10; // @[RegisterRouter.scala 42:29]
  wire  _T_54_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 290:17]
  wire [29:0] _T_17; // @[RegisterRouter.scala 48:19]
  wire  _T_11; // @[RegisterRouter.scala 42:26]
  wire [1:0] _T_20; // @[OneHot.scala 65:12]
  wire [1:0] _T_22; // @[Misc.scala 200:81]
  wire  _T_23; // @[Misc.scala 204:21]
  wire  _T_26; // @[Misc.scala 209:20]
  wire  _T_28; // @[Misc.scala 213:38]
  wire  _T_29; // @[Misc.scala 213:29]
  wire  _T_31; // @[Misc.scala 213:38]
  wire  _T_32; // @[Misc.scala 213:29]
  wire  _T_35; // @[Misc.scala 209:20]
  wire  _T_36; // @[Misc.scala 212:27]
  wire  _T_37; // @[Misc.scala 213:38]
  wire  _T_38; // @[Misc.scala 213:29]
  wire  _T_39; // @[Misc.scala 212:27]
  wire  _T_40; // @[Misc.scala 213:38]
  wire  _T_41; // @[Misc.scala 213:29]
  wire  _T_42; // @[Misc.scala 212:27]
  wire  _T_43; // @[Misc.scala 213:38]
  wire  _T_44; // @[Misc.scala 213:29]
  wire  _T_45; // @[Misc.scala 212:27]
  wire  _T_46; // @[Misc.scala 213:38]
  wire  _T_47; // @[Misc.scala 213:29]
  wire [3:0] _T_50; // @[Cat.scala 29:58]
  wire  _T_178_bits_read; // @[Decoupled.scala 308:19 Decoupled.scala 309:14]
  wire  _T_178_valid; // @[Decoupled.scala 308:19 Decoupled.scala 310:15]
  wire  _T_181; // @[RegisterRouter.scala 65:29]
  Queue_22 queuedStream ( // @[Decoupled.scala 287:21]
    .clock(queuedStream_clock),
    .reset(queuedStream_reset),
    .io_enq_ready(queuedStream_io_enq_ready),
    .io_enq_valid(queuedStream_io_enq_valid),
    .io_enq_bits_data(queuedStream_io_enq_bits_data),
    .io_enq_bits_last(queuedStream_io_enq_bits_last),
    .io_deq_ready(queuedStream_io_deq_ready),
    .io_deq_valid(queuedStream_io_deq_valid),
    .io_deq_bits_data(queuedStream_io_deq_bits_data),
    .io_deq_bits_last(queuedStream_io_deq_bits_last)
  );
  Queue_23 Queue ( // @[Decoupled.scala 287:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_read(Queue_io_enq_bits_read),
    .io_enq_bits_index(Queue_io_enq_bits_index),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_mask(Queue_io_enq_bits_mask),
    .io_enq_bits_extra(Queue_io_enq_bits_extra),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_read(Queue_io_deq_bits_read),
    .io_deq_bits_index(Queue_io_deq_bits_index),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_mask(Queue_io_deq_bits_mask),
    .io_deq_bits_extra(Queue_io_deq_bits_extra)
  );
  Queue Queue_1 ( // @[Decoupled.scala 287:21]
    .clock(Queue_1_clock),
    .reset(Queue_1_reset),
    .io_enq_ready(Queue_1_io_enq_ready),
    .io_enq_valid(Queue_1_io_enq_valid),
    .io_enq_bits_read(Queue_1_io_enq_bits_read),
    .io_enq_bits_data(Queue_1_io_enq_bits_data),
    .io_enq_bits_extra(Queue_1_io_enq_bits_extra),
    .io_deq_ready(Queue_1_io_deq_ready),
    .io_deq_valid(Queue_1_io_deq_valid),
    .io_deq_bits_read(Queue_1_io_deq_bits_read),
    .io_deq_bits_data(Queue_1_io_deq_bits_data),
    .io_deq_bits_extra(Queue_1_io_deq_bits_extra)
  );
  assign _T_53_ready = Queue_1_io_enq_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 290:17]
  assign _T_154 = Queue_io_deq_valid & _T_53_ready; // @[RegisterRouter.scala 59:16]
  assign _T_155 = ~Queue_io_deq_bits_read; // @[RegisterRouter.scala 59:16]
  assign _T_156 = _T_154 & _T_155; // @[RegisterRouter.scala 59:16]
  assign _T_57 = Queue_io_deq_bits_index; // @[RegisterRouter.scala 59:16]
  assign _T_59 = _T_57 == 10'h0; // @[RegisterRouter.scala 59:16]
  assign _T_159 = _T_156 & _T_59; // @[RegisterRouter.scala 59:16]
  assign _T_90 = Queue_io_deq_bits_mask[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_88 = Queue_io_deq_bits_mask[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_86 = Queue_io_deq_bits_mask[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_84 = Queue_io_deq_bits_mask[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_93 = {_T_90,_T_88,_T_86,_T_84}; // @[Cat.scala 29:58]
  assign _T_101 = _T_93 == 32'hffffffff; // @[RegisterRouter.scala 59:16]
  assign _T_105 = _T_159 & _T_101; // @[RegisterRouter.scala 59:16]
  assign _T_106 = Queue_io_deq_bits_data; // @[RegisterRouter.scala 59:16]
  assign queueThreshold = _T_105 ? _T_106 : 32'h40; // @[RegField.scala 134:88]
  assign _T_8 = auto_in_aw_valid & auto_in_w_valid; // @[RegisterRouter.scala 40:39]
  assign _T_10 = ~auto_in_ar_valid; // @[RegisterRouter.scala 42:29]
  assign _T_54_ready = Queue_io_enq_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 290:17]
  assign _T_17 = auto_in_ar_valid ? auto_in_ar_bits_addr : auto_in_aw_bits_addr; // @[RegisterRouter.scala 48:19]
  assign _T_11 = _T_54_ready & _T_10; // @[RegisterRouter.scala 42:26]
  assign _T_20 = 2'h1 << auto_in_ar_bits_size[0]; // @[OneHot.scala 65:12]
  assign _T_22 = _T_20 | 2'h1; // @[Misc.scala 200:81]
  assign _T_23 = auto_in_ar_bits_size >= 3'h2; // @[Misc.scala 204:21]
  assign _T_26 = ~auto_in_ar_bits_addr[1]; // @[Misc.scala 209:20]
  assign _T_28 = _T_22[1] & _T_26; // @[Misc.scala 213:38]
  assign _T_29 = _T_23 | _T_28; // @[Misc.scala 213:29]
  assign _T_31 = _T_22[1] & auto_in_ar_bits_addr[1]; // @[Misc.scala 213:38]
  assign _T_32 = _T_23 | _T_31; // @[Misc.scala 213:29]
  assign _T_35 = ~auto_in_ar_bits_addr[0]; // @[Misc.scala 209:20]
  assign _T_36 = _T_26 & _T_35; // @[Misc.scala 212:27]
  assign _T_37 = _T_22[0] & _T_36; // @[Misc.scala 213:38]
  assign _T_38 = _T_29 | _T_37; // @[Misc.scala 213:29]
  assign _T_39 = _T_26 & auto_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  assign _T_40 = _T_22[0] & _T_39; // @[Misc.scala 213:38]
  assign _T_41 = _T_29 | _T_40; // @[Misc.scala 213:29]
  assign _T_42 = auto_in_ar_bits_addr[1] & _T_35; // @[Misc.scala 212:27]
  assign _T_43 = _T_22[0] & _T_42; // @[Misc.scala 213:38]
  assign _T_44 = _T_32 | _T_43; // @[Misc.scala 213:29]
  assign _T_45 = auto_in_ar_bits_addr[1] & auto_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  assign _T_46 = _T_22[0] & _T_45; // @[Misc.scala 213:38]
  assign _T_47 = _T_32 | _T_46; // @[Misc.scala 213:29]
  assign _T_50 = {_T_47,_T_44,_T_41,_T_38}; // @[Cat.scala 29:58]
  assign _T_178_bits_read = Queue_1_io_deq_bits_read; // @[Decoupled.scala 308:19 Decoupled.scala 309:14]
  assign _T_178_valid = Queue_1_io_deq_valid; // @[Decoupled.scala 308:19 Decoupled.scala 310:15]
  assign _T_181 = ~_T_178_bits_read; // @[RegisterRouter.scala 65:29]
  assign auto_stream_in_ready = queuedStream_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_stream_out_valid = queuedStream_io_deq_valid; // @[LazyModule.scala 173:49]
  assign auto_stream_out_bits_data = queuedStream_io_deq_bits_data; // @[LazyModule.scala 173:49]
  assign auto_stream_out_bits_last = queuedStream_io_deq_bits_last; // @[LazyModule.scala 173:49]
  assign auto_in_aw_ready = _T_11 & auto_in_w_valid; // @[LazyModule.scala 173:31]
  assign auto_in_w_ready = _T_11 & auto_in_aw_valid; // @[LazyModule.scala 173:31]
  assign auto_in_b_valid = _T_178_valid & _T_181; // @[LazyModule.scala 173:31]
  assign auto_in_b_bits_id = Queue_1_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_in_ar_ready = Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_in_r_valid = _T_178_valid & _T_178_bits_read; // @[LazyModule.scala 173:31]
  assign auto_in_r_bits_id = Queue_1_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_in_r_bits_data = Queue_1_io_deq_bits_data; // @[LazyModule.scala 173:31]
  assign queuedStream_clock = clock;
  assign queuedStream_reset = reset;
  assign queuedStream_io_enq_valid = auto_stream_in_valid; // @[Decoupled.scala 288:22]
  assign queuedStream_io_enq_bits_data = auto_stream_in_bits_data; // @[Decoupled.scala 289:21]
  assign queuedStream_io_enq_bits_last = auto_stream_in_bits_last; // @[Decoupled.scala 289:21]
  assign queuedStream_io_deq_ready = auto_stream_out_ready; // @[DspQueueBlock.scala 25:13]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_in_ar_valid | _T_8; // @[Decoupled.scala 288:22]
  assign Queue_io_enq_bits_read = auto_in_ar_valid; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_index = _T_17[11:2]; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_data = auto_in_w_bits_data; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_mask = auto_in_ar_valid ? _T_50 : auto_in_w_bits_strb; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_extra = auto_in_ar_valid ? auto_in_ar_bits_id : auto_in_aw_bits_id; // @[Decoupled.scala 289:21]
  assign Queue_io_deq_ready = Queue_1_io_enq_ready; // @[RegisterRouter.scala 59:16]
  assign Queue_1_clock = clock;
  assign Queue_1_reset = reset;
  assign Queue_1_io_enq_valid = Queue_io_deq_valid; // @[Decoupled.scala 288:22]
  assign Queue_1_io_enq_bits_read = Queue_io_deq_bits_read; // @[Decoupled.scala 289:21]
  assign Queue_1_io_enq_bits_data = _T_59 ? queueThreshold : 32'h0; // @[Decoupled.scala 289:21]
  assign Queue_1_io_enq_bits_extra = Queue_io_deq_bits_extra; // @[Decoupled.scala 289:21]
  assign Queue_1_io_deq_ready = _T_178_bits_read ? auto_in_r_ready : auto_in_b_ready; // @[Decoupled.scala 311:15]
endmodule
module AXI4Xbar_1(
  input         clock,
  input         reset,
  output        auto_in_aw_ready,
  input         auto_in_aw_valid,
  input         auto_in_aw_bits_id,
  input  [29:0] auto_in_aw_bits_addr,
  input  [2:0]  auto_in_aw_bits_size,
  output        auto_in_w_ready,
  input         auto_in_w_valid,
  input  [31:0] auto_in_w_bits_data,
  input  [3:0]  auto_in_w_bits_strb,
  input         auto_in_w_bits_last,
  input         auto_in_b_ready,
  output        auto_in_b_valid,
  output [1:0]  auto_in_b_bits_resp,
  output        auto_in_ar_ready,
  input         auto_in_ar_valid,
  input         auto_in_ar_bits_id,
  input  [29:0] auto_in_ar_bits_addr,
  input  [2:0]  auto_in_ar_bits_size,
  input         auto_in_r_ready,
  output        auto_in_r_valid,
  output [31:0] auto_in_r_bits_data,
  output [1:0]  auto_in_r_bits_resp,
  output        auto_in_r_bits_last,
  input         auto_out_1_aw_ready,
  output        auto_out_1_aw_valid,
  output        auto_out_1_aw_bits_id,
  output [29:0] auto_out_1_aw_bits_addr,
  output [2:0]  auto_out_1_aw_bits_size,
  input         auto_out_1_w_ready,
  output        auto_out_1_w_valid,
  output [31:0] auto_out_1_w_bits_data,
  output [3:0]  auto_out_1_w_bits_strb,
  output        auto_out_1_w_bits_last,
  output        auto_out_1_b_ready,
  input         auto_out_1_b_valid,
  input         auto_out_1_b_bits_id,
  input  [1:0]  auto_out_1_b_bits_resp,
  input         auto_out_1_ar_ready,
  output        auto_out_1_ar_valid,
  output        auto_out_1_ar_bits_id,
  output [29:0] auto_out_1_ar_bits_addr,
  output [2:0]  auto_out_1_ar_bits_size,
  output        auto_out_1_r_ready,
  input         auto_out_1_r_valid,
  input         auto_out_1_r_bits_id,
  input  [31:0] auto_out_1_r_bits_data,
  input  [1:0]  auto_out_1_r_bits_resp,
  input         auto_out_1_r_bits_last,
  input         auto_out_0_aw_ready,
  output        auto_out_0_aw_valid,
  output        auto_out_0_aw_bits_id,
  output [29:0] auto_out_0_aw_bits_addr,
  output [2:0]  auto_out_0_aw_bits_size,
  input         auto_out_0_w_ready,
  output        auto_out_0_w_valid,
  output [31:0] auto_out_0_w_bits_data,
  output [3:0]  auto_out_0_w_bits_strb,
  output        auto_out_0_w_bits_last,
  output        auto_out_0_b_ready,
  input         auto_out_0_b_valid,
  input         auto_out_0_b_bits_id,
  input  [1:0]  auto_out_0_b_bits_resp,
  input         auto_out_0_ar_ready,
  output        auto_out_0_ar_valid,
  output        auto_out_0_ar_bits_id,
  output [29:0] auto_out_0_ar_bits_addr,
  output [2:0]  auto_out_0_ar_bits_size,
  output        auto_out_0_r_ready,
  input         auto_out_0_r_valid,
  input         auto_out_0_r_bits_id,
  input  [31:0] auto_out_0_r_bits_data,
  input  [1:0]  auto_out_0_r_bits_resp,
  input         auto_out_0_r_bits_last
);
  wire  awIn_0_clock; // @[Xbar.scala 55:47]
  wire  awIn_0_reset; // @[Xbar.scala 55:47]
  wire  awIn_0_io_enq_ready; // @[Xbar.scala 55:47]
  wire  awIn_0_io_enq_valid; // @[Xbar.scala 55:47]
  wire [1:0] awIn_0_io_enq_bits; // @[Xbar.scala 55:47]
  wire  awIn_0_io_deq_ready; // @[Xbar.scala 55:47]
  wire  awIn_0_io_deq_valid; // @[Xbar.scala 55:47]
  wire [1:0] awIn_0_io_deq_bits; // @[Xbar.scala 55:47]
  wire [30:0] _T_1; // @[Parameters.scala 137:49]
  wire [30:0] _T_3; // @[Parameters.scala 137:52]
  wire  requestARIO_0_0; // @[Parameters.scala 137:67]
  wire [29:0] _T_5; // @[Parameters.scala 137:31]
  wire [30:0] _T_6; // @[Parameters.scala 137:49]
  wire [30:0] _T_8; // @[Parameters.scala 137:52]
  wire  requestARIO_0_1; // @[Parameters.scala 137:67]
  wire [30:0] _T_11; // @[Parameters.scala 137:49]
  wire [30:0] _T_13; // @[Parameters.scala 137:52]
  wire  requestAWIO_0_0; // @[Parameters.scala 137:67]
  wire [29:0] _T_15; // @[Parameters.scala 137:31]
  wire [30:0] _T_16; // @[Parameters.scala 137:49]
  wire [30:0] _T_18; // @[Parameters.scala 137:52]
  wire  requestAWIO_0_1; // @[Parameters.scala 137:67]
  wire  requestROI_0_0; // @[Parameters.scala 47:9]
  wire  requestROI_1_0; // @[Parameters.scala 47:9]
  wire  requestBOI_0_0; // @[Parameters.scala 47:9]
  wire  requestBOI_1_0; // @[Parameters.scala 47:9]
  wire [1:0] _T_20; // @[Xbar.scala 64:75]
  wire  requestWIO_0_0; // @[Xbar.scala 65:73]
  wire  requestWIO_0_1; // @[Xbar.scala 65:73]
  wire [1:0] _T_27; // @[Xbar.scala 93:45]
  wire  _T_108; // @[Mux.scala 27:72]
  wire  _T_109; // @[Mux.scala 27:72]
  wire  in_0_ar_ready; // @[Mux.scala 27:72]
  reg [2:0] _T_36; // @[Xbar.scala 104:34]
  reg [31:0] _RAND_0;
  wire  _T_55; // @[Xbar.scala 112:22]
  reg  _T_37; // @[Xbar.scala 105:29]
  reg [31:0] _RAND_1;
  wire  _T_54; // @[Xbar.scala 111:75]
  wire  _T_56; // @[Xbar.scala 112:34]
  wire  _T_57; // @[Xbar.scala 112:80]
  wire  _T_59; // @[Xbar.scala 112:48]
  wire  io_in_0_ar_ready; // @[Xbar.scala 130:45]
  wire  _T_31; // @[Decoupled.scala 40:37]
  reg  _T_222; // @[Xbar.scala 242:23]
  reg [31:0] _RAND_2;
  wire  _T_127; // @[Xbar.scala 222:40]
  wire  _T_129; // @[Xbar.scala 222:40]
  wire  _T_223; // @[Xbar.scala 246:36]
  reg  _T_278_0; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_3;
  wire  _T_284; // @[Mux.scala 27:72]
  reg  _T_278_1; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_4;
  wire  _T_285; // @[Mux.scala 27:72]
  wire  _T_286; // @[Mux.scala 27:72]
  wire  in_0_r_valid; // @[Xbar.scala 278:22]
  wire  _T_33; // @[Decoupled.scala 40:37]
  wire [1:0] _T_224; // @[Cat.scala 29:58]
  reg [1:0] _T_231; // @[Arbiter.scala 20:23]
  reg [31:0] _RAND_5;
  wire [1:0] _T_232; // @[Arbiter.scala 21:30]
  wire [1:0] _T_233; // @[Arbiter.scala 21:28]
  wire [3:0] _T_234; // @[Cat.scala 29:58]
  wire [3:0] _GEN_18; // @[package.scala 208:43]
  wire [3:0] _T_236; // @[package.scala 208:43]
  wire [3:0] _T_239; // @[Arbiter.scala 22:66]
  wire [3:0] _GEN_19; // @[Arbiter.scala 22:58]
  wire [3:0] _T_240; // @[Arbiter.scala 22:58]
  wire [1:0] _T_243; // @[Arbiter.scala 23:39]
  wire [1:0] _T_244; // @[Arbiter.scala 23:18]
  wire  _T_256; // @[Xbar.scala 250:63]
  wire  _T_279_0; // @[Xbar.scala 262:23]
  wire [35:0] _T_291; // @[Mux.scala 27:72]
  wire [35:0] _T_292; // @[Mux.scala 27:72]
  wire  _T_257; // @[Xbar.scala 250:63]
  wire  _T_279_1; // @[Xbar.scala 262:23]
  wire [35:0] _T_295; // @[Mux.scala 27:72]
  wire [35:0] _T_296; // @[Mux.scala 27:72]
  wire [35:0] _T_297; // @[Mux.scala 27:72]
  wire  in_0_r_bits_last; // @[Mux.scala 27:72]
  wire  _T_35; // @[Xbar.scala 120:45]
  wire [2:0] _GEN_20; // @[Xbar.scala 106:30]
  wire [2:0] _T_39; // @[Xbar.scala 106:30]
  wire [2:0] _GEN_21; // @[Xbar.scala 106:48]
  wire [2:0] _T_41; // @[Xbar.scala 106:48]
  wire  _T_42; // @[Xbar.scala 107:23]
  wire  _T_43; // @[Xbar.scala 107:43]
  wire  _T_44; // @[Xbar.scala 107:34]
  wire  _T_46; // @[Xbar.scala 107:22]
  wire  _T_47; // @[Xbar.scala 107:22]
  wire  _T_48; // @[Xbar.scala 108:23]
  wire  _T_50; // @[Xbar.scala 108:34]
  wire  _T_52; // @[Xbar.scala 108:22]
  wire  _T_53; // @[Xbar.scala 108:22]
  wire  _T_115; // @[Mux.scala 27:72]
  wire  _T_116; // @[Mux.scala 27:72]
  wire  in_0_aw_ready; // @[Mux.scala 27:72]
  reg  _T_90; // @[Xbar.scala 137:30]
  reg [31:0] _RAND_6;
  wire  _T_94; // @[Xbar.scala 139:57]
  wire  _T_95; // @[Xbar.scala 139:45]
  reg [2:0] _T_64; // @[Xbar.scala 104:34]
  reg [31:0] _RAND_7;
  wire  _T_83; // @[Xbar.scala 112:22]
  reg  _T_65; // @[Xbar.scala 105:29]
  reg [31:0] _RAND_8;
  wire  _T_82; // @[Xbar.scala 111:75]
  wire  _T_84; // @[Xbar.scala 112:34]
  wire  _T_85; // @[Xbar.scala 112:80]
  wire  _T_87; // @[Xbar.scala 112:48]
  wire  io_in_0_aw_ready; // @[Xbar.scala 139:82]
  wire  _T_60; // @[Decoupled.scala 40:37]
  reg  _T_304; // @[Xbar.scala 242:23]
  reg [31:0] _RAND_9;
  wire  _T_131; // @[Xbar.scala 222:40]
  wire  _T_133; // @[Xbar.scala 222:40]
  wire  _T_305; // @[Xbar.scala 246:36]
  reg  _T_360_0; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_10;
  wire  _T_366; // @[Mux.scala 27:72]
  reg  _T_360_1; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_11;
  wire  _T_367; // @[Mux.scala 27:72]
  wire  _T_368; // @[Mux.scala 27:72]
  wire  in_0_b_valid; // @[Xbar.scala 278:22]
  wire  _T_62; // @[Decoupled.scala 40:37]
  wire [2:0] _GEN_22; // @[Xbar.scala 106:30]
  wire [2:0] _T_67; // @[Xbar.scala 106:30]
  wire [2:0] _GEN_23; // @[Xbar.scala 106:48]
  wire [2:0] _T_69; // @[Xbar.scala 106:48]
  wire  _T_70; // @[Xbar.scala 107:23]
  wire  _T_71; // @[Xbar.scala 107:43]
  wire  _T_72; // @[Xbar.scala 107:34]
  wire  _T_74; // @[Xbar.scala 107:22]
  wire  _T_75; // @[Xbar.scala 107:22]
  wire  _T_76; // @[Xbar.scala 108:23]
  wire  _T_78; // @[Xbar.scala 108:34]
  wire  _T_80; // @[Xbar.scala 108:22]
  wire  _T_81; // @[Xbar.scala 108:22]
  wire  in_0_ar_valid; // @[Xbar.scala 129:45]
  wire  _T_92; // @[Xbar.scala 138:45]
  wire  in_0_aw_valid; // @[Xbar.scala 138:82]
  wire  _T_97; // @[Xbar.scala 140:54]
  wire  _T_99; // @[Decoupled.scala 40:37]
  wire  _GEN_2; // @[Xbar.scala 141:38]
  wire  _T_100; // @[Decoupled.scala 40:37]
  wire  in_0_w_valid; // @[Xbar.scala 145:43]
  wire  _T_122; // @[Mux.scala 27:72]
  wire  _T_123; // @[Mux.scala 27:72]
  wire  in_0_w_ready; // @[Mux.scala 27:72]
  wire  _T_103; // @[Xbar.scala 147:50]
  wire  out_0_ar_valid; // @[Xbar.scala 222:40]
  wire  out_1_ar_valid; // @[Xbar.scala 222:40]
  wire  out_0_aw_valid; // @[Xbar.scala 222:40]
  wire  out_1_aw_valid; // @[Xbar.scala 222:40]
  wire  _T_140; // @[Xbar.scala 256:60]
  wire  _T_146; // @[Xbar.scala 258:23]
  wire  _T_148; // @[Xbar.scala 258:12]
  wire  _T_149; // @[Xbar.scala 258:12]
  wire  _T_161; // @[Xbar.scala 256:60]
  wire  _T_167; // @[Xbar.scala 258:23]
  wire  _T_169; // @[Xbar.scala 258:12]
  wire  _T_170; // @[Xbar.scala 258:12]
  wire  _T_184; // @[Xbar.scala 256:60]
  wire  _T_190; // @[Xbar.scala 258:23]
  wire  _T_192; // @[Xbar.scala 258:12]
  wire  _T_193; // @[Xbar.scala 258:12]
  wire  _T_205; // @[Xbar.scala 256:60]
  wire  _T_211; // @[Xbar.scala 258:23]
  wire  _T_213; // @[Xbar.scala 258:12]
  wire  _T_214; // @[Xbar.scala 258:12]
  wire  _T_245; // @[Arbiter.scala 24:27]
  wire  _T_246; // @[Arbiter.scala 24:18]
  wire [1:0] _T_247; // @[Arbiter.scala 25:29]
  wire [2:0] _T_248; // @[package.scala 199:48]
  wire [1:0] _T_250; // @[package.scala 199:43]
  wire  _T_260; // @[Xbar.scala 255:50]
  wire  _T_262; // @[Xbar.scala 256:60]
  wire  _T_265; // @[Xbar.scala 256:60]
  wire  _T_266; // @[Xbar.scala 256:57]
  wire  _T_269; // @[Xbar.scala 256:11]
  wire  _T_270; // @[Xbar.scala 256:11]
  wire  _T_271; // @[Xbar.scala 258:13]
  wire  _T_273; // @[Xbar.scala 258:23]
  wire  _T_275; // @[Xbar.scala 258:12]
  wire  _T_276; // @[Xbar.scala 258:12]
  wire  _GEN_13; // @[Xbar.scala 266:21]
  wire  _GEN_14; // @[Xbar.scala 267:24]
  wire  _T_281_0; // @[Xbar.scala 270:24]
  wire  _T_281_1; // @[Xbar.scala 270:24]
  wire [1:0] _T_306; // @[Cat.scala 29:58]
  reg [1:0] _T_313; // @[Arbiter.scala 20:23]
  reg [31:0] _RAND_12;
  wire [1:0] _T_314; // @[Arbiter.scala 21:30]
  wire [1:0] _T_315; // @[Arbiter.scala 21:28]
  wire [3:0] _T_316; // @[Cat.scala 29:58]
  wire [3:0] _GEN_24; // @[package.scala 208:43]
  wire [3:0] _T_318; // @[package.scala 208:43]
  wire [3:0] _T_321; // @[Arbiter.scala 22:66]
  wire [3:0] _GEN_25; // @[Arbiter.scala 22:58]
  wire [3:0] _T_322; // @[Arbiter.scala 22:58]
  wire [1:0] _T_325; // @[Arbiter.scala 23:39]
  wire [1:0] _T_326; // @[Arbiter.scala 23:18]
  wire  _T_327; // @[Arbiter.scala 24:27]
  wire  _T_328; // @[Arbiter.scala 24:18]
  wire [1:0] _T_329; // @[Arbiter.scala 25:29]
  wire [2:0] _T_330; // @[package.scala 199:48]
  wire [1:0] _T_332; // @[package.scala 199:43]
  wire  _T_338; // @[Xbar.scala 250:63]
  wire  _T_339; // @[Xbar.scala 250:63]
  wire  _T_342; // @[Xbar.scala 255:50]
  wire  _T_344; // @[Xbar.scala 256:60]
  wire  _T_347; // @[Xbar.scala 256:60]
  wire  _T_348; // @[Xbar.scala 256:57]
  wire  _T_351; // @[Xbar.scala 256:11]
  wire  _T_352; // @[Xbar.scala 256:11]
  wire  _T_353; // @[Xbar.scala 258:13]
  wire  _T_355; // @[Xbar.scala 258:23]
  wire  _T_357; // @[Xbar.scala 258:12]
  wire  _T_358; // @[Xbar.scala 258:12]
  wire  _T_361_0; // @[Xbar.scala 262:23]
  wire  _T_361_1; // @[Xbar.scala 262:23]
  wire  _GEN_16; // @[Xbar.scala 266:21]
  wire  _GEN_17; // @[Xbar.scala 267:24]
  wire  _T_363_0; // @[Xbar.scala 270:24]
  wire  _T_363_1; // @[Xbar.scala 270:24]
  wire [2:0] _T_371; // @[Mux.scala 27:72]
  wire [2:0] _T_372; // @[Mux.scala 27:72]
  wire [2:0] _T_373; // @[Mux.scala 27:72]
  wire [2:0] _T_374; // @[Mux.scala 27:72]
  wire [2:0] _T_375; // @[Mux.scala 27:72]
  QueueCompatibility awIn_0 ( // @[Xbar.scala 55:47]
    .clock(awIn_0_clock),
    .reset(awIn_0_reset),
    .io_enq_ready(awIn_0_io_enq_ready),
    .io_enq_valid(awIn_0_io_enq_valid),
    .io_enq_bits(awIn_0_io_enq_bits),
    .io_deq_ready(awIn_0_io_deq_ready),
    .io_deq_valid(awIn_0_io_deq_valid),
    .io_deq_bits(awIn_0_io_deq_bits)
  );
  assign _T_1 = {1'b0,$signed(auto_in_ar_bits_addr)}; // @[Parameters.scala 137:49]
  assign _T_3 = $signed(_T_1) & 31'sh1000; // @[Parameters.scala 137:52]
  assign requestARIO_0_0 = $signed(_T_3) == 31'sh0; // @[Parameters.scala 137:67]
  assign _T_5 = auto_in_ar_bits_addr ^ 30'h1000; // @[Parameters.scala 137:31]
  assign _T_6 = {1'b0,$signed(_T_5)}; // @[Parameters.scala 137:49]
  assign _T_8 = $signed(_T_6) & 31'sh1000; // @[Parameters.scala 137:52]
  assign requestARIO_0_1 = $signed(_T_8) == 31'sh0; // @[Parameters.scala 137:67]
  assign _T_11 = {1'b0,$signed(auto_in_aw_bits_addr)}; // @[Parameters.scala 137:49]
  assign _T_13 = $signed(_T_11) & 31'sh1000; // @[Parameters.scala 137:52]
  assign requestAWIO_0_0 = $signed(_T_13) == 31'sh0; // @[Parameters.scala 137:67]
  assign _T_15 = auto_in_aw_bits_addr ^ 30'h1000; // @[Parameters.scala 137:31]
  assign _T_16 = {1'b0,$signed(_T_15)}; // @[Parameters.scala 137:49]
  assign _T_18 = $signed(_T_16) & 31'sh1000; // @[Parameters.scala 137:52]
  assign requestAWIO_0_1 = $signed(_T_18) == 31'sh0; // @[Parameters.scala 137:67]
  assign requestROI_0_0 = ~auto_out_0_r_bits_id; // @[Parameters.scala 47:9]
  assign requestROI_1_0 = ~auto_out_1_r_bits_id; // @[Parameters.scala 47:9]
  assign requestBOI_0_0 = ~auto_out_0_b_bits_id; // @[Parameters.scala 47:9]
  assign requestBOI_1_0 = ~auto_out_1_b_bits_id; // @[Parameters.scala 47:9]
  assign _T_20 = {requestAWIO_0_1,requestAWIO_0_0}; // @[Xbar.scala 64:75]
  assign requestWIO_0_0 = awIn_0_io_deq_bits[0]; // @[Xbar.scala 65:73]
  assign requestWIO_0_1 = awIn_0_io_deq_bits[1]; // @[Xbar.scala 65:73]
  assign _T_27 = {requestARIO_0_1,requestARIO_0_0}; // @[Xbar.scala 93:45]
  assign _T_108 = requestARIO_0_0 & auto_out_0_ar_ready; // @[Mux.scala 27:72]
  assign _T_109 = requestARIO_0_1 & auto_out_1_ar_ready; // @[Mux.scala 27:72]
  assign in_0_ar_ready = _T_108 | _T_109; // @[Mux.scala 27:72]
  assign _T_55 = _T_36 == 3'h0; // @[Xbar.scala 112:22]
  assign _T_54 = _T_37 == _T_27[1]; // @[Xbar.scala 111:75]
  assign _T_56 = _T_55 | _T_54; // @[Xbar.scala 112:34]
  assign _T_57 = _T_36 != 3'h7; // @[Xbar.scala 112:80]
  assign _T_59 = _T_56 & _T_57; // @[Xbar.scala 112:48]
  assign io_in_0_ar_ready = in_0_ar_ready & _T_59; // @[Xbar.scala 130:45]
  assign _T_31 = io_in_0_ar_ready & auto_in_ar_valid; // @[Decoupled.scala 40:37]
  assign _T_127 = auto_out_0_r_valid & requestROI_0_0; // @[Xbar.scala 222:40]
  assign _T_129 = auto_out_1_r_valid & requestROI_1_0; // @[Xbar.scala 222:40]
  assign _T_223 = _T_127 | _T_129; // @[Xbar.scala 246:36]
  assign _T_284 = _T_278_0 & _T_127; // @[Mux.scala 27:72]
  assign _T_285 = _T_278_1 & _T_129; // @[Mux.scala 27:72]
  assign _T_286 = _T_284 | _T_285; // @[Mux.scala 27:72]
  assign in_0_r_valid = _T_222 ? _T_223 : _T_286; // @[Xbar.scala 278:22]
  assign _T_33 = auto_in_r_ready & in_0_r_valid; // @[Decoupled.scala 40:37]
  assign _T_224 = {_T_129,_T_127}; // @[Cat.scala 29:58]
  assign _T_232 = ~_T_231; // @[Arbiter.scala 21:30]
  assign _T_233 = _T_224 & _T_232; // @[Arbiter.scala 21:28]
  assign _T_234 = {_T_233,_T_129,_T_127}; // @[Cat.scala 29:58]
  assign _GEN_18 = {{1'd0}, _T_234[3:1]}; // @[package.scala 208:43]
  assign _T_236 = _T_234 | _GEN_18; // @[package.scala 208:43]
  assign _T_239 = {_T_231, 2'h0}; // @[Arbiter.scala 22:66]
  assign _GEN_19 = {{1'd0}, _T_236[3:1]}; // @[Arbiter.scala 22:58]
  assign _T_240 = _GEN_19 | _T_239; // @[Arbiter.scala 22:58]
  assign _T_243 = _T_240[3:2] & _T_240[1:0]; // @[Arbiter.scala 23:39]
  assign _T_244 = ~_T_243; // @[Arbiter.scala 23:18]
  assign _T_256 = _T_244[0] & _T_127; // @[Xbar.scala 250:63]
  assign _T_279_0 = _T_222 ? _T_256 : _T_278_0; // @[Xbar.scala 262:23]
  assign _T_291 = {auto_out_0_r_bits_id,auto_out_0_r_bits_data,auto_out_0_r_bits_resp,auto_out_0_r_bits_last}; // @[Mux.scala 27:72]
  assign _T_292 = _T_279_0 ? _T_291 : 36'h0; // @[Mux.scala 27:72]
  assign _T_257 = _T_244[1] & _T_129; // @[Xbar.scala 250:63]
  assign _T_279_1 = _T_222 ? _T_257 : _T_278_1; // @[Xbar.scala 262:23]
  assign _T_295 = {auto_out_1_r_bits_id,auto_out_1_r_bits_data,auto_out_1_r_bits_resp,auto_out_1_r_bits_last}; // @[Mux.scala 27:72]
  assign _T_296 = _T_279_1 ? _T_295 : 36'h0; // @[Mux.scala 27:72]
  assign _T_297 = _T_292 | _T_296; // @[Mux.scala 27:72]
  assign in_0_r_bits_last = _T_297[0]; // @[Mux.scala 27:72]
  assign _T_35 = _T_33 & in_0_r_bits_last; // @[Xbar.scala 120:45]
  assign _GEN_20 = {{2'd0}, _T_31}; // @[Xbar.scala 106:30]
  assign _T_39 = _T_36 + _GEN_20; // @[Xbar.scala 106:30]
  assign _GEN_21 = {{2'd0}, _T_35}; // @[Xbar.scala 106:48]
  assign _T_41 = _T_39 - _GEN_21; // @[Xbar.scala 106:48]
  assign _T_42 = ~_T_35; // @[Xbar.scala 107:23]
  assign _T_43 = _T_36 != 3'h0; // @[Xbar.scala 107:43]
  assign _T_44 = _T_42 | _T_43; // @[Xbar.scala 107:34]
  assign _T_46 = _T_44 | reset; // @[Xbar.scala 107:22]
  assign _T_47 = ~_T_46; // @[Xbar.scala 107:22]
  assign _T_48 = ~_T_31; // @[Xbar.scala 108:23]
  assign _T_50 = _T_48 | _T_57; // @[Xbar.scala 108:34]
  assign _T_52 = _T_50 | reset; // @[Xbar.scala 108:22]
  assign _T_53 = ~_T_52; // @[Xbar.scala 108:22]
  assign _T_115 = requestAWIO_0_0 & auto_out_0_aw_ready; // @[Mux.scala 27:72]
  assign _T_116 = requestAWIO_0_1 & auto_out_1_aw_ready; // @[Mux.scala 27:72]
  assign in_0_aw_ready = _T_115 | _T_116; // @[Mux.scala 27:72]
  assign _T_94 = _T_90 | awIn_0_io_enq_ready; // @[Xbar.scala 139:57]
  assign _T_95 = in_0_aw_ready & _T_94; // @[Xbar.scala 139:45]
  assign _T_83 = _T_64 == 3'h0; // @[Xbar.scala 112:22]
  assign _T_82 = _T_65 == _T_20[1]; // @[Xbar.scala 111:75]
  assign _T_84 = _T_83 | _T_82; // @[Xbar.scala 112:34]
  assign _T_85 = _T_64 != 3'h7; // @[Xbar.scala 112:80]
  assign _T_87 = _T_84 & _T_85; // @[Xbar.scala 112:48]
  assign io_in_0_aw_ready = _T_95 & _T_87; // @[Xbar.scala 139:82]
  assign _T_60 = io_in_0_aw_ready & auto_in_aw_valid; // @[Decoupled.scala 40:37]
  assign _T_131 = auto_out_0_b_valid & requestBOI_0_0; // @[Xbar.scala 222:40]
  assign _T_133 = auto_out_1_b_valid & requestBOI_1_0; // @[Xbar.scala 222:40]
  assign _T_305 = _T_131 | _T_133; // @[Xbar.scala 246:36]
  assign _T_366 = _T_360_0 & _T_131; // @[Mux.scala 27:72]
  assign _T_367 = _T_360_1 & _T_133; // @[Mux.scala 27:72]
  assign _T_368 = _T_366 | _T_367; // @[Mux.scala 27:72]
  assign in_0_b_valid = _T_304 ? _T_305 : _T_368; // @[Xbar.scala 278:22]
  assign _T_62 = auto_in_b_ready & in_0_b_valid; // @[Decoupled.scala 40:37]
  assign _GEN_22 = {{2'd0}, _T_60}; // @[Xbar.scala 106:30]
  assign _T_67 = _T_64 + _GEN_22; // @[Xbar.scala 106:30]
  assign _GEN_23 = {{2'd0}, _T_62}; // @[Xbar.scala 106:48]
  assign _T_69 = _T_67 - _GEN_23; // @[Xbar.scala 106:48]
  assign _T_70 = ~_T_62; // @[Xbar.scala 107:23]
  assign _T_71 = _T_64 != 3'h0; // @[Xbar.scala 107:43]
  assign _T_72 = _T_70 | _T_71; // @[Xbar.scala 107:34]
  assign _T_74 = _T_72 | reset; // @[Xbar.scala 107:22]
  assign _T_75 = ~_T_74; // @[Xbar.scala 107:22]
  assign _T_76 = ~_T_60; // @[Xbar.scala 108:23]
  assign _T_78 = _T_76 | _T_85; // @[Xbar.scala 108:34]
  assign _T_80 = _T_78 | reset; // @[Xbar.scala 108:22]
  assign _T_81 = ~_T_80; // @[Xbar.scala 108:22]
  assign in_0_ar_valid = auto_in_ar_valid & _T_59; // @[Xbar.scala 129:45]
  assign _T_92 = auto_in_aw_valid & _T_94; // @[Xbar.scala 138:45]
  assign in_0_aw_valid = _T_92 & _T_87; // @[Xbar.scala 138:82]
  assign _T_97 = ~_T_90; // @[Xbar.scala 140:54]
  assign _T_99 = awIn_0_io_enq_ready & awIn_0_io_enq_valid; // @[Decoupled.scala 40:37]
  assign _GEN_2 = _T_99 | _T_90; // @[Xbar.scala 141:38]
  assign _T_100 = in_0_aw_ready & in_0_aw_valid; // @[Decoupled.scala 40:37]
  assign in_0_w_valid = auto_in_w_valid & awIn_0_io_deq_valid; // @[Xbar.scala 145:43]
  assign _T_122 = requestWIO_0_0 & auto_out_0_w_ready; // @[Mux.scala 27:72]
  assign _T_123 = requestWIO_0_1 & auto_out_1_w_ready; // @[Mux.scala 27:72]
  assign in_0_w_ready = _T_122 | _T_123; // @[Mux.scala 27:72]
  assign _T_103 = auto_in_w_valid & auto_in_w_bits_last; // @[Xbar.scala 147:50]
  assign out_0_ar_valid = in_0_ar_valid & requestARIO_0_0; // @[Xbar.scala 222:40]
  assign out_1_ar_valid = in_0_ar_valid & requestARIO_0_1; // @[Xbar.scala 222:40]
  assign out_0_aw_valid = in_0_aw_valid & requestAWIO_0_0; // @[Xbar.scala 222:40]
  assign out_1_aw_valid = in_0_aw_valid & requestAWIO_0_1; // @[Xbar.scala 222:40]
  assign _T_140 = ~out_0_aw_valid; // @[Xbar.scala 256:60]
  assign _T_146 = _T_140 | out_0_aw_valid; // @[Xbar.scala 258:23]
  assign _T_148 = _T_146 | reset; // @[Xbar.scala 258:12]
  assign _T_149 = ~_T_148; // @[Xbar.scala 258:12]
  assign _T_161 = ~out_0_ar_valid; // @[Xbar.scala 256:60]
  assign _T_167 = _T_161 | out_0_ar_valid; // @[Xbar.scala 258:23]
  assign _T_169 = _T_167 | reset; // @[Xbar.scala 258:12]
  assign _T_170 = ~_T_169; // @[Xbar.scala 258:12]
  assign _T_184 = ~out_1_aw_valid; // @[Xbar.scala 256:60]
  assign _T_190 = _T_184 | out_1_aw_valid; // @[Xbar.scala 258:23]
  assign _T_192 = _T_190 | reset; // @[Xbar.scala 258:12]
  assign _T_193 = ~_T_192; // @[Xbar.scala 258:12]
  assign _T_205 = ~out_1_ar_valid; // @[Xbar.scala 256:60]
  assign _T_211 = _T_205 | out_1_ar_valid; // @[Xbar.scala 258:23]
  assign _T_213 = _T_211 | reset; // @[Xbar.scala 258:12]
  assign _T_214 = ~_T_213; // @[Xbar.scala 258:12]
  assign _T_245 = _T_224 != 2'h0; // @[Arbiter.scala 24:27]
  assign _T_246 = _T_222 & _T_245; // @[Arbiter.scala 24:18]
  assign _T_247 = _T_244 & _T_224; // @[Arbiter.scala 25:29]
  assign _T_248 = {_T_247, 1'h0}; // @[package.scala 199:48]
  assign _T_250 = _T_247 | _T_248[1:0]; // @[package.scala 199:43]
  assign _T_260 = _T_256 | _T_257; // @[Xbar.scala 255:50]
  assign _T_262 = ~_T_256; // @[Xbar.scala 256:60]
  assign _T_265 = ~_T_257; // @[Xbar.scala 256:60]
  assign _T_266 = _T_262 | _T_265; // @[Xbar.scala 256:57]
  assign _T_269 = _T_266 | reset; // @[Xbar.scala 256:11]
  assign _T_270 = ~_T_269; // @[Xbar.scala 256:11]
  assign _T_271 = ~_T_223; // @[Xbar.scala 258:13]
  assign _T_273 = _T_271 | _T_260; // @[Xbar.scala 258:23]
  assign _T_275 = _T_273 | reset; // @[Xbar.scala 258:12]
  assign _T_276 = ~_T_275; // @[Xbar.scala 258:12]
  assign _GEN_13 = _T_223 ? 1'h0 : _T_222; // @[Xbar.scala 266:21]
  assign _GEN_14 = _T_33 | _GEN_13; // @[Xbar.scala 267:24]
  assign _T_281_0 = _T_222 ? _T_244[0] : _T_278_0; // @[Xbar.scala 270:24]
  assign _T_281_1 = _T_222 ? _T_244[1] : _T_278_1; // @[Xbar.scala 270:24]
  assign _T_306 = {_T_133,_T_131}; // @[Cat.scala 29:58]
  assign _T_314 = ~_T_313; // @[Arbiter.scala 21:30]
  assign _T_315 = _T_306 & _T_314; // @[Arbiter.scala 21:28]
  assign _T_316 = {_T_315,_T_133,_T_131}; // @[Cat.scala 29:58]
  assign _GEN_24 = {{1'd0}, _T_316[3:1]}; // @[package.scala 208:43]
  assign _T_318 = _T_316 | _GEN_24; // @[package.scala 208:43]
  assign _T_321 = {_T_313, 2'h0}; // @[Arbiter.scala 22:66]
  assign _GEN_25 = {{1'd0}, _T_318[3:1]}; // @[Arbiter.scala 22:58]
  assign _T_322 = _GEN_25 | _T_321; // @[Arbiter.scala 22:58]
  assign _T_325 = _T_322[3:2] & _T_322[1:0]; // @[Arbiter.scala 23:39]
  assign _T_326 = ~_T_325; // @[Arbiter.scala 23:18]
  assign _T_327 = _T_306 != 2'h0; // @[Arbiter.scala 24:27]
  assign _T_328 = _T_304 & _T_327; // @[Arbiter.scala 24:18]
  assign _T_329 = _T_326 & _T_306; // @[Arbiter.scala 25:29]
  assign _T_330 = {_T_329, 1'h0}; // @[package.scala 199:48]
  assign _T_332 = _T_329 | _T_330[1:0]; // @[package.scala 199:43]
  assign _T_338 = _T_326[0] & _T_131; // @[Xbar.scala 250:63]
  assign _T_339 = _T_326[1] & _T_133; // @[Xbar.scala 250:63]
  assign _T_342 = _T_338 | _T_339; // @[Xbar.scala 255:50]
  assign _T_344 = ~_T_338; // @[Xbar.scala 256:60]
  assign _T_347 = ~_T_339; // @[Xbar.scala 256:60]
  assign _T_348 = _T_344 | _T_347; // @[Xbar.scala 256:57]
  assign _T_351 = _T_348 | reset; // @[Xbar.scala 256:11]
  assign _T_352 = ~_T_351; // @[Xbar.scala 256:11]
  assign _T_353 = ~_T_305; // @[Xbar.scala 258:13]
  assign _T_355 = _T_353 | _T_342; // @[Xbar.scala 258:23]
  assign _T_357 = _T_355 | reset; // @[Xbar.scala 258:12]
  assign _T_358 = ~_T_357; // @[Xbar.scala 258:12]
  assign _T_361_0 = _T_304 ? _T_338 : _T_360_0; // @[Xbar.scala 262:23]
  assign _T_361_1 = _T_304 ? _T_339 : _T_360_1; // @[Xbar.scala 262:23]
  assign _GEN_16 = _T_305 ? 1'h0 : _T_304; // @[Xbar.scala 266:21]
  assign _GEN_17 = _T_62 | _GEN_16; // @[Xbar.scala 267:24]
  assign _T_363_0 = _T_304 ? _T_326[0] : _T_360_0; // @[Xbar.scala 270:24]
  assign _T_363_1 = _T_304 ? _T_326[1] : _T_360_1; // @[Xbar.scala 270:24]
  assign _T_371 = {auto_out_0_b_bits_id,auto_out_0_b_bits_resp}; // @[Mux.scala 27:72]
  assign _T_372 = _T_361_0 ? _T_371 : 3'h0; // @[Mux.scala 27:72]
  assign _T_373 = {auto_out_1_b_bits_id,auto_out_1_b_bits_resp}; // @[Mux.scala 27:72]
  assign _T_374 = _T_361_1 ? _T_373 : 3'h0; // @[Mux.scala 27:72]
  assign _T_375 = _T_372 | _T_374; // @[Mux.scala 27:72]
  assign auto_in_aw_ready = _T_95 & _T_87; // @[LazyModule.scala 173:31]
  assign auto_in_w_ready = in_0_w_ready & awIn_0_io_deq_valid; // @[LazyModule.scala 173:31]
  assign auto_in_b_valid = _T_304 ? _T_305 : _T_368; // @[LazyModule.scala 173:31]
  assign auto_in_b_bits_resp = _T_375[1:0]; // @[LazyModule.scala 173:31]
  assign auto_in_ar_ready = in_0_ar_ready & _T_59; // @[LazyModule.scala 173:31]
  assign auto_in_r_valid = _T_222 ? _T_223 : _T_286; // @[LazyModule.scala 173:31]
  assign auto_in_r_bits_data = _T_297[34:3]; // @[LazyModule.scala 173:31]
  assign auto_in_r_bits_resp = _T_297[2:1]; // @[LazyModule.scala 173:31]
  assign auto_in_r_bits_last = _T_297[0]; // @[LazyModule.scala 173:31]
  assign auto_out_1_aw_valid = in_0_aw_valid & requestAWIO_0_1; // @[LazyModule.scala 173:49]
  assign auto_out_1_aw_bits_id = auto_in_aw_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_1_aw_bits_addr = auto_in_aw_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_1_aw_bits_size = auto_in_aw_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_1_w_valid = in_0_w_valid & requestWIO_0_1; // @[LazyModule.scala 173:49]
  assign auto_out_1_w_bits_data = auto_in_w_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_1_w_bits_strb = auto_in_w_bits_strb; // @[LazyModule.scala 173:49]
  assign auto_out_1_w_bits_last = auto_in_w_bits_last; // @[LazyModule.scala 173:49]
  assign auto_out_1_b_ready = auto_in_b_ready & _T_363_1; // @[LazyModule.scala 173:49]
  assign auto_out_1_ar_valid = in_0_ar_valid & requestARIO_0_1; // @[LazyModule.scala 173:49]
  assign auto_out_1_ar_bits_id = auto_in_ar_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_1_ar_bits_addr = auto_in_ar_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_1_ar_bits_size = auto_in_ar_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_1_r_ready = auto_in_r_ready & _T_281_1; // @[LazyModule.scala 173:49]
  assign auto_out_0_aw_valid = in_0_aw_valid & requestAWIO_0_0; // @[LazyModule.scala 173:49]
  assign auto_out_0_aw_bits_id = auto_in_aw_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_0_aw_bits_addr = auto_in_aw_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_0_aw_bits_size = auto_in_aw_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_0_w_valid = in_0_w_valid & requestWIO_0_0; // @[LazyModule.scala 173:49]
  assign auto_out_0_w_bits_data = auto_in_w_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_0_w_bits_strb = auto_in_w_bits_strb; // @[LazyModule.scala 173:49]
  assign auto_out_0_w_bits_last = auto_in_w_bits_last; // @[LazyModule.scala 173:49]
  assign auto_out_0_b_ready = auto_in_b_ready & _T_363_0; // @[LazyModule.scala 173:49]
  assign auto_out_0_ar_valid = in_0_ar_valid & requestARIO_0_0; // @[LazyModule.scala 173:49]
  assign auto_out_0_ar_bits_id = auto_in_ar_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_0_ar_bits_addr = auto_in_ar_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_0_ar_bits_size = auto_in_ar_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_0_r_ready = auto_in_r_ready & _T_281_0; // @[LazyModule.scala 173:49]
  assign awIn_0_clock = clock;
  assign awIn_0_reset = reset;
  assign awIn_0_io_enq_valid = auto_in_aw_valid & _T_97; // @[Xbar.scala 140:30]
  assign awIn_0_io_enq_bits = {requestAWIO_0_1,requestAWIO_0_0}; // @[Xbar.scala 64:57]
  assign awIn_0_io_deq_ready = _T_103 & in_0_w_ready; // @[Xbar.scala 147:30]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_36 = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_37 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_222 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_278_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_278_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_231 = _RAND_5[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_90 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_64 = _RAND_7[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_65 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_304 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_360_0 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_360_1 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_313 = _RAND_12[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      _T_36 <= 3'h0;
    end else begin
      _T_36 <= _T_41;
    end
    if (_T_31) begin
      _T_37 <= _T_27[1];
    end
    _T_222 <= reset | _GEN_14;
    if (reset) begin
      _T_278_0 <= 1'h0;
    end else if (_T_222) begin
      _T_278_0 <= _T_256;
    end
    if (reset) begin
      _T_278_1 <= 1'h0;
    end else if (_T_222) begin
      _T_278_1 <= _T_257;
    end
    if (reset) begin
      _T_231 <= 2'h3;
    end else if (_T_246) begin
      _T_231 <= _T_250;
    end
    if (reset) begin
      _T_90 <= 1'h0;
    end else if (_T_100) begin
      _T_90 <= 1'h0;
    end else begin
      _T_90 <= _GEN_2;
    end
    if (reset) begin
      _T_64 <= 3'h0;
    end else begin
      _T_64 <= _T_69;
    end
    if (_T_60) begin
      _T_65 <= _T_20[1];
    end
    _T_304 <= reset | _GEN_17;
    if (reset) begin
      _T_360_0 <= 1'h0;
    end else if (_T_304) begin
      _T_360_0 <= _T_338;
    end
    if (reset) begin
      _T_360_1 <= 1'h0;
    end else if (_T_304) begin
      _T_360_1 <= _T_339;
    end
    if (reset) begin
      _T_313 <= 2'h3;
    end else if (_T_328) begin
      _T_313 <= _T_332;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_47) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:107 assert (!resp_fire || count =/= UInt(0))\n"); // @[Xbar.scala 107:22]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_47) begin
          $fatal; // @[Xbar.scala 107:22]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_53) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:108 assert (!req_fire  || count =/= UInt(flight))\n"); // @[Xbar.scala 108:22]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_53) begin
          $fatal; // @[Xbar.scala 108:22]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_75) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:107 assert (!resp_fire || count =/= UInt(0))\n"); // @[Xbar.scala 107:22]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_75) begin
          $fatal; // @[Xbar.scala 107:22]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_81) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:108 assert (!req_fire  || count =/= UInt(flight))\n"); // @[Xbar.scala 108:22]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_81) begin
          $fatal; // @[Xbar.scala 108:22]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_149) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_149) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_170) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_170) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_193) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_193) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_214) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_214) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_270) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:256 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n"); // @[Xbar.scala 256:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_270) begin
          $fatal; // @[Xbar.scala 256:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_276) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_276) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_352) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:256 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n"); // @[Xbar.scala 256:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_352) begin
          $fatal; // @[Xbar.scala 256:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_358) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_358) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module Queue_25(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input         io_enq_bits_id,
  input  [29:0] io_enq_bits_addr,
  input  [2:0]  io_enq_bits_size,
  input         io_deq_ready,
  output        io_deq_valid,
  output        io_deq_bits_id,
  output [29:0] io_deq_bits_addr,
  output [2:0]  io_deq_bits_size
);
  reg  _T_id [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_0;
  wire  _T_id__T_18_data; // @[Decoupled.scala 209:24]
  wire  _T_id__T_18_addr; // @[Decoupled.scala 209:24]
  wire  _T_id__T_10_data; // @[Decoupled.scala 209:24]
  wire  _T_id__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T_id__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T_id__T_10_en; // @[Decoupled.scala 209:24]
  reg [29:0] _T_addr [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_1;
  wire [29:0] _T_addr__T_18_data; // @[Decoupled.scala 209:24]
  wire  _T_addr__T_18_addr; // @[Decoupled.scala 209:24]
  wire [29:0] _T_addr__T_10_data; // @[Decoupled.scala 209:24]
  wire  _T_addr__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T_addr__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T_addr__T_10_en; // @[Decoupled.scala 209:24]
  reg [2:0] _T_size [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_2;
  wire [2:0] _T_size__T_18_data; // @[Decoupled.scala 209:24]
  wire  _T_size__T_18_addr; // @[Decoupled.scala 209:24]
  wire [2:0] _T_size__T_10_data; // @[Decoupled.scala 209:24]
  wire  _T_size__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T_size__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T_size__T_10_en; // @[Decoupled.scala 209:24]
  reg  value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_3;
  reg  value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_4;
  reg  _T_1; // @[Decoupled.scala 212:35]
  reg [31:0] _RAND_5;
  wire  _T_2; // @[Decoupled.scala 214:41]
  wire  _T_3; // @[Decoupled.scala 215:36]
  wire  _T_4; // @[Decoupled.scala 215:33]
  wire  _T_5; // @[Decoupled.scala 216:32]
  wire  _T_6; // @[Decoupled.scala 40:37]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _T_12; // @[Counter.scala 39:22]
  wire  _T_14; // @[Counter.scala 39:22]
  wire  _T_15; // @[Decoupled.scala 227:16]
  assign _T_id__T_18_addr = value_1;
  assign _T_id__T_18_data = _T_id[_T_id__T_18_addr]; // @[Decoupled.scala 209:24]
  assign _T_id__T_10_data = io_enq_bits_id;
  assign _T_id__T_10_addr = value;
  assign _T_id__T_10_mask = 1'h1;
  assign _T_id__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_addr__T_18_addr = value_1;
  assign _T_addr__T_18_data = _T_addr[_T_addr__T_18_addr]; // @[Decoupled.scala 209:24]
  assign _T_addr__T_10_data = io_enq_bits_addr;
  assign _T_addr__T_10_addr = value;
  assign _T_addr__T_10_mask = 1'h1;
  assign _T_addr__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_size__T_18_addr = value_1;
  assign _T_size__T_18_data = _T_size[_T_size__T_18_addr]; // @[Decoupled.scala 209:24]
  assign _T_size__T_10_data = io_enq_bits_size;
  assign _T_size__T_10_addr = value;
  assign _T_size__T_10_mask = 1'h1;
  assign _T_size__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_2 = value == value_1; // @[Decoupled.scala 214:41]
  assign _T_3 = ~_T_1; // @[Decoupled.scala 215:36]
  assign _T_4 = _T_2 & _T_3; // @[Decoupled.scala 215:33]
  assign _T_5 = _T_2 & _T_1; // @[Decoupled.scala 216:32]
  assign _T_6 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  assign _T_8 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  assign _T_12 = value + 1'h1; // @[Counter.scala 39:22]
  assign _T_14 = value_1 + 1'h1; // @[Counter.scala 39:22]
  assign _T_15 = _T_6 != _T_8; // @[Decoupled.scala 227:16]
  assign io_enq_ready = ~_T_5; // @[Decoupled.scala 232:16]
  assign io_deq_valid = ~_T_4; // @[Decoupled.scala 231:16]
  assign io_deq_bits_id = _T_id__T_18_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_addr = _T_addr__T_18_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_size = _T_size__T_18_data; // @[Decoupled.scala 233:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_id[initvar] = _RAND_0[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_addr[initvar] = _RAND_1[29:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_size[initvar] = _RAND_2[2:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  value = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  value_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_1 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T_id__T_10_en & _T_id__T_10_mask) begin
      _T_id[_T_id__T_10_addr] <= _T_id__T_10_data; // @[Decoupled.scala 209:24]
    end
    if(_T_addr__T_10_en & _T_addr__T_10_mask) begin
      _T_addr[_T_addr__T_10_addr] <= _T_addr__T_10_data; // @[Decoupled.scala 209:24]
    end
    if(_T_size__T_10_en & _T_size__T_10_mask) begin
      _T_size[_T_size__T_10_addr] <= _T_size__T_10_data; // @[Decoupled.scala 209:24]
    end
    if (reset) begin
      value <= 1'h0;
    end else if (_T_6) begin
      value <= _T_12;
    end
    if (reset) begin
      value_1 <= 1'h0;
    end else if (_T_8) begin
      value_1 <= _T_14;
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else if (_T_15) begin
      _T_1 <= _T_6;
    end
  end
endmodule
module Queue_26(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [31:0] io_enq_bits_data,
  input  [3:0]  io_enq_bits_strb,
  input         io_enq_bits_last,
  input         io_deq_ready,
  output        io_deq_valid,
  output [31:0] io_deq_bits_data,
  output [3:0]  io_deq_bits_strb,
  output        io_deq_bits_last
);
  reg [31:0] _T_data [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_0;
  wire [31:0] _T_data__T_18_data; // @[Decoupled.scala 209:24]
  wire  _T_data__T_18_addr; // @[Decoupled.scala 209:24]
  wire [31:0] _T_data__T_10_data; // @[Decoupled.scala 209:24]
  wire  _T_data__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T_data__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T_data__T_10_en; // @[Decoupled.scala 209:24]
  reg [3:0] _T_strb [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_1;
  wire [3:0] _T_strb__T_18_data; // @[Decoupled.scala 209:24]
  wire  _T_strb__T_18_addr; // @[Decoupled.scala 209:24]
  wire [3:0] _T_strb__T_10_data; // @[Decoupled.scala 209:24]
  wire  _T_strb__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T_strb__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T_strb__T_10_en; // @[Decoupled.scala 209:24]
  reg  _T_last [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_2;
  wire  _T_last__T_18_data; // @[Decoupled.scala 209:24]
  wire  _T_last__T_18_addr; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_data; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_en; // @[Decoupled.scala 209:24]
  reg  value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_3;
  reg  value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_4;
  reg  _T_1; // @[Decoupled.scala 212:35]
  reg [31:0] _RAND_5;
  wire  _T_2; // @[Decoupled.scala 214:41]
  wire  _T_3; // @[Decoupled.scala 215:36]
  wire  _T_4; // @[Decoupled.scala 215:33]
  wire  _T_5; // @[Decoupled.scala 216:32]
  wire  _T_6; // @[Decoupled.scala 40:37]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _T_12; // @[Counter.scala 39:22]
  wire  _T_14; // @[Counter.scala 39:22]
  wire  _T_15; // @[Decoupled.scala 227:16]
  assign _T_data__T_18_addr = value_1;
  assign _T_data__T_18_data = _T_data[_T_data__T_18_addr]; // @[Decoupled.scala 209:24]
  assign _T_data__T_10_data = io_enq_bits_data;
  assign _T_data__T_10_addr = value;
  assign _T_data__T_10_mask = 1'h1;
  assign _T_data__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_strb__T_18_addr = value_1;
  assign _T_strb__T_18_data = _T_strb[_T_strb__T_18_addr]; // @[Decoupled.scala 209:24]
  assign _T_strb__T_10_data = io_enq_bits_strb;
  assign _T_strb__T_10_addr = value;
  assign _T_strb__T_10_mask = 1'h1;
  assign _T_strb__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_last__T_18_addr = value_1;
  assign _T_last__T_18_data = _T_last[_T_last__T_18_addr]; // @[Decoupled.scala 209:24]
  assign _T_last__T_10_data = io_enq_bits_last;
  assign _T_last__T_10_addr = value;
  assign _T_last__T_10_mask = 1'h1;
  assign _T_last__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_2 = value == value_1; // @[Decoupled.scala 214:41]
  assign _T_3 = ~_T_1; // @[Decoupled.scala 215:36]
  assign _T_4 = _T_2 & _T_3; // @[Decoupled.scala 215:33]
  assign _T_5 = _T_2 & _T_1; // @[Decoupled.scala 216:32]
  assign _T_6 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  assign _T_8 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  assign _T_12 = value + 1'h1; // @[Counter.scala 39:22]
  assign _T_14 = value_1 + 1'h1; // @[Counter.scala 39:22]
  assign _T_15 = _T_6 != _T_8; // @[Decoupled.scala 227:16]
  assign io_enq_ready = ~_T_5; // @[Decoupled.scala 232:16]
  assign io_deq_valid = ~_T_4; // @[Decoupled.scala 231:16]
  assign io_deq_bits_data = _T_data__T_18_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_strb = _T_strb__T_18_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_last = _T_last__T_18_data; // @[Decoupled.scala 233:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_data[initvar] = _RAND_0[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_strb[initvar] = _RAND_1[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_last[initvar] = _RAND_2[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  value = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  value_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_1 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T_data__T_10_en & _T_data__T_10_mask) begin
      _T_data[_T_data__T_10_addr] <= _T_data__T_10_data; // @[Decoupled.scala 209:24]
    end
    if(_T_strb__T_10_en & _T_strb__T_10_mask) begin
      _T_strb[_T_strb__T_10_addr] <= _T_strb__T_10_data; // @[Decoupled.scala 209:24]
    end
    if(_T_last__T_10_en & _T_last__T_10_mask) begin
      _T_last[_T_last__T_10_addr] <= _T_last__T_10_data; // @[Decoupled.scala 209:24]
    end
    if (reset) begin
      value <= 1'h0;
    end else if (_T_6) begin
      value <= _T_12;
    end
    if (reset) begin
      value_1 <= 1'h0;
    end else if (_T_8) begin
      value_1 <= _T_14;
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else if (_T_15) begin
      _T_1 <= _T_6;
    end
  end
endmodule
module Queue_27(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input        io_enq_bits_id,
  input  [1:0] io_enq_bits_resp,
  input        io_deq_ready,
  output       io_deq_valid,
  output       io_deq_bits_id,
  output [1:0] io_deq_bits_resp
);
  reg  _T_id [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_0;
  wire  _T_id__T_18_data; // @[Decoupled.scala 209:24]
  wire  _T_id__T_18_addr; // @[Decoupled.scala 209:24]
  wire  _T_id__T_10_data; // @[Decoupled.scala 209:24]
  wire  _T_id__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T_id__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T_id__T_10_en; // @[Decoupled.scala 209:24]
  reg [1:0] _T_resp [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_1;
  wire [1:0] _T_resp__T_18_data; // @[Decoupled.scala 209:24]
  wire  _T_resp__T_18_addr; // @[Decoupled.scala 209:24]
  wire [1:0] _T_resp__T_10_data; // @[Decoupled.scala 209:24]
  wire  _T_resp__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T_resp__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T_resp__T_10_en; // @[Decoupled.scala 209:24]
  reg  value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_2;
  reg  value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_3;
  reg  _T_1; // @[Decoupled.scala 212:35]
  reg [31:0] _RAND_4;
  wire  _T_2; // @[Decoupled.scala 214:41]
  wire  _T_3; // @[Decoupled.scala 215:36]
  wire  _T_4; // @[Decoupled.scala 215:33]
  wire  _T_5; // @[Decoupled.scala 216:32]
  wire  _T_6; // @[Decoupled.scala 40:37]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _T_12; // @[Counter.scala 39:22]
  wire  _T_14; // @[Counter.scala 39:22]
  wire  _T_15; // @[Decoupled.scala 227:16]
  assign _T_id__T_18_addr = value_1;
  assign _T_id__T_18_data = _T_id[_T_id__T_18_addr]; // @[Decoupled.scala 209:24]
  assign _T_id__T_10_data = io_enq_bits_id;
  assign _T_id__T_10_addr = value;
  assign _T_id__T_10_mask = 1'h1;
  assign _T_id__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_resp__T_18_addr = value_1;
  assign _T_resp__T_18_data = _T_resp[_T_resp__T_18_addr]; // @[Decoupled.scala 209:24]
  assign _T_resp__T_10_data = io_enq_bits_resp;
  assign _T_resp__T_10_addr = value;
  assign _T_resp__T_10_mask = 1'h1;
  assign _T_resp__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_2 = value == value_1; // @[Decoupled.scala 214:41]
  assign _T_3 = ~_T_1; // @[Decoupled.scala 215:36]
  assign _T_4 = _T_2 & _T_3; // @[Decoupled.scala 215:33]
  assign _T_5 = _T_2 & _T_1; // @[Decoupled.scala 216:32]
  assign _T_6 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  assign _T_8 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  assign _T_12 = value + 1'h1; // @[Counter.scala 39:22]
  assign _T_14 = value_1 + 1'h1; // @[Counter.scala 39:22]
  assign _T_15 = _T_6 != _T_8; // @[Decoupled.scala 227:16]
  assign io_enq_ready = ~_T_5; // @[Decoupled.scala 232:16]
  assign io_deq_valid = ~_T_4; // @[Decoupled.scala 231:16]
  assign io_deq_bits_id = _T_id__T_18_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_resp = _T_resp__T_18_data; // @[Decoupled.scala 233:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_id[initvar] = _RAND_0[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_resp[initvar] = _RAND_1[1:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  value = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  value_1 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T_id__T_10_en & _T_id__T_10_mask) begin
      _T_id[_T_id__T_10_addr] <= _T_id__T_10_data; // @[Decoupled.scala 209:24]
    end
    if(_T_resp__T_10_en & _T_resp__T_10_mask) begin
      _T_resp[_T_resp__T_10_addr] <= _T_resp__T_10_data; // @[Decoupled.scala 209:24]
    end
    if (reset) begin
      value <= 1'h0;
    end else if (_T_6) begin
      value <= _T_12;
    end
    if (reset) begin
      value_1 <= 1'h0;
    end else if (_T_8) begin
      value_1 <= _T_14;
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else if (_T_15) begin
      _T_1 <= _T_6;
    end
  end
endmodule
module Queue_29(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input         io_enq_bits_id,
  input  [31:0] io_enq_bits_data,
  input  [1:0]  io_enq_bits_resp,
  input         io_enq_bits_last,
  input         io_deq_ready,
  output        io_deq_valid,
  output        io_deq_bits_id,
  output [31:0] io_deq_bits_data,
  output [1:0]  io_deq_bits_resp,
  output        io_deq_bits_last
);
  reg  _T_id [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_0;
  wire  _T_id__T_18_data; // @[Decoupled.scala 209:24]
  wire  _T_id__T_18_addr; // @[Decoupled.scala 209:24]
  wire  _T_id__T_10_data; // @[Decoupled.scala 209:24]
  wire  _T_id__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T_id__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T_id__T_10_en; // @[Decoupled.scala 209:24]
  reg [31:0] _T_data [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_1;
  wire [31:0] _T_data__T_18_data; // @[Decoupled.scala 209:24]
  wire  _T_data__T_18_addr; // @[Decoupled.scala 209:24]
  wire [31:0] _T_data__T_10_data; // @[Decoupled.scala 209:24]
  wire  _T_data__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T_data__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T_data__T_10_en; // @[Decoupled.scala 209:24]
  reg [1:0] _T_resp [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_2;
  wire [1:0] _T_resp__T_18_data; // @[Decoupled.scala 209:24]
  wire  _T_resp__T_18_addr; // @[Decoupled.scala 209:24]
  wire [1:0] _T_resp__T_10_data; // @[Decoupled.scala 209:24]
  wire  _T_resp__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T_resp__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T_resp__T_10_en; // @[Decoupled.scala 209:24]
  reg  _T_last [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_3;
  wire  _T_last__T_18_data; // @[Decoupled.scala 209:24]
  wire  _T_last__T_18_addr; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_data; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_en; // @[Decoupled.scala 209:24]
  reg  value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_4;
  reg  value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  reg  _T_1; // @[Decoupled.scala 212:35]
  reg [31:0] _RAND_6;
  wire  _T_2; // @[Decoupled.scala 214:41]
  wire  _T_3; // @[Decoupled.scala 215:36]
  wire  _T_4; // @[Decoupled.scala 215:33]
  wire  _T_5; // @[Decoupled.scala 216:32]
  wire  _T_6; // @[Decoupled.scala 40:37]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _T_12; // @[Counter.scala 39:22]
  wire  _T_14; // @[Counter.scala 39:22]
  wire  _T_15; // @[Decoupled.scala 227:16]
  assign _T_id__T_18_addr = value_1;
  assign _T_id__T_18_data = _T_id[_T_id__T_18_addr]; // @[Decoupled.scala 209:24]
  assign _T_id__T_10_data = io_enq_bits_id;
  assign _T_id__T_10_addr = value;
  assign _T_id__T_10_mask = 1'h1;
  assign _T_id__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_data__T_18_addr = value_1;
  assign _T_data__T_18_data = _T_data[_T_data__T_18_addr]; // @[Decoupled.scala 209:24]
  assign _T_data__T_10_data = io_enq_bits_data;
  assign _T_data__T_10_addr = value;
  assign _T_data__T_10_mask = 1'h1;
  assign _T_data__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_resp__T_18_addr = value_1;
  assign _T_resp__T_18_data = _T_resp[_T_resp__T_18_addr]; // @[Decoupled.scala 209:24]
  assign _T_resp__T_10_data = io_enq_bits_resp;
  assign _T_resp__T_10_addr = value;
  assign _T_resp__T_10_mask = 1'h1;
  assign _T_resp__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_last__T_18_addr = value_1;
  assign _T_last__T_18_data = _T_last[_T_last__T_18_addr]; // @[Decoupled.scala 209:24]
  assign _T_last__T_10_data = io_enq_bits_last;
  assign _T_last__T_10_addr = value;
  assign _T_last__T_10_mask = 1'h1;
  assign _T_last__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_2 = value == value_1; // @[Decoupled.scala 214:41]
  assign _T_3 = ~_T_1; // @[Decoupled.scala 215:36]
  assign _T_4 = _T_2 & _T_3; // @[Decoupled.scala 215:33]
  assign _T_5 = _T_2 & _T_1; // @[Decoupled.scala 216:32]
  assign _T_6 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  assign _T_8 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  assign _T_12 = value + 1'h1; // @[Counter.scala 39:22]
  assign _T_14 = value_1 + 1'h1; // @[Counter.scala 39:22]
  assign _T_15 = _T_6 != _T_8; // @[Decoupled.scala 227:16]
  assign io_enq_ready = ~_T_5; // @[Decoupled.scala 232:16]
  assign io_deq_valid = ~_T_4; // @[Decoupled.scala 231:16]
  assign io_deq_bits_id = _T_id__T_18_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_data = _T_data__T_18_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_resp = _T_resp__T_18_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_last = _T_last__T_18_data; // @[Decoupled.scala 233:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_id[initvar] = _RAND_0[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_data[initvar] = _RAND_1[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_resp[initvar] = _RAND_2[1:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_last[initvar] = _RAND_3[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  value = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value_1 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_1 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T_id__T_10_en & _T_id__T_10_mask) begin
      _T_id[_T_id__T_10_addr] <= _T_id__T_10_data; // @[Decoupled.scala 209:24]
    end
    if(_T_data__T_10_en & _T_data__T_10_mask) begin
      _T_data[_T_data__T_10_addr] <= _T_data__T_10_data; // @[Decoupled.scala 209:24]
    end
    if(_T_resp__T_10_en & _T_resp__T_10_mask) begin
      _T_resp[_T_resp__T_10_addr] <= _T_resp__T_10_data; // @[Decoupled.scala 209:24]
    end
    if(_T_last__T_10_en & _T_last__T_10_mask) begin
      _T_last[_T_last__T_10_addr] <= _T_last__T_10_data; // @[Decoupled.scala 209:24]
    end
    if (reset) begin
      value <= 1'h0;
    end else if (_T_6) begin
      value <= _T_12;
    end
    if (reset) begin
      value_1 <= 1'h0;
    end else if (_T_8) begin
      value_1 <= _T_14;
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else if (_T_15) begin
      _T_1 <= _T_6;
    end
  end
endmodule
module AXI4Buffer(
  input         clock,
  input         reset,
  output        auto_in_aw_ready,
  input         auto_in_aw_valid,
  input         auto_in_aw_bits_id,
  input  [29:0] auto_in_aw_bits_addr,
  input  [2:0]  auto_in_aw_bits_size,
  output        auto_in_w_ready,
  input         auto_in_w_valid,
  input  [31:0] auto_in_w_bits_data,
  input  [3:0]  auto_in_w_bits_strb,
  input         auto_in_w_bits_last,
  input         auto_in_b_ready,
  output        auto_in_b_valid,
  output        auto_in_b_bits_id,
  output [1:0]  auto_in_b_bits_resp,
  output        auto_in_ar_ready,
  input         auto_in_ar_valid,
  input         auto_in_ar_bits_id,
  input  [29:0] auto_in_ar_bits_addr,
  input  [2:0]  auto_in_ar_bits_size,
  input         auto_in_r_ready,
  output        auto_in_r_valid,
  output        auto_in_r_bits_id,
  output [31:0] auto_in_r_bits_data,
  output [1:0]  auto_in_r_bits_resp,
  output        auto_in_r_bits_last,
  input         auto_out_aw_ready,
  output        auto_out_aw_valid,
  output        auto_out_aw_bits_id,
  output [29:0] auto_out_aw_bits_addr,
  input         auto_out_w_ready,
  output        auto_out_w_valid,
  output [31:0] auto_out_w_bits_data,
  output [3:0]  auto_out_w_bits_strb,
  output        auto_out_w_bits_last,
  output        auto_out_b_ready,
  input         auto_out_b_valid,
  input         auto_out_b_bits_id,
  input  [1:0]  auto_out_b_bits_resp,
  input         auto_out_ar_ready,
  output        auto_out_ar_valid,
  output        auto_out_ar_bits_id,
  output [29:0] auto_out_ar_bits_addr,
  output [2:0]  auto_out_ar_bits_size,
  output        auto_out_r_ready,
  input         auto_out_r_valid,
  input         auto_out_r_bits_id,
  input  [31:0] auto_out_r_bits_data,
  input  [1:0]  auto_out_r_bits_resp,
  input         auto_out_r_bits_last
);
  wire  Queue_clock; // @[Decoupled.scala 287:21]
  wire  Queue_reset; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_id; // @[Decoupled.scala 287:21]
  wire [29:0] Queue_io_enq_bits_addr; // @[Decoupled.scala 287:21]
  wire [2:0] Queue_io_enq_bits_size; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_id; // @[Decoupled.scala 287:21]
  wire [29:0] Queue_io_deq_bits_addr; // @[Decoupled.scala 287:21]
  wire [2:0] Queue_io_deq_bits_size; // @[Decoupled.scala 287:21]
  wire  Queue_1_clock; // @[Decoupled.scala 287:21]
  wire  Queue_1_reset; // @[Decoupled.scala 287:21]
  wire  Queue_1_io_enq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_1_io_enq_valid; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_1_io_enq_bits_data; // @[Decoupled.scala 287:21]
  wire [3:0] Queue_1_io_enq_bits_strb; // @[Decoupled.scala 287:21]
  wire  Queue_1_io_enq_bits_last; // @[Decoupled.scala 287:21]
  wire  Queue_1_io_deq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_1_io_deq_valid; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_1_io_deq_bits_data; // @[Decoupled.scala 287:21]
  wire [3:0] Queue_1_io_deq_bits_strb; // @[Decoupled.scala 287:21]
  wire  Queue_1_io_deq_bits_last; // @[Decoupled.scala 287:21]
  wire  Queue_2_clock; // @[Decoupled.scala 287:21]
  wire  Queue_2_reset; // @[Decoupled.scala 287:21]
  wire  Queue_2_io_enq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_2_io_enq_valid; // @[Decoupled.scala 287:21]
  wire  Queue_2_io_enq_bits_id; // @[Decoupled.scala 287:21]
  wire [1:0] Queue_2_io_enq_bits_resp; // @[Decoupled.scala 287:21]
  wire  Queue_2_io_deq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_2_io_deq_valid; // @[Decoupled.scala 287:21]
  wire  Queue_2_io_deq_bits_id; // @[Decoupled.scala 287:21]
  wire [1:0] Queue_2_io_deq_bits_resp; // @[Decoupled.scala 287:21]
  wire  Queue_3_clock; // @[Decoupled.scala 287:21]
  wire  Queue_3_reset; // @[Decoupled.scala 287:21]
  wire  Queue_3_io_enq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_3_io_enq_valid; // @[Decoupled.scala 287:21]
  wire  Queue_3_io_enq_bits_id; // @[Decoupled.scala 287:21]
  wire [29:0] Queue_3_io_enq_bits_addr; // @[Decoupled.scala 287:21]
  wire [2:0] Queue_3_io_enq_bits_size; // @[Decoupled.scala 287:21]
  wire  Queue_3_io_deq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_3_io_deq_valid; // @[Decoupled.scala 287:21]
  wire  Queue_3_io_deq_bits_id; // @[Decoupled.scala 287:21]
  wire [29:0] Queue_3_io_deq_bits_addr; // @[Decoupled.scala 287:21]
  wire [2:0] Queue_3_io_deq_bits_size; // @[Decoupled.scala 287:21]
  wire  Queue_4_clock; // @[Decoupled.scala 287:21]
  wire  Queue_4_reset; // @[Decoupled.scala 287:21]
  wire  Queue_4_io_enq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_4_io_enq_valid; // @[Decoupled.scala 287:21]
  wire  Queue_4_io_enq_bits_id; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_4_io_enq_bits_data; // @[Decoupled.scala 287:21]
  wire [1:0] Queue_4_io_enq_bits_resp; // @[Decoupled.scala 287:21]
  wire  Queue_4_io_enq_bits_last; // @[Decoupled.scala 287:21]
  wire  Queue_4_io_deq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_4_io_deq_valid; // @[Decoupled.scala 287:21]
  wire  Queue_4_io_deq_bits_id; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_4_io_deq_bits_data; // @[Decoupled.scala 287:21]
  wire [1:0] Queue_4_io_deq_bits_resp; // @[Decoupled.scala 287:21]
  wire  Queue_4_io_deq_bits_last; // @[Decoupled.scala 287:21]
  Queue_25 Queue ( // @[Decoupled.scala 287:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_id(Queue_io_enq_bits_id),
    .io_enq_bits_addr(Queue_io_enq_bits_addr),
    .io_enq_bits_size(Queue_io_enq_bits_size),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_id(Queue_io_deq_bits_id),
    .io_deq_bits_addr(Queue_io_deq_bits_addr),
    .io_deq_bits_size(Queue_io_deq_bits_size)
  );
  Queue_26 Queue_1 ( // @[Decoupled.scala 287:21]
    .clock(Queue_1_clock),
    .reset(Queue_1_reset),
    .io_enq_ready(Queue_1_io_enq_ready),
    .io_enq_valid(Queue_1_io_enq_valid),
    .io_enq_bits_data(Queue_1_io_enq_bits_data),
    .io_enq_bits_strb(Queue_1_io_enq_bits_strb),
    .io_enq_bits_last(Queue_1_io_enq_bits_last),
    .io_deq_ready(Queue_1_io_deq_ready),
    .io_deq_valid(Queue_1_io_deq_valid),
    .io_deq_bits_data(Queue_1_io_deq_bits_data),
    .io_deq_bits_strb(Queue_1_io_deq_bits_strb),
    .io_deq_bits_last(Queue_1_io_deq_bits_last)
  );
  Queue_27 Queue_2 ( // @[Decoupled.scala 287:21]
    .clock(Queue_2_clock),
    .reset(Queue_2_reset),
    .io_enq_ready(Queue_2_io_enq_ready),
    .io_enq_valid(Queue_2_io_enq_valid),
    .io_enq_bits_id(Queue_2_io_enq_bits_id),
    .io_enq_bits_resp(Queue_2_io_enq_bits_resp),
    .io_deq_ready(Queue_2_io_deq_ready),
    .io_deq_valid(Queue_2_io_deq_valid),
    .io_deq_bits_id(Queue_2_io_deq_bits_id),
    .io_deq_bits_resp(Queue_2_io_deq_bits_resp)
  );
  Queue_25 Queue_3 ( // @[Decoupled.scala 287:21]
    .clock(Queue_3_clock),
    .reset(Queue_3_reset),
    .io_enq_ready(Queue_3_io_enq_ready),
    .io_enq_valid(Queue_3_io_enq_valid),
    .io_enq_bits_id(Queue_3_io_enq_bits_id),
    .io_enq_bits_addr(Queue_3_io_enq_bits_addr),
    .io_enq_bits_size(Queue_3_io_enq_bits_size),
    .io_deq_ready(Queue_3_io_deq_ready),
    .io_deq_valid(Queue_3_io_deq_valid),
    .io_deq_bits_id(Queue_3_io_deq_bits_id),
    .io_deq_bits_addr(Queue_3_io_deq_bits_addr),
    .io_deq_bits_size(Queue_3_io_deq_bits_size)
  );
  Queue_29 Queue_4 ( // @[Decoupled.scala 287:21]
    .clock(Queue_4_clock),
    .reset(Queue_4_reset),
    .io_enq_ready(Queue_4_io_enq_ready),
    .io_enq_valid(Queue_4_io_enq_valid),
    .io_enq_bits_id(Queue_4_io_enq_bits_id),
    .io_enq_bits_data(Queue_4_io_enq_bits_data),
    .io_enq_bits_resp(Queue_4_io_enq_bits_resp),
    .io_enq_bits_last(Queue_4_io_enq_bits_last),
    .io_deq_ready(Queue_4_io_deq_ready),
    .io_deq_valid(Queue_4_io_deq_valid),
    .io_deq_bits_id(Queue_4_io_deq_bits_id),
    .io_deq_bits_data(Queue_4_io_deq_bits_data),
    .io_deq_bits_resp(Queue_4_io_deq_bits_resp),
    .io_deq_bits_last(Queue_4_io_deq_bits_last)
  );
  assign auto_in_aw_ready = Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_in_w_ready = Queue_1_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_in_b_valid = Queue_2_io_deq_valid; // @[LazyModule.scala 173:31]
  assign auto_in_b_bits_id = Queue_2_io_deq_bits_id; // @[LazyModule.scala 173:31]
  assign auto_in_b_bits_resp = Queue_2_io_deq_bits_resp; // @[LazyModule.scala 173:31]
  assign auto_in_ar_ready = Queue_3_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_in_r_valid = Queue_4_io_deq_valid; // @[LazyModule.scala 173:31]
  assign auto_in_r_bits_id = Queue_4_io_deq_bits_id; // @[LazyModule.scala 173:31]
  assign auto_in_r_bits_data = Queue_4_io_deq_bits_data; // @[LazyModule.scala 173:31]
  assign auto_in_r_bits_resp = Queue_4_io_deq_bits_resp; // @[LazyModule.scala 173:31]
  assign auto_in_r_bits_last = Queue_4_io_deq_bits_last; // @[LazyModule.scala 173:31]
  assign auto_out_aw_valid = Queue_io_deq_valid; // @[LazyModule.scala 173:49]
  assign auto_out_aw_bits_id = Queue_io_deq_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_aw_bits_addr = Queue_io_deq_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_w_valid = Queue_1_io_deq_valid; // @[LazyModule.scala 173:49]
  assign auto_out_w_bits_data = Queue_1_io_deq_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_w_bits_strb = Queue_1_io_deq_bits_strb; // @[LazyModule.scala 173:49]
  assign auto_out_w_bits_last = Queue_1_io_deq_bits_last; // @[LazyModule.scala 173:49]
  assign auto_out_b_ready = Queue_2_io_enq_ready; // @[LazyModule.scala 173:49]
  assign auto_out_ar_valid = Queue_3_io_deq_valid; // @[LazyModule.scala 173:49]
  assign auto_out_ar_bits_id = Queue_3_io_deq_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_ar_bits_addr = Queue_3_io_deq_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_ar_bits_size = Queue_3_io_deq_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_r_ready = Queue_4_io_enq_ready; // @[LazyModule.scala 173:49]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_in_aw_valid; // @[Decoupled.scala 288:22]
  assign Queue_io_enq_bits_id = auto_in_aw_bits_id; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_addr = auto_in_aw_bits_addr; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_size = auto_in_aw_bits_size; // @[Decoupled.scala 289:21]
  assign Queue_io_deq_ready = auto_out_aw_ready; // @[Decoupled.scala 311:15]
  assign Queue_1_clock = clock;
  assign Queue_1_reset = reset;
  assign Queue_1_io_enq_valid = auto_in_w_valid; // @[Decoupled.scala 288:22]
  assign Queue_1_io_enq_bits_data = auto_in_w_bits_data; // @[Decoupled.scala 289:21]
  assign Queue_1_io_enq_bits_strb = auto_in_w_bits_strb; // @[Decoupled.scala 289:21]
  assign Queue_1_io_enq_bits_last = auto_in_w_bits_last; // @[Decoupled.scala 289:21]
  assign Queue_1_io_deq_ready = auto_out_w_ready; // @[Decoupled.scala 311:15]
  assign Queue_2_clock = clock;
  assign Queue_2_reset = reset;
  assign Queue_2_io_enq_valid = auto_out_b_valid; // @[Decoupled.scala 288:22]
  assign Queue_2_io_enq_bits_id = auto_out_b_bits_id; // @[Decoupled.scala 289:21]
  assign Queue_2_io_enq_bits_resp = auto_out_b_bits_resp; // @[Decoupled.scala 289:21]
  assign Queue_2_io_deq_ready = auto_in_b_ready; // @[Decoupled.scala 311:15]
  assign Queue_3_clock = clock;
  assign Queue_3_reset = reset;
  assign Queue_3_io_enq_valid = auto_in_ar_valid; // @[Decoupled.scala 288:22]
  assign Queue_3_io_enq_bits_id = auto_in_ar_bits_id; // @[Decoupled.scala 289:21]
  assign Queue_3_io_enq_bits_addr = auto_in_ar_bits_addr; // @[Decoupled.scala 289:21]
  assign Queue_3_io_enq_bits_size = auto_in_ar_bits_size; // @[Decoupled.scala 289:21]
  assign Queue_3_io_deq_ready = auto_out_ar_ready; // @[Decoupled.scala 311:15]
  assign Queue_4_clock = clock;
  assign Queue_4_reset = reset;
  assign Queue_4_io_enq_valid = auto_out_r_valid; // @[Decoupled.scala 288:22]
  assign Queue_4_io_enq_bits_id = auto_out_r_bits_id; // @[Decoupled.scala 289:21]
  assign Queue_4_io_enq_bits_data = auto_out_r_bits_data; // @[Decoupled.scala 289:21]
  assign Queue_4_io_enq_bits_resp = auto_out_r_bits_resp; // @[Decoupled.scala 289:21]
  assign Queue_4_io_enq_bits_last = auto_out_r_bits_last; // @[Decoupled.scala 289:21]
  assign Queue_4_io_deq_ready = auto_in_r_ready; // @[Decoupled.scala 311:15]
endmodule
module AccumulatorChain(
  input         clock,
  input         reset,
  output        auto_bus_in_aw_ready,
  input         auto_bus_in_aw_valid,
  input         auto_bus_in_aw_bits_id,
  input  [29:0] auto_bus_in_aw_bits_addr,
  input  [2:0]  auto_bus_in_aw_bits_size,
  output        auto_bus_in_w_ready,
  input         auto_bus_in_w_valid,
  input  [31:0] auto_bus_in_w_bits_data,
  input  [3:0]  auto_bus_in_w_bits_strb,
  input         auto_bus_in_w_bits_last,
  input         auto_bus_in_b_ready,
  output        auto_bus_in_b_valid,
  output [1:0]  auto_bus_in_b_bits_resp,
  output        auto_bus_in_ar_ready,
  input         auto_bus_in_ar_valid,
  input         auto_bus_in_ar_bits_id,
  input  [29:0] auto_bus_in_ar_bits_addr,
  input  [2:0]  auto_bus_in_ar_bits_size,
  input         auto_bus_in_r_ready,
  output        auto_bus_in_r_valid,
  output [31:0] auto_bus_in_r_bits_data,
  output [1:0]  auto_bus_in_r_bits_resp,
  output        auto_bus_in_r_bits_last,
  input         auto_dspQueue_stream_out_ready,
  output        auto_dspQueue_stream_out_valid,
  output [15:0] auto_dspQueue_stream_out_bits_data,
  output        auto_dspQueue_stream_out_bits_last,
  output        auto_accumulator_slave_in_ready,
  input         auto_accumulator_slave_in_valid,
  input  [31:0] auto_accumulator_slave_in_bits_data,
  input         auto_accumulator_slave_in_bits_last
);
  wire  accumulator_clock; // @[AccChain.scala 27:30]
  wire  accumulator_reset; // @[AccChain.scala 27:30]
  wire  accumulator_auto_mem_in_aw_ready; // @[AccChain.scala 27:30]
  wire  accumulator_auto_mem_in_aw_valid; // @[AccChain.scala 27:30]
  wire  accumulator_auto_mem_in_aw_bits_id; // @[AccChain.scala 27:30]
  wire [29:0] accumulator_auto_mem_in_aw_bits_addr; // @[AccChain.scala 27:30]
  wire  accumulator_auto_mem_in_w_ready; // @[AccChain.scala 27:30]
  wire  accumulator_auto_mem_in_w_valid; // @[AccChain.scala 27:30]
  wire [31:0] accumulator_auto_mem_in_w_bits_data; // @[AccChain.scala 27:30]
  wire [3:0] accumulator_auto_mem_in_w_bits_strb; // @[AccChain.scala 27:30]
  wire  accumulator_auto_mem_in_b_ready; // @[AccChain.scala 27:30]
  wire  accumulator_auto_mem_in_b_valid; // @[AccChain.scala 27:30]
  wire  accumulator_auto_mem_in_b_bits_id; // @[AccChain.scala 27:30]
  wire  accumulator_auto_mem_in_ar_ready; // @[AccChain.scala 27:30]
  wire  accumulator_auto_mem_in_ar_valid; // @[AccChain.scala 27:30]
  wire  accumulator_auto_mem_in_ar_bits_id; // @[AccChain.scala 27:30]
  wire [29:0] accumulator_auto_mem_in_ar_bits_addr; // @[AccChain.scala 27:30]
  wire [2:0] accumulator_auto_mem_in_ar_bits_size; // @[AccChain.scala 27:30]
  wire  accumulator_auto_mem_in_r_ready; // @[AccChain.scala 27:30]
  wire  accumulator_auto_mem_in_r_valid; // @[AccChain.scala 27:30]
  wire  accumulator_auto_mem_in_r_bits_id; // @[AccChain.scala 27:30]
  wire [31:0] accumulator_auto_mem_in_r_bits_data; // @[AccChain.scala 27:30]
  wire  accumulator_auto_master_out_ready; // @[AccChain.scala 27:30]
  wire  accumulator_auto_master_out_valid; // @[AccChain.scala 27:30]
  wire [15:0] accumulator_auto_master_out_bits_data; // @[AccChain.scala 27:30]
  wire  accumulator_auto_master_out_bits_last; // @[AccChain.scala 27:30]
  wire  accumulator_auto_slave_in_ready; // @[AccChain.scala 27:30]
  wire  accumulator_auto_slave_in_valid; // @[AccChain.scala 27:30]
  wire [31:0] accumulator_auto_slave_in_bits_data; // @[AccChain.scala 27:30]
  wire  accumulator_auto_slave_in_bits_last; // @[AccChain.scala 27:30]
  wire  dspQueue_clock; // @[AccChain.scala 29:27]
  wire  dspQueue_reset; // @[AccChain.scala 29:27]
  wire  dspQueue_auto_stream_in_ready; // @[AccChain.scala 29:27]
  wire  dspQueue_auto_stream_in_valid; // @[AccChain.scala 29:27]
  wire [15:0] dspQueue_auto_stream_in_bits_data; // @[AccChain.scala 29:27]
  wire  dspQueue_auto_stream_in_bits_last; // @[AccChain.scala 29:27]
  wire  dspQueue_auto_stream_out_ready; // @[AccChain.scala 29:27]
  wire  dspQueue_auto_stream_out_valid; // @[AccChain.scala 29:27]
  wire [15:0] dspQueue_auto_stream_out_bits_data; // @[AccChain.scala 29:27]
  wire  dspQueue_auto_stream_out_bits_last; // @[AccChain.scala 29:27]
  wire  dspQueue_auto_in_aw_ready; // @[AccChain.scala 29:27]
  wire  dspQueue_auto_in_aw_valid; // @[AccChain.scala 29:27]
  wire  dspQueue_auto_in_aw_bits_id; // @[AccChain.scala 29:27]
  wire [29:0] dspQueue_auto_in_aw_bits_addr; // @[AccChain.scala 29:27]
  wire  dspQueue_auto_in_w_ready; // @[AccChain.scala 29:27]
  wire  dspQueue_auto_in_w_valid; // @[AccChain.scala 29:27]
  wire [31:0] dspQueue_auto_in_w_bits_data; // @[AccChain.scala 29:27]
  wire [3:0] dspQueue_auto_in_w_bits_strb; // @[AccChain.scala 29:27]
  wire  dspQueue_auto_in_b_ready; // @[AccChain.scala 29:27]
  wire  dspQueue_auto_in_b_valid; // @[AccChain.scala 29:27]
  wire  dspQueue_auto_in_b_bits_id; // @[AccChain.scala 29:27]
  wire  dspQueue_auto_in_ar_ready; // @[AccChain.scala 29:27]
  wire  dspQueue_auto_in_ar_valid; // @[AccChain.scala 29:27]
  wire  dspQueue_auto_in_ar_bits_id; // @[AccChain.scala 29:27]
  wire [29:0] dspQueue_auto_in_ar_bits_addr; // @[AccChain.scala 29:27]
  wire [2:0] dspQueue_auto_in_ar_bits_size; // @[AccChain.scala 29:27]
  wire  dspQueue_auto_in_r_ready; // @[AccChain.scala 29:27]
  wire  dspQueue_auto_in_r_valid; // @[AccChain.scala 29:27]
  wire  dspQueue_auto_in_r_bits_id; // @[AccChain.scala 29:27]
  wire [31:0] dspQueue_auto_in_r_bits_data; // @[AccChain.scala 29:27]
  wire  bus_clock; // @[AccChain.scala 44:23]
  wire  bus_reset; // @[AccChain.scala 44:23]
  wire  bus_auto_in_aw_ready; // @[AccChain.scala 44:23]
  wire  bus_auto_in_aw_valid; // @[AccChain.scala 44:23]
  wire  bus_auto_in_aw_bits_id; // @[AccChain.scala 44:23]
  wire [29:0] bus_auto_in_aw_bits_addr; // @[AccChain.scala 44:23]
  wire [2:0] bus_auto_in_aw_bits_size; // @[AccChain.scala 44:23]
  wire  bus_auto_in_w_ready; // @[AccChain.scala 44:23]
  wire  bus_auto_in_w_valid; // @[AccChain.scala 44:23]
  wire [31:0] bus_auto_in_w_bits_data; // @[AccChain.scala 44:23]
  wire [3:0] bus_auto_in_w_bits_strb; // @[AccChain.scala 44:23]
  wire  bus_auto_in_w_bits_last; // @[AccChain.scala 44:23]
  wire  bus_auto_in_b_ready; // @[AccChain.scala 44:23]
  wire  bus_auto_in_b_valid; // @[AccChain.scala 44:23]
  wire [1:0] bus_auto_in_b_bits_resp; // @[AccChain.scala 44:23]
  wire  bus_auto_in_ar_ready; // @[AccChain.scala 44:23]
  wire  bus_auto_in_ar_valid; // @[AccChain.scala 44:23]
  wire  bus_auto_in_ar_bits_id; // @[AccChain.scala 44:23]
  wire [29:0] bus_auto_in_ar_bits_addr; // @[AccChain.scala 44:23]
  wire [2:0] bus_auto_in_ar_bits_size; // @[AccChain.scala 44:23]
  wire  bus_auto_in_r_ready; // @[AccChain.scala 44:23]
  wire  bus_auto_in_r_valid; // @[AccChain.scala 44:23]
  wire [31:0] bus_auto_in_r_bits_data; // @[AccChain.scala 44:23]
  wire [1:0] bus_auto_in_r_bits_resp; // @[AccChain.scala 44:23]
  wire  bus_auto_in_r_bits_last; // @[AccChain.scala 44:23]
  wire  bus_auto_out_1_aw_ready; // @[AccChain.scala 44:23]
  wire  bus_auto_out_1_aw_valid; // @[AccChain.scala 44:23]
  wire  bus_auto_out_1_aw_bits_id; // @[AccChain.scala 44:23]
  wire [29:0] bus_auto_out_1_aw_bits_addr; // @[AccChain.scala 44:23]
  wire [2:0] bus_auto_out_1_aw_bits_size; // @[AccChain.scala 44:23]
  wire  bus_auto_out_1_w_ready; // @[AccChain.scala 44:23]
  wire  bus_auto_out_1_w_valid; // @[AccChain.scala 44:23]
  wire [31:0] bus_auto_out_1_w_bits_data; // @[AccChain.scala 44:23]
  wire [3:0] bus_auto_out_1_w_bits_strb; // @[AccChain.scala 44:23]
  wire  bus_auto_out_1_w_bits_last; // @[AccChain.scala 44:23]
  wire  bus_auto_out_1_b_ready; // @[AccChain.scala 44:23]
  wire  bus_auto_out_1_b_valid; // @[AccChain.scala 44:23]
  wire  bus_auto_out_1_b_bits_id; // @[AccChain.scala 44:23]
  wire [1:0] bus_auto_out_1_b_bits_resp; // @[AccChain.scala 44:23]
  wire  bus_auto_out_1_ar_ready; // @[AccChain.scala 44:23]
  wire  bus_auto_out_1_ar_valid; // @[AccChain.scala 44:23]
  wire  bus_auto_out_1_ar_bits_id; // @[AccChain.scala 44:23]
  wire [29:0] bus_auto_out_1_ar_bits_addr; // @[AccChain.scala 44:23]
  wire [2:0] bus_auto_out_1_ar_bits_size; // @[AccChain.scala 44:23]
  wire  bus_auto_out_1_r_ready; // @[AccChain.scala 44:23]
  wire  bus_auto_out_1_r_valid; // @[AccChain.scala 44:23]
  wire  bus_auto_out_1_r_bits_id; // @[AccChain.scala 44:23]
  wire [31:0] bus_auto_out_1_r_bits_data; // @[AccChain.scala 44:23]
  wire [1:0] bus_auto_out_1_r_bits_resp; // @[AccChain.scala 44:23]
  wire  bus_auto_out_1_r_bits_last; // @[AccChain.scala 44:23]
  wire  bus_auto_out_0_aw_ready; // @[AccChain.scala 44:23]
  wire  bus_auto_out_0_aw_valid; // @[AccChain.scala 44:23]
  wire  bus_auto_out_0_aw_bits_id; // @[AccChain.scala 44:23]
  wire [29:0] bus_auto_out_0_aw_bits_addr; // @[AccChain.scala 44:23]
  wire [2:0] bus_auto_out_0_aw_bits_size; // @[AccChain.scala 44:23]
  wire  bus_auto_out_0_w_ready; // @[AccChain.scala 44:23]
  wire  bus_auto_out_0_w_valid; // @[AccChain.scala 44:23]
  wire [31:0] bus_auto_out_0_w_bits_data; // @[AccChain.scala 44:23]
  wire [3:0] bus_auto_out_0_w_bits_strb; // @[AccChain.scala 44:23]
  wire  bus_auto_out_0_w_bits_last; // @[AccChain.scala 44:23]
  wire  bus_auto_out_0_b_ready; // @[AccChain.scala 44:23]
  wire  bus_auto_out_0_b_valid; // @[AccChain.scala 44:23]
  wire  bus_auto_out_0_b_bits_id; // @[AccChain.scala 44:23]
  wire [1:0] bus_auto_out_0_b_bits_resp; // @[AccChain.scala 44:23]
  wire  bus_auto_out_0_ar_ready; // @[AccChain.scala 44:23]
  wire  bus_auto_out_0_ar_valid; // @[AccChain.scala 44:23]
  wire  bus_auto_out_0_ar_bits_id; // @[AccChain.scala 44:23]
  wire [29:0] bus_auto_out_0_ar_bits_addr; // @[AccChain.scala 44:23]
  wire [2:0] bus_auto_out_0_ar_bits_size; // @[AccChain.scala 44:23]
  wire  bus_auto_out_0_r_ready; // @[AccChain.scala 44:23]
  wire  bus_auto_out_0_r_valid; // @[AccChain.scala 44:23]
  wire  bus_auto_out_0_r_bits_id; // @[AccChain.scala 44:23]
  wire [31:0] bus_auto_out_0_r_bits_data; // @[AccChain.scala 44:23]
  wire [1:0] bus_auto_out_0_r_bits_resp; // @[AccChain.scala 44:23]
  wire  bus_auto_out_0_r_bits_last; // @[AccChain.scala 44:23]
  wire  axi4buf_clock; // @[Buffer.scala 58:29]
  wire  axi4buf_reset; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_in_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_in_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_in_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_auto_in_aw_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_auto_in_aw_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_in_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_in_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_auto_in_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_auto_in_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_in_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_in_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_in_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_in_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_auto_in_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_in_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_in_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_in_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_auto_in_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_auto_in_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_in_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_in_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_in_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_auto_in_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_auto_in_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_in_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_out_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_out_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_out_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_auto_out_aw_bits_addr; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_out_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_out_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_auto_out_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_auto_out_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_out_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_out_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_out_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_out_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_auto_out_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_out_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_out_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_out_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_auto_out_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_auto_out_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_out_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_out_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_out_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_auto_out_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_auto_out_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_out_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_1_clock; // @[Buffer.scala 58:29]
  wire  axi4buf_1_reset; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_in_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_in_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_in_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_1_auto_in_aw_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_1_auto_in_aw_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_in_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_in_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_1_auto_in_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_1_auto_in_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_in_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_in_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_in_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_in_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_1_auto_in_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_in_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_in_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_in_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_1_auto_in_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_1_auto_in_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_in_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_in_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_in_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_1_auto_in_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_1_auto_in_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_in_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_out_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_out_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_out_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_1_auto_out_aw_bits_addr; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_out_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_out_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_1_auto_out_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_1_auto_out_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_out_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_out_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_out_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_out_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_1_auto_out_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_out_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_out_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_out_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_1_auto_out_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_1_auto_out_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_out_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_out_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_out_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_1_auto_out_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_1_auto_out_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_out_r_bits_last; // @[Buffer.scala 58:29]
  AXI4AccumulatorBlock accumulator ( // @[AccChain.scala 27:30]
    .clock(accumulator_clock),
    .reset(accumulator_reset),
    .auto_mem_in_aw_ready(accumulator_auto_mem_in_aw_ready),
    .auto_mem_in_aw_valid(accumulator_auto_mem_in_aw_valid),
    .auto_mem_in_aw_bits_id(accumulator_auto_mem_in_aw_bits_id),
    .auto_mem_in_aw_bits_addr(accumulator_auto_mem_in_aw_bits_addr),
    .auto_mem_in_w_ready(accumulator_auto_mem_in_w_ready),
    .auto_mem_in_w_valid(accumulator_auto_mem_in_w_valid),
    .auto_mem_in_w_bits_data(accumulator_auto_mem_in_w_bits_data),
    .auto_mem_in_w_bits_strb(accumulator_auto_mem_in_w_bits_strb),
    .auto_mem_in_b_ready(accumulator_auto_mem_in_b_ready),
    .auto_mem_in_b_valid(accumulator_auto_mem_in_b_valid),
    .auto_mem_in_b_bits_id(accumulator_auto_mem_in_b_bits_id),
    .auto_mem_in_ar_ready(accumulator_auto_mem_in_ar_ready),
    .auto_mem_in_ar_valid(accumulator_auto_mem_in_ar_valid),
    .auto_mem_in_ar_bits_id(accumulator_auto_mem_in_ar_bits_id),
    .auto_mem_in_ar_bits_addr(accumulator_auto_mem_in_ar_bits_addr),
    .auto_mem_in_ar_bits_size(accumulator_auto_mem_in_ar_bits_size),
    .auto_mem_in_r_ready(accumulator_auto_mem_in_r_ready),
    .auto_mem_in_r_valid(accumulator_auto_mem_in_r_valid),
    .auto_mem_in_r_bits_id(accumulator_auto_mem_in_r_bits_id),
    .auto_mem_in_r_bits_data(accumulator_auto_mem_in_r_bits_data),
    .auto_master_out_ready(accumulator_auto_master_out_ready),
    .auto_master_out_valid(accumulator_auto_master_out_valid),
    .auto_master_out_bits_data(accumulator_auto_master_out_bits_data),
    .auto_master_out_bits_last(accumulator_auto_master_out_bits_last),
    .auto_slave_in_ready(accumulator_auto_slave_in_ready),
    .auto_slave_in_valid(accumulator_auto_slave_in_valid),
    .auto_slave_in_bits_data(accumulator_auto_slave_in_bits_data),
    .auto_slave_in_bits_last(accumulator_auto_slave_in_bits_last)
  );
  AXI4DspQueueBlock dspQueue ( // @[AccChain.scala 29:27]
    .clock(dspQueue_clock),
    .reset(dspQueue_reset),
    .auto_stream_in_ready(dspQueue_auto_stream_in_ready),
    .auto_stream_in_valid(dspQueue_auto_stream_in_valid),
    .auto_stream_in_bits_data(dspQueue_auto_stream_in_bits_data),
    .auto_stream_in_bits_last(dspQueue_auto_stream_in_bits_last),
    .auto_stream_out_ready(dspQueue_auto_stream_out_ready),
    .auto_stream_out_valid(dspQueue_auto_stream_out_valid),
    .auto_stream_out_bits_data(dspQueue_auto_stream_out_bits_data),
    .auto_stream_out_bits_last(dspQueue_auto_stream_out_bits_last),
    .auto_in_aw_ready(dspQueue_auto_in_aw_ready),
    .auto_in_aw_valid(dspQueue_auto_in_aw_valid),
    .auto_in_aw_bits_id(dspQueue_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(dspQueue_auto_in_aw_bits_addr),
    .auto_in_w_ready(dspQueue_auto_in_w_ready),
    .auto_in_w_valid(dspQueue_auto_in_w_valid),
    .auto_in_w_bits_data(dspQueue_auto_in_w_bits_data),
    .auto_in_w_bits_strb(dspQueue_auto_in_w_bits_strb),
    .auto_in_b_ready(dspQueue_auto_in_b_ready),
    .auto_in_b_valid(dspQueue_auto_in_b_valid),
    .auto_in_b_bits_id(dspQueue_auto_in_b_bits_id),
    .auto_in_ar_ready(dspQueue_auto_in_ar_ready),
    .auto_in_ar_valid(dspQueue_auto_in_ar_valid),
    .auto_in_ar_bits_id(dspQueue_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(dspQueue_auto_in_ar_bits_addr),
    .auto_in_ar_bits_size(dspQueue_auto_in_ar_bits_size),
    .auto_in_r_ready(dspQueue_auto_in_r_ready),
    .auto_in_r_valid(dspQueue_auto_in_r_valid),
    .auto_in_r_bits_id(dspQueue_auto_in_r_bits_id),
    .auto_in_r_bits_data(dspQueue_auto_in_r_bits_data)
  );
  AXI4Xbar_1 bus ( // @[AccChain.scala 44:23]
    .clock(bus_clock),
    .reset(bus_reset),
    .auto_in_aw_ready(bus_auto_in_aw_ready),
    .auto_in_aw_valid(bus_auto_in_aw_valid),
    .auto_in_aw_bits_id(bus_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(bus_auto_in_aw_bits_addr),
    .auto_in_aw_bits_size(bus_auto_in_aw_bits_size),
    .auto_in_w_ready(bus_auto_in_w_ready),
    .auto_in_w_valid(bus_auto_in_w_valid),
    .auto_in_w_bits_data(bus_auto_in_w_bits_data),
    .auto_in_w_bits_strb(bus_auto_in_w_bits_strb),
    .auto_in_w_bits_last(bus_auto_in_w_bits_last),
    .auto_in_b_ready(bus_auto_in_b_ready),
    .auto_in_b_valid(bus_auto_in_b_valid),
    .auto_in_b_bits_resp(bus_auto_in_b_bits_resp),
    .auto_in_ar_ready(bus_auto_in_ar_ready),
    .auto_in_ar_valid(bus_auto_in_ar_valid),
    .auto_in_ar_bits_id(bus_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(bus_auto_in_ar_bits_addr),
    .auto_in_ar_bits_size(bus_auto_in_ar_bits_size),
    .auto_in_r_ready(bus_auto_in_r_ready),
    .auto_in_r_valid(bus_auto_in_r_valid),
    .auto_in_r_bits_data(bus_auto_in_r_bits_data),
    .auto_in_r_bits_resp(bus_auto_in_r_bits_resp),
    .auto_in_r_bits_last(bus_auto_in_r_bits_last),
    .auto_out_1_aw_ready(bus_auto_out_1_aw_ready),
    .auto_out_1_aw_valid(bus_auto_out_1_aw_valid),
    .auto_out_1_aw_bits_id(bus_auto_out_1_aw_bits_id),
    .auto_out_1_aw_bits_addr(bus_auto_out_1_aw_bits_addr),
    .auto_out_1_aw_bits_size(bus_auto_out_1_aw_bits_size),
    .auto_out_1_w_ready(bus_auto_out_1_w_ready),
    .auto_out_1_w_valid(bus_auto_out_1_w_valid),
    .auto_out_1_w_bits_data(bus_auto_out_1_w_bits_data),
    .auto_out_1_w_bits_strb(bus_auto_out_1_w_bits_strb),
    .auto_out_1_w_bits_last(bus_auto_out_1_w_bits_last),
    .auto_out_1_b_ready(bus_auto_out_1_b_ready),
    .auto_out_1_b_valid(bus_auto_out_1_b_valid),
    .auto_out_1_b_bits_id(bus_auto_out_1_b_bits_id),
    .auto_out_1_b_bits_resp(bus_auto_out_1_b_bits_resp),
    .auto_out_1_ar_ready(bus_auto_out_1_ar_ready),
    .auto_out_1_ar_valid(bus_auto_out_1_ar_valid),
    .auto_out_1_ar_bits_id(bus_auto_out_1_ar_bits_id),
    .auto_out_1_ar_bits_addr(bus_auto_out_1_ar_bits_addr),
    .auto_out_1_ar_bits_size(bus_auto_out_1_ar_bits_size),
    .auto_out_1_r_ready(bus_auto_out_1_r_ready),
    .auto_out_1_r_valid(bus_auto_out_1_r_valid),
    .auto_out_1_r_bits_id(bus_auto_out_1_r_bits_id),
    .auto_out_1_r_bits_data(bus_auto_out_1_r_bits_data),
    .auto_out_1_r_bits_resp(bus_auto_out_1_r_bits_resp),
    .auto_out_1_r_bits_last(bus_auto_out_1_r_bits_last),
    .auto_out_0_aw_ready(bus_auto_out_0_aw_ready),
    .auto_out_0_aw_valid(bus_auto_out_0_aw_valid),
    .auto_out_0_aw_bits_id(bus_auto_out_0_aw_bits_id),
    .auto_out_0_aw_bits_addr(bus_auto_out_0_aw_bits_addr),
    .auto_out_0_aw_bits_size(bus_auto_out_0_aw_bits_size),
    .auto_out_0_w_ready(bus_auto_out_0_w_ready),
    .auto_out_0_w_valid(bus_auto_out_0_w_valid),
    .auto_out_0_w_bits_data(bus_auto_out_0_w_bits_data),
    .auto_out_0_w_bits_strb(bus_auto_out_0_w_bits_strb),
    .auto_out_0_w_bits_last(bus_auto_out_0_w_bits_last),
    .auto_out_0_b_ready(bus_auto_out_0_b_ready),
    .auto_out_0_b_valid(bus_auto_out_0_b_valid),
    .auto_out_0_b_bits_id(bus_auto_out_0_b_bits_id),
    .auto_out_0_b_bits_resp(bus_auto_out_0_b_bits_resp),
    .auto_out_0_ar_ready(bus_auto_out_0_ar_ready),
    .auto_out_0_ar_valid(bus_auto_out_0_ar_valid),
    .auto_out_0_ar_bits_id(bus_auto_out_0_ar_bits_id),
    .auto_out_0_ar_bits_addr(bus_auto_out_0_ar_bits_addr),
    .auto_out_0_ar_bits_size(bus_auto_out_0_ar_bits_size),
    .auto_out_0_r_ready(bus_auto_out_0_r_ready),
    .auto_out_0_r_valid(bus_auto_out_0_r_valid),
    .auto_out_0_r_bits_id(bus_auto_out_0_r_bits_id),
    .auto_out_0_r_bits_data(bus_auto_out_0_r_bits_data),
    .auto_out_0_r_bits_resp(bus_auto_out_0_r_bits_resp),
    .auto_out_0_r_bits_last(bus_auto_out_0_r_bits_last)
  );
  AXI4Buffer axi4buf ( // @[Buffer.scala 58:29]
    .clock(axi4buf_clock),
    .reset(axi4buf_reset),
    .auto_in_aw_ready(axi4buf_auto_in_aw_ready),
    .auto_in_aw_valid(axi4buf_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4buf_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4buf_auto_in_aw_bits_addr),
    .auto_in_aw_bits_size(axi4buf_auto_in_aw_bits_size),
    .auto_in_w_ready(axi4buf_auto_in_w_ready),
    .auto_in_w_valid(axi4buf_auto_in_w_valid),
    .auto_in_w_bits_data(axi4buf_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi4buf_auto_in_w_bits_strb),
    .auto_in_w_bits_last(axi4buf_auto_in_w_bits_last),
    .auto_in_b_ready(axi4buf_auto_in_b_ready),
    .auto_in_b_valid(axi4buf_auto_in_b_valid),
    .auto_in_b_bits_id(axi4buf_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi4buf_auto_in_b_bits_resp),
    .auto_in_ar_ready(axi4buf_auto_in_ar_ready),
    .auto_in_ar_valid(axi4buf_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4buf_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4buf_auto_in_ar_bits_addr),
    .auto_in_ar_bits_size(axi4buf_auto_in_ar_bits_size),
    .auto_in_r_ready(axi4buf_auto_in_r_ready),
    .auto_in_r_valid(axi4buf_auto_in_r_valid),
    .auto_in_r_bits_id(axi4buf_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4buf_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4buf_auto_in_r_bits_resp),
    .auto_in_r_bits_last(axi4buf_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4buf_auto_out_aw_ready),
    .auto_out_aw_valid(axi4buf_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4buf_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4buf_auto_out_aw_bits_addr),
    .auto_out_w_ready(axi4buf_auto_out_w_ready),
    .auto_out_w_valid(axi4buf_auto_out_w_valid),
    .auto_out_w_bits_data(axi4buf_auto_out_w_bits_data),
    .auto_out_w_bits_strb(axi4buf_auto_out_w_bits_strb),
    .auto_out_w_bits_last(axi4buf_auto_out_w_bits_last),
    .auto_out_b_ready(axi4buf_auto_out_b_ready),
    .auto_out_b_valid(axi4buf_auto_out_b_valid),
    .auto_out_b_bits_id(axi4buf_auto_out_b_bits_id),
    .auto_out_b_bits_resp(axi4buf_auto_out_b_bits_resp),
    .auto_out_ar_ready(axi4buf_auto_out_ar_ready),
    .auto_out_ar_valid(axi4buf_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4buf_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4buf_auto_out_ar_bits_addr),
    .auto_out_ar_bits_size(axi4buf_auto_out_ar_bits_size),
    .auto_out_r_ready(axi4buf_auto_out_r_ready),
    .auto_out_r_valid(axi4buf_auto_out_r_valid),
    .auto_out_r_bits_id(axi4buf_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4buf_auto_out_r_bits_data),
    .auto_out_r_bits_resp(axi4buf_auto_out_r_bits_resp),
    .auto_out_r_bits_last(axi4buf_auto_out_r_bits_last)
  );
  AXI4Buffer axi4buf_1 ( // @[Buffer.scala 58:29]
    .clock(axi4buf_1_clock),
    .reset(axi4buf_1_reset),
    .auto_in_aw_ready(axi4buf_1_auto_in_aw_ready),
    .auto_in_aw_valid(axi4buf_1_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4buf_1_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4buf_1_auto_in_aw_bits_addr),
    .auto_in_aw_bits_size(axi4buf_1_auto_in_aw_bits_size),
    .auto_in_w_ready(axi4buf_1_auto_in_w_ready),
    .auto_in_w_valid(axi4buf_1_auto_in_w_valid),
    .auto_in_w_bits_data(axi4buf_1_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi4buf_1_auto_in_w_bits_strb),
    .auto_in_w_bits_last(axi4buf_1_auto_in_w_bits_last),
    .auto_in_b_ready(axi4buf_1_auto_in_b_ready),
    .auto_in_b_valid(axi4buf_1_auto_in_b_valid),
    .auto_in_b_bits_id(axi4buf_1_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi4buf_1_auto_in_b_bits_resp),
    .auto_in_ar_ready(axi4buf_1_auto_in_ar_ready),
    .auto_in_ar_valid(axi4buf_1_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4buf_1_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4buf_1_auto_in_ar_bits_addr),
    .auto_in_ar_bits_size(axi4buf_1_auto_in_ar_bits_size),
    .auto_in_r_ready(axi4buf_1_auto_in_r_ready),
    .auto_in_r_valid(axi4buf_1_auto_in_r_valid),
    .auto_in_r_bits_id(axi4buf_1_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4buf_1_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4buf_1_auto_in_r_bits_resp),
    .auto_in_r_bits_last(axi4buf_1_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4buf_1_auto_out_aw_ready),
    .auto_out_aw_valid(axi4buf_1_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4buf_1_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4buf_1_auto_out_aw_bits_addr),
    .auto_out_w_ready(axi4buf_1_auto_out_w_ready),
    .auto_out_w_valid(axi4buf_1_auto_out_w_valid),
    .auto_out_w_bits_data(axi4buf_1_auto_out_w_bits_data),
    .auto_out_w_bits_strb(axi4buf_1_auto_out_w_bits_strb),
    .auto_out_w_bits_last(axi4buf_1_auto_out_w_bits_last),
    .auto_out_b_ready(axi4buf_1_auto_out_b_ready),
    .auto_out_b_valid(axi4buf_1_auto_out_b_valid),
    .auto_out_b_bits_id(axi4buf_1_auto_out_b_bits_id),
    .auto_out_b_bits_resp(axi4buf_1_auto_out_b_bits_resp),
    .auto_out_ar_ready(axi4buf_1_auto_out_ar_ready),
    .auto_out_ar_valid(axi4buf_1_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4buf_1_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4buf_1_auto_out_ar_bits_addr),
    .auto_out_ar_bits_size(axi4buf_1_auto_out_ar_bits_size),
    .auto_out_r_ready(axi4buf_1_auto_out_r_ready),
    .auto_out_r_valid(axi4buf_1_auto_out_r_valid),
    .auto_out_r_bits_id(axi4buf_1_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4buf_1_auto_out_r_bits_data),
    .auto_out_r_bits_resp(axi4buf_1_auto_out_r_bits_resp),
    .auto_out_r_bits_last(axi4buf_1_auto_out_r_bits_last)
  );
  assign auto_bus_in_aw_ready = bus_auto_in_aw_ready; // @[LazyModule.scala 173:31]
  assign auto_bus_in_w_ready = bus_auto_in_w_ready; // @[LazyModule.scala 173:31]
  assign auto_bus_in_b_valid = bus_auto_in_b_valid; // @[LazyModule.scala 173:31]
  assign auto_bus_in_b_bits_resp = bus_auto_in_b_bits_resp; // @[LazyModule.scala 173:31]
  assign auto_bus_in_ar_ready = bus_auto_in_ar_ready; // @[LazyModule.scala 173:31]
  assign auto_bus_in_r_valid = bus_auto_in_r_valid; // @[LazyModule.scala 173:31]
  assign auto_bus_in_r_bits_data = bus_auto_in_r_bits_data; // @[LazyModule.scala 173:31]
  assign auto_bus_in_r_bits_resp = bus_auto_in_r_bits_resp; // @[LazyModule.scala 173:31]
  assign auto_bus_in_r_bits_last = bus_auto_in_r_bits_last; // @[LazyModule.scala 173:31]
  assign auto_dspQueue_stream_out_valid = dspQueue_auto_stream_out_valid; // @[LazyModule.scala 173:49]
  assign auto_dspQueue_stream_out_bits_data = dspQueue_auto_stream_out_bits_data; // @[LazyModule.scala 173:49]
  assign auto_dspQueue_stream_out_bits_last = dspQueue_auto_stream_out_bits_last; // @[LazyModule.scala 173:49]
  assign auto_accumulator_slave_in_ready = accumulator_auto_slave_in_ready; // @[LazyModule.scala 173:31]
  assign accumulator_clock = clock;
  assign accumulator_reset = reset;
  assign accumulator_auto_mem_in_aw_valid = axi4buf_1_auto_out_aw_valid; // @[LazyModule.scala 167:31]
  assign accumulator_auto_mem_in_aw_bits_id = axi4buf_1_auto_out_aw_bits_id; // @[LazyModule.scala 167:31]
  assign accumulator_auto_mem_in_aw_bits_addr = axi4buf_1_auto_out_aw_bits_addr; // @[LazyModule.scala 167:31]
  assign accumulator_auto_mem_in_w_valid = axi4buf_1_auto_out_w_valid; // @[LazyModule.scala 167:31]
  assign accumulator_auto_mem_in_w_bits_data = axi4buf_1_auto_out_w_bits_data; // @[LazyModule.scala 167:31]
  assign accumulator_auto_mem_in_w_bits_strb = axi4buf_1_auto_out_w_bits_strb; // @[LazyModule.scala 167:31]
  assign accumulator_auto_mem_in_b_ready = axi4buf_1_auto_out_b_ready; // @[LazyModule.scala 167:31]
  assign accumulator_auto_mem_in_ar_valid = axi4buf_1_auto_out_ar_valid; // @[LazyModule.scala 167:31]
  assign accumulator_auto_mem_in_ar_bits_id = axi4buf_1_auto_out_ar_bits_id; // @[LazyModule.scala 167:31]
  assign accumulator_auto_mem_in_ar_bits_addr = axi4buf_1_auto_out_ar_bits_addr; // @[LazyModule.scala 167:31]
  assign accumulator_auto_mem_in_ar_bits_size = axi4buf_1_auto_out_ar_bits_size; // @[LazyModule.scala 167:31]
  assign accumulator_auto_mem_in_r_ready = axi4buf_1_auto_out_r_ready; // @[LazyModule.scala 167:31]
  assign accumulator_auto_master_out_ready = dspQueue_auto_stream_in_ready; // @[LazyModule.scala 167:57]
  assign accumulator_auto_slave_in_valid = auto_accumulator_slave_in_valid; // @[LazyModule.scala 173:31]
  assign accumulator_auto_slave_in_bits_data = auto_accumulator_slave_in_bits_data; // @[LazyModule.scala 173:31]
  assign accumulator_auto_slave_in_bits_last = auto_accumulator_slave_in_bits_last; // @[LazyModule.scala 173:31]
  assign dspQueue_clock = clock;
  assign dspQueue_reset = reset;
  assign dspQueue_auto_stream_in_valid = accumulator_auto_master_out_valid; // @[LazyModule.scala 167:57]
  assign dspQueue_auto_stream_in_bits_data = accumulator_auto_master_out_bits_data; // @[LazyModule.scala 167:57]
  assign dspQueue_auto_stream_in_bits_last = accumulator_auto_master_out_bits_last; // @[LazyModule.scala 167:57]
  assign dspQueue_auto_stream_out_ready = auto_dspQueue_stream_out_ready; // @[LazyModule.scala 173:49]
  assign dspQueue_auto_in_aw_valid = axi4buf_auto_out_aw_valid; // @[LazyModule.scala 167:31]
  assign dspQueue_auto_in_aw_bits_id = axi4buf_auto_out_aw_bits_id; // @[LazyModule.scala 167:31]
  assign dspQueue_auto_in_aw_bits_addr = axi4buf_auto_out_aw_bits_addr; // @[LazyModule.scala 167:31]
  assign dspQueue_auto_in_w_valid = axi4buf_auto_out_w_valid; // @[LazyModule.scala 167:31]
  assign dspQueue_auto_in_w_bits_data = axi4buf_auto_out_w_bits_data; // @[LazyModule.scala 167:31]
  assign dspQueue_auto_in_w_bits_strb = axi4buf_auto_out_w_bits_strb; // @[LazyModule.scala 167:31]
  assign dspQueue_auto_in_b_ready = axi4buf_auto_out_b_ready; // @[LazyModule.scala 167:31]
  assign dspQueue_auto_in_ar_valid = axi4buf_auto_out_ar_valid; // @[LazyModule.scala 167:31]
  assign dspQueue_auto_in_ar_bits_id = axi4buf_auto_out_ar_bits_id; // @[LazyModule.scala 167:31]
  assign dspQueue_auto_in_ar_bits_addr = axi4buf_auto_out_ar_bits_addr; // @[LazyModule.scala 167:31]
  assign dspQueue_auto_in_ar_bits_size = axi4buf_auto_out_ar_bits_size; // @[LazyModule.scala 167:31]
  assign dspQueue_auto_in_r_ready = axi4buf_auto_out_r_ready; // @[LazyModule.scala 167:31]
  assign bus_clock = clock;
  assign bus_reset = reset;
  assign bus_auto_in_aw_valid = auto_bus_in_aw_valid; // @[LazyModule.scala 173:31]
  assign bus_auto_in_aw_bits_id = auto_bus_in_aw_bits_id; // @[LazyModule.scala 173:31]
  assign bus_auto_in_aw_bits_addr = auto_bus_in_aw_bits_addr; // @[LazyModule.scala 173:31]
  assign bus_auto_in_aw_bits_size = auto_bus_in_aw_bits_size; // @[LazyModule.scala 173:31]
  assign bus_auto_in_w_valid = auto_bus_in_w_valid; // @[LazyModule.scala 173:31]
  assign bus_auto_in_w_bits_data = auto_bus_in_w_bits_data; // @[LazyModule.scala 173:31]
  assign bus_auto_in_w_bits_strb = auto_bus_in_w_bits_strb; // @[LazyModule.scala 173:31]
  assign bus_auto_in_w_bits_last = auto_bus_in_w_bits_last; // @[LazyModule.scala 173:31]
  assign bus_auto_in_b_ready = auto_bus_in_b_ready; // @[LazyModule.scala 173:31]
  assign bus_auto_in_ar_valid = auto_bus_in_ar_valid; // @[LazyModule.scala 173:31]
  assign bus_auto_in_ar_bits_id = auto_bus_in_ar_bits_id; // @[LazyModule.scala 173:31]
  assign bus_auto_in_ar_bits_addr = auto_bus_in_ar_bits_addr; // @[LazyModule.scala 173:31]
  assign bus_auto_in_ar_bits_size = auto_bus_in_ar_bits_size; // @[LazyModule.scala 173:31]
  assign bus_auto_in_r_ready = auto_bus_in_r_ready; // @[LazyModule.scala 173:31]
  assign bus_auto_out_1_aw_ready = axi4buf_1_auto_in_aw_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_1_w_ready = axi4buf_1_auto_in_w_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_1_b_valid = axi4buf_1_auto_in_b_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_1_b_bits_id = axi4buf_1_auto_in_b_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_1_b_bits_resp = axi4buf_1_auto_in_b_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_1_ar_ready = axi4buf_1_auto_in_ar_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_1_r_valid = axi4buf_1_auto_in_r_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_1_r_bits_id = axi4buf_1_auto_in_r_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_1_r_bits_data = axi4buf_1_auto_in_r_bits_data; // @[LazyModule.scala 167:57]
  assign bus_auto_out_1_r_bits_resp = axi4buf_1_auto_in_r_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_1_r_bits_last = axi4buf_1_auto_in_r_bits_last; // @[LazyModule.scala 167:57]
  assign bus_auto_out_0_aw_ready = axi4buf_auto_in_aw_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_0_w_ready = axi4buf_auto_in_w_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_0_b_valid = axi4buf_auto_in_b_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_0_b_bits_id = axi4buf_auto_in_b_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_0_b_bits_resp = axi4buf_auto_in_b_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_0_ar_ready = axi4buf_auto_in_ar_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_0_r_valid = axi4buf_auto_in_r_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_0_r_bits_id = axi4buf_auto_in_r_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_0_r_bits_data = axi4buf_auto_in_r_bits_data; // @[LazyModule.scala 167:57]
  assign bus_auto_out_0_r_bits_resp = axi4buf_auto_in_r_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_0_r_bits_last = axi4buf_auto_in_r_bits_last; // @[LazyModule.scala 167:57]
  assign axi4buf_clock = clock;
  assign axi4buf_reset = reset;
  assign axi4buf_auto_in_aw_valid = bus_auto_out_0_aw_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_auto_in_aw_bits_id = bus_auto_out_0_aw_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_auto_in_aw_bits_addr = bus_auto_out_0_aw_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_auto_in_aw_bits_size = bus_auto_out_0_aw_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_auto_in_w_valid = bus_auto_out_0_w_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_auto_in_w_bits_data = bus_auto_out_0_w_bits_data; // @[LazyModule.scala 167:57]
  assign axi4buf_auto_in_w_bits_strb = bus_auto_out_0_w_bits_strb; // @[LazyModule.scala 167:57]
  assign axi4buf_auto_in_w_bits_last = bus_auto_out_0_w_bits_last; // @[LazyModule.scala 167:57]
  assign axi4buf_auto_in_b_ready = bus_auto_out_0_b_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_auto_in_ar_valid = bus_auto_out_0_ar_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_auto_in_ar_bits_id = bus_auto_out_0_ar_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_auto_in_ar_bits_addr = bus_auto_out_0_ar_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_auto_in_ar_bits_size = bus_auto_out_0_ar_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_auto_in_r_ready = bus_auto_out_0_r_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_auto_out_aw_ready = dspQueue_auto_in_aw_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_auto_out_w_ready = dspQueue_auto_in_w_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_auto_out_b_valid = dspQueue_auto_in_b_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_auto_out_b_bits_id = dspQueue_auto_in_b_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_auto_out_b_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_auto_out_ar_ready = dspQueue_auto_in_ar_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_auto_out_r_valid = dspQueue_auto_in_r_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_auto_out_r_bits_id = dspQueue_auto_in_r_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_auto_out_r_bits_data = dspQueue_auto_in_r_bits_data; // @[LazyModule.scala 167:31]
  assign axi4buf_auto_out_r_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_auto_out_r_bits_last = 1'h1; // @[LazyModule.scala 167:31]
  assign axi4buf_1_clock = clock;
  assign axi4buf_1_reset = reset;
  assign axi4buf_1_auto_in_aw_valid = bus_auto_out_1_aw_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_1_auto_in_aw_bits_id = bus_auto_out_1_aw_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_1_auto_in_aw_bits_addr = bus_auto_out_1_aw_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_1_auto_in_aw_bits_size = bus_auto_out_1_aw_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_1_auto_in_w_valid = bus_auto_out_1_w_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_1_auto_in_w_bits_data = bus_auto_out_1_w_bits_data; // @[LazyModule.scala 167:57]
  assign axi4buf_1_auto_in_w_bits_strb = bus_auto_out_1_w_bits_strb; // @[LazyModule.scala 167:57]
  assign axi4buf_1_auto_in_w_bits_last = bus_auto_out_1_w_bits_last; // @[LazyModule.scala 167:57]
  assign axi4buf_1_auto_in_b_ready = bus_auto_out_1_b_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_1_auto_in_ar_valid = bus_auto_out_1_ar_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_1_auto_in_ar_bits_id = bus_auto_out_1_ar_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_1_auto_in_ar_bits_addr = bus_auto_out_1_ar_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_1_auto_in_ar_bits_size = bus_auto_out_1_ar_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_1_auto_in_r_ready = bus_auto_out_1_r_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_1_auto_out_aw_ready = accumulator_auto_mem_in_aw_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_1_auto_out_w_ready = accumulator_auto_mem_in_w_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_1_auto_out_b_valid = accumulator_auto_mem_in_b_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_1_auto_out_b_bits_id = accumulator_auto_mem_in_b_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_1_auto_out_b_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_1_auto_out_ar_ready = accumulator_auto_mem_in_ar_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_1_auto_out_r_valid = accumulator_auto_mem_in_r_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_1_auto_out_r_bits_id = accumulator_auto_mem_in_r_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_1_auto_out_r_bits_data = accumulator_auto_mem_in_r_bits_data; // @[LazyModule.scala 167:31]
  assign axi4buf_1_auto_out_r_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_1_auto_out_r_bits_last = 1'h1; // @[LazyModule.scala 167:31]
endmodule
module AXI4StreamWidthAdapater_2_to_1(
  input         clock,
  input         reset,
  output        auto_in_ready,
  input         auto_in_valid,
  input  [15:0] auto_in_bits_data,
  input         auto_in_bits_last,
  input         auto_out_ready,
  output        auto_out_valid,
  output [31:0] auto_out_bits_data,
  output        auto_out_bits_last
);
  reg [15:0] _T; // @[AXI4StreamWidthAdapter.scala 101:37]
  reg [31:0] _RAND_0;
  reg  _T_1; // @[AXI4StreamWidthAdapter.scala 102:22]
  reg [31:0] _RAND_1;
  wire  _T_2; // @[AXI4StreamWidthAdapter.scala 103:14]
  wire [1:0] _T_4; // @[AXI4StreamWidthAdapter.scala 103:60]
  wire [1:0] _T_5; // @[AXI4StreamWidthAdapter.scala 103:33]
  wire [1:0] _GEN_0; // @[AXI4StreamWidthAdapter.scala 103:21]
  wire  _T_7; // @[AXI4StreamWidthAdapter.scala 106:29]
  wire  _T_8; // @[AXI4StreamWidthAdapter.scala 106:22]
  wire  ov0; // @[AXI4StreamWidthAdapter.scala 112:32]
  reg  _T_10; // @[AXI4StreamWidthAdapter.scala 101:37]
  reg [31:0] _RAND_2;
  reg  _T_11; // @[AXI4StreamWidthAdapter.scala 102:22]
  reg [31:0] _RAND_3;
  wire [1:0] _T_14; // @[AXI4StreamWidthAdapter.scala 103:60]
  wire [1:0] _T_15; // @[AXI4StreamWidthAdapter.scala 103:33]
  wire [1:0] _GEN_2; // @[AXI4StreamWidthAdapter.scala 103:21]
  wire  _T_17; // @[AXI4StreamWidthAdapter.scala 106:29]
  wire  _T_18; // @[AXI4StreamWidthAdapter.scala 106:22]
  wire [1:0] _T_19; // @[Cat.scala 29:58]
  wire  ov1; // @[AXI4StreamWidthAdapter.scala 112:32]
  reg  _T_22; // @[AXI4StreamWidthAdapter.scala 102:22]
  reg [31:0] _RAND_4;
  wire [1:0] _T_25; // @[AXI4StreamWidthAdapter.scala 103:60]
  wire [1:0] _T_26; // @[AXI4StreamWidthAdapter.scala 103:33]
  wire [1:0] _GEN_4; // @[AXI4StreamWidthAdapter.scala 103:21]
  wire  ov2; // @[AXI4StreamWidthAdapter.scala 112:32]
  reg  _T_32; // @[AXI4StreamWidthAdapter.scala 102:22]
  reg [31:0] _RAND_5;
  wire [1:0] _T_35; // @[AXI4StreamWidthAdapter.scala 103:60]
  wire [1:0] _T_36; // @[AXI4StreamWidthAdapter.scala 103:33]
  wire [1:0] _GEN_6; // @[AXI4StreamWidthAdapter.scala 103:21]
  wire  ov3; // @[AXI4StreamWidthAdapter.scala 112:32]
  reg  _T_42; // @[AXI4StreamWidthAdapter.scala 102:22]
  reg [31:0] _RAND_6;
  wire [1:0] _T_45; // @[AXI4StreamWidthAdapter.scala 103:60]
  wire [1:0] _T_46; // @[AXI4StreamWidthAdapter.scala 103:33]
  wire [1:0] _GEN_8; // @[AXI4StreamWidthAdapter.scala 103:21]
  wire  ov4; // @[AXI4StreamWidthAdapter.scala 112:32]
  wire  _T_51; // @[AXI4StreamWidthAdapter.scala 42:16]
  wire  _T_53; // @[AXI4StreamWidthAdapter.scala 42:11]
  wire  _T_54; // @[AXI4StreamWidthAdapter.scala 42:11]
  wire  _T_55; // @[AXI4StreamWidthAdapter.scala 43:16]
  wire  _T_57; // @[AXI4StreamWidthAdapter.scala 43:11]
  wire  _T_58; // @[AXI4StreamWidthAdapter.scala 43:11]
  wire  _T_59; // @[AXI4StreamWidthAdapter.scala 44:16]
  wire  _T_61; // @[AXI4StreamWidthAdapter.scala 44:11]
  wire  _T_62; // @[AXI4StreamWidthAdapter.scala 44:11]
  wire  _T_63; // @[AXI4StreamWidthAdapter.scala 45:16]
  wire  _T_65; // @[AXI4StreamWidthAdapter.scala 45:11]
  wire  _T_66; // @[AXI4StreamWidthAdapter.scala 45:11]
  assign _T_2 = auto_in_valid & auto_out_ready; // @[AXI4StreamWidthAdapter.scala 103:14]
  assign _T_4 = _T_1 + 1'h1; // @[AXI4StreamWidthAdapter.scala 103:60]
  assign _T_5 = _T_1 ? 2'h0 : _T_4; // @[AXI4StreamWidthAdapter.scala 103:33]
  assign _GEN_0 = _T_2 ? _T_5 : {{1'd0}, _T_1}; // @[AXI4StreamWidthAdapter.scala 103:21]
  assign _T_7 = ~_T_1; // @[AXI4StreamWidthAdapter.scala 106:29]
  assign _T_8 = _T_2 & _T_7; // @[AXI4StreamWidthAdapter.scala 106:22]
  assign ov0 = _T_1 & auto_in_valid; // @[AXI4StreamWidthAdapter.scala 112:32]
  assign _T_14 = _T_11 + 1'h1; // @[AXI4StreamWidthAdapter.scala 103:60]
  assign _T_15 = _T_11 ? 2'h0 : _T_14; // @[AXI4StreamWidthAdapter.scala 103:33]
  assign _GEN_2 = _T_2 ? _T_15 : {{1'd0}, _T_11}; // @[AXI4StreamWidthAdapter.scala 103:21]
  assign _T_17 = ~_T_11; // @[AXI4StreamWidthAdapter.scala 106:29]
  assign _T_18 = _T_2 & _T_17; // @[AXI4StreamWidthAdapter.scala 106:22]
  assign _T_19 = {auto_in_bits_last,_T_10}; // @[Cat.scala 29:58]
  assign ov1 = _T_11 & auto_in_valid; // @[AXI4StreamWidthAdapter.scala 112:32]
  assign _T_25 = _T_22 + 1'h1; // @[AXI4StreamWidthAdapter.scala 103:60]
  assign _T_26 = _T_22 ? 2'h0 : _T_25; // @[AXI4StreamWidthAdapter.scala 103:33]
  assign _GEN_4 = _T_2 ? _T_26 : {{1'd0}, _T_22}; // @[AXI4StreamWidthAdapter.scala 103:21]
  assign ov2 = _T_22 & auto_in_valid; // @[AXI4StreamWidthAdapter.scala 112:32]
  assign _T_35 = _T_32 + 1'h1; // @[AXI4StreamWidthAdapter.scala 103:60]
  assign _T_36 = _T_32 ? 2'h0 : _T_35; // @[AXI4StreamWidthAdapter.scala 103:33]
  assign _GEN_6 = _T_2 ? _T_36 : {{1'd0}, _T_32}; // @[AXI4StreamWidthAdapter.scala 103:21]
  assign ov3 = _T_32 & auto_in_valid; // @[AXI4StreamWidthAdapter.scala 112:32]
  assign _T_45 = _T_42 + 1'h1; // @[AXI4StreamWidthAdapter.scala 103:60]
  assign _T_46 = _T_42 ? 2'h0 : _T_45; // @[AXI4StreamWidthAdapter.scala 103:33]
  assign _GEN_8 = _T_2 ? _T_46 : {{1'd0}, _T_42}; // @[AXI4StreamWidthAdapter.scala 103:21]
  assign ov4 = _T_42 & auto_in_valid; // @[AXI4StreamWidthAdapter.scala 112:32]
  assign _T_51 = ov0 == ov1; // @[AXI4StreamWidthAdapter.scala 42:16]
  assign _T_53 = _T_51 | reset; // @[AXI4StreamWidthAdapter.scala 42:11]
  assign _T_54 = ~_T_53; // @[AXI4StreamWidthAdapter.scala 42:11]
  assign _T_55 = ov0 == ov2; // @[AXI4StreamWidthAdapter.scala 43:16]
  assign _T_57 = _T_55 | reset; // @[AXI4StreamWidthAdapter.scala 43:11]
  assign _T_58 = ~_T_57; // @[AXI4StreamWidthAdapter.scala 43:11]
  assign _T_59 = ov0 == ov3; // @[AXI4StreamWidthAdapter.scala 44:16]
  assign _T_61 = _T_59 | reset; // @[AXI4StreamWidthAdapter.scala 44:11]
  assign _T_62 = ~_T_61; // @[AXI4StreamWidthAdapter.scala 44:11]
  assign _T_63 = ov0 == ov4; // @[AXI4StreamWidthAdapter.scala 45:16]
  assign _T_65 = _T_63 | reset; // @[AXI4StreamWidthAdapter.scala 45:11]
  assign _T_66 = ~_T_65; // @[AXI4StreamWidthAdapter.scala 45:11]
  assign auto_in_ready = auto_out_ready; // @[LazyModule.scala 173:31]
  assign auto_out_valid = _T_1 & auto_in_valid; // @[LazyModule.scala 173:49]
  assign auto_out_bits_data = {auto_in_bits_data,_T}; // @[LazyModule.scala 173:49]
  assign auto_out_bits_last = _T_19 != 2'h0; // @[LazyModule.scala 173:49]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_10 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_11 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_22 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_32 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_42 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (_T_8) begin
      _T <= auto_in_bits_data;
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else begin
      _T_1 <= _GEN_0[0];
    end
    if (_T_18) begin
      _T_10 <= auto_in_bits_last;
    end
    if (reset) begin
      _T_11 <= 1'h0;
    end else begin
      _T_11 <= _GEN_2[0];
    end
    if (reset) begin
      _T_22 <= 1'h0;
    end else begin
      _T_22 <= _GEN_4[0];
    end
    if (reset) begin
      _T_32 <= 1'h0;
    end else begin
      _T_32 <= _GEN_6[0];
    end
    if (reset) begin
      _T_42 <= 1'h0;
    end else begin
      _T_42 <= _GEN_8[0];
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_54) begin
          $fwrite(32'h80000002,"Assertion failed\n    at AXI4StreamWidthAdapter.scala:42 assert(ov0 === ov1)\n"); // @[AXI4StreamWidthAdapter.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_54) begin
          $fatal; // @[AXI4StreamWidthAdapter.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_58) begin
          $fwrite(32'h80000002,"Assertion failed\n    at AXI4StreamWidthAdapter.scala:43 assert(ov0 === ov2)\n"); // @[AXI4StreamWidthAdapter.scala 43:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_58) begin
          $fatal; // @[AXI4StreamWidthAdapter.scala 43:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_62) begin
          $fwrite(32'h80000002,"Assertion failed\n    at AXI4StreamWidthAdapter.scala:44 assert(ov0 === ov3)\n"); // @[AXI4StreamWidthAdapter.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_62) begin
          $fatal; // @[AXI4StreamWidthAdapter.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_66) begin
          $fwrite(32'h80000002,"Assertion failed\n    at AXI4StreamWidthAdapter.scala:45 assert(ov0 === ov4)\n"); // @[AXI4StreamWidthAdapter.scala 45:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_66) begin
          $fatal; // @[AXI4StreamWidthAdapter.scala 45:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module Queue_35(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [31:0] io_enq_bits_data,
  input         io_enq_bits_last,
  input         io_deq_ready,
  output        io_deq_valid,
  output [31:0] io_deq_bits_data,
  output        io_deq_bits_last
);
  reg [31:0] _T_data [0:0]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_0;
  wire [31:0] _T_data__T_14_data; // @[Decoupled.scala 209:24]
  wire  _T_data__T_14_addr; // @[Decoupled.scala 209:24]
  wire [31:0] _T_data__T_10_data; // @[Decoupled.scala 209:24]
  wire  _T_data__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T_data__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T_data__T_10_en; // @[Decoupled.scala 209:24]
  reg  _T_last [0:0]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_1;
  wire  _T_last__T_14_data; // @[Decoupled.scala 209:24]
  wire  _T_last__T_14_addr; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_data; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_en; // @[Decoupled.scala 209:24]
  reg  _T_1; // @[Decoupled.scala 212:35]
  reg [31:0] _RAND_2;
  wire  _T_3; // @[Decoupled.scala 215:36]
  wire  _T_6; // @[Decoupled.scala 40:37]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[Decoupled.scala 240:27]
  wire  _GEN_22; // @[Decoupled.scala 237:18]
  wire  _GEN_21; // @[Decoupled.scala 237:18]
  wire  _T_11; // @[Decoupled.scala 227:16]
  wire  _T_12; // @[Decoupled.scala 231:19]
  assign _T_data__T_14_addr = 1'h0;
  assign _T_data__T_14_data = _T_data[_T_data__T_14_addr]; // @[Decoupled.scala 209:24]
  assign _T_data__T_10_data = io_enq_bits_data;
  assign _T_data__T_10_addr = 1'h0;
  assign _T_data__T_10_mask = 1'h1;
  assign _T_data__T_10_en = _T_3 ? _GEN_13 : _T_6;
  assign _T_last__T_14_addr = 1'h0;
  assign _T_last__T_14_data = _T_last[_T_last__T_14_addr]; // @[Decoupled.scala 209:24]
  assign _T_last__T_10_data = io_enq_bits_last;
  assign _T_last__T_10_addr = 1'h0;
  assign _T_last__T_10_mask = 1'h1;
  assign _T_last__T_10_en = _T_3 ? _GEN_13 : _T_6;
  assign _T_3 = ~_T_1; // @[Decoupled.scala 215:36]
  assign _T_6 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  assign _T_8 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = io_deq_ready ? 1'h0 : _T_6; // @[Decoupled.scala 240:27]
  assign _GEN_22 = _T_3 ? _GEN_13 : _T_6; // @[Decoupled.scala 237:18]
  assign _GEN_21 = _T_3 ? 1'h0 : _T_8; // @[Decoupled.scala 237:18]
  assign _T_11 = _GEN_22 != _GEN_21; // @[Decoupled.scala 227:16]
  assign _T_12 = ~_T_3; // @[Decoupled.scala 231:19]
  assign io_enq_ready = io_deq_ready | _T_3; // @[Decoupled.scala 232:16 Decoupled.scala 245:40]
  assign io_deq_valid = io_enq_valid | _T_12; // @[Decoupled.scala 231:16 Decoupled.scala 236:40]
  assign io_deq_bits_data = _T_3 ? io_enq_bits_data : _T_data__T_14_data; // @[Decoupled.scala 233:15 Decoupled.scala 238:19]
  assign io_deq_bits_last = _T_3 ? io_enq_bits_last : _T_last__T_14_data; // @[Decoupled.scala 233:15 Decoupled.scala 238:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_data[initvar] = _RAND_0[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_last[initvar] = _RAND_1[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_1 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T_data__T_10_en & _T_data__T_10_mask) begin
      _T_data[_T_data__T_10_addr] <= _T_data__T_10_data; // @[Decoupled.scala 209:24]
    end
    if(_T_last__T_10_en & _T_last__T_10_mask) begin
      _T_last[_T_last__T_10_addr] <= _T_last__T_10_data; // @[Decoupled.scala 209:24]
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else if (_T_11) begin
      if (_T_3) begin
        if (io_deq_ready) begin
          _T_1 <= 1'h0;
        end else begin
          _T_1 <= _T_6;
        end
      end else begin
        _T_1 <= _T_6;
      end
    end
  end
endmodule
module StreamBuffer_1(
  input         clock,
  input         reset,
  input         auto_out_out_ready,
  output        auto_out_out_valid,
  output [31:0] auto_out_out_bits_data,
  output        auto_out_out_bits_last,
  output        auto_in_in_ready,
  input         auto_in_in_valid,
  input  [31:0] auto_in_in_bits_data,
  input         auto_in_in_bits_last
);
  wire  Queue_clock; // @[Decoupled.scala 287:21]
  wire  Queue_reset; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_enq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_last; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_deq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_last; // @[Decoupled.scala 287:21]
  Queue_35 Queue ( // @[Decoupled.scala 287:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_last(Queue_io_enq_bits_last),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_last(Queue_io_deq_bits_last)
  );
  assign auto_out_out_valid = Queue_io_deq_valid; // @[LazyModule.scala 173:49]
  assign auto_out_out_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_out_bits_last = Queue_io_deq_bits_last; // @[LazyModule.scala 173:49]
  assign auto_in_in_ready = Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_in_in_valid; // @[Decoupled.scala 288:22]
  assign Queue_io_enq_bits_data = auto_in_in_bits_data; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_last = auto_in_in_bits_last; // @[Decoupled.scala 289:21]
  assign Queue_io_deq_ready = auto_out_out_ready; // @[Decoupled.scala 311:15]
endmodule
module AXI4StreamMux_8(
  input         clock,
  input         reset,
  output        auto_register_in_aw_ready,
  input         auto_register_in_aw_valid,
  input         auto_register_in_aw_bits_id,
  input  [29:0] auto_register_in_aw_bits_addr,
  output        auto_register_in_w_ready,
  input         auto_register_in_w_valid,
  input  [31:0] auto_register_in_w_bits_data,
  input  [3:0]  auto_register_in_w_bits_strb,
  input         auto_register_in_b_ready,
  output        auto_register_in_b_valid,
  output        auto_register_in_b_bits_id,
  output        auto_register_in_ar_ready,
  input         auto_register_in_ar_valid,
  input         auto_register_in_ar_bits_id,
  input  [29:0] auto_register_in_ar_bits_addr,
  input  [2:0]  auto_register_in_ar_bits_size,
  input         auto_register_in_r_ready,
  output        auto_register_in_r_valid,
  output        auto_register_in_r_bits_id,
  output [31:0] auto_register_in_r_bits_data,
  output        auto_stream_in_6_ready,
  input         auto_stream_in_6_valid,
  input  [31:0] auto_stream_in_6_bits_data,
  input         auto_stream_in_6_bits_last,
  output        auto_stream_in_5_ready,
  input         auto_stream_in_5_valid,
  input  [31:0] auto_stream_in_5_bits_data,
  input         auto_stream_in_5_bits_last,
  output        auto_stream_in_4_ready,
  input         auto_stream_in_4_valid,
  input  [31:0] auto_stream_in_4_bits_data,
  input         auto_stream_in_4_bits_last,
  output        auto_stream_in_3_ready,
  input         auto_stream_in_3_valid,
  input  [31:0] auto_stream_in_3_bits_data,
  input         auto_stream_in_3_bits_last,
  output        auto_stream_in_2_ready,
  input         auto_stream_in_2_valid,
  input  [31:0] auto_stream_in_2_bits_data,
  input         auto_stream_in_2_bits_last,
  output        auto_stream_in_1_ready,
  input         auto_stream_in_1_valid,
  input  [31:0] auto_stream_in_1_bits_data,
  input         auto_stream_in_1_bits_last,
  output        auto_stream_in_0_ready,
  input         auto_stream_in_0_valid,
  input  [31:0] auto_stream_in_0_bits_data,
  input         auto_stream_in_0_bits_last,
  input         auto_stream_out_1_ready,
  output        auto_stream_out_1_valid,
  output [31:0] auto_stream_out_1_bits_data,
  output        auto_stream_out_1_bits_last,
  input         auto_stream_out_0_ready,
  output        auto_stream_out_0_valid,
  output [31:0] auto_stream_out_0_bits_data,
  output        auto_stream_out_0_bits_last
);
  wire  Queue_clock; // @[Decoupled.scala 287:21]
  wire  Queue_reset; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_read; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_enq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_extra; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_read; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_deq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_extra; // @[Decoupled.scala 287:21]
  reg [2:0] sels_0; // @[Mux.scala 32:23]
  reg [31:0] _RAND_0;
  reg [2:0] sels_1; // @[Mux.scala 32:23]
  reg [31:0] _RAND_1;
  reg [2:0] sels_2; // @[Mux.scala 32:23]
  reg [31:0] _RAND_2;
  wire  _T_3; // @[Mux.scala 45:28]
  wire  _GEN_7; // @[Mux.scala 45:41]
  wire  _GEN_8; // @[Mux.scala 45:41]
  wire  _T_4; // @[Mux.scala 45:28]
  wire  _GEN_12; // @[Mux.scala 45:41]
  wire [31:0] _GEN_15; // @[Mux.scala 45:41]
  wire  _GEN_16; // @[Mux.scala 45:41]
  wire  _GEN_17; // @[Mux.scala 45:41]
  wire  _T_5; // @[Mux.scala 45:28]
  wire  _GEN_21; // @[Mux.scala 45:41]
  wire [31:0] _GEN_24; // @[Mux.scala 45:41]
  wire  _GEN_25; // @[Mux.scala 45:41]
  wire  _GEN_26; // @[Mux.scala 45:41]
  wire  _T_6; // @[Mux.scala 45:28]
  wire  _GEN_30; // @[Mux.scala 45:41]
  wire [31:0] _GEN_33; // @[Mux.scala 45:41]
  wire  _GEN_34; // @[Mux.scala 45:41]
  wire  _GEN_35; // @[Mux.scala 45:41]
  wire  _T_7; // @[Mux.scala 45:28]
  wire  _GEN_39; // @[Mux.scala 45:41]
  wire [31:0] _GEN_42; // @[Mux.scala 45:41]
  wire  _GEN_43; // @[Mux.scala 45:41]
  wire  _GEN_44; // @[Mux.scala 45:41]
  wire  _T_8; // @[Mux.scala 45:28]
  wire  _GEN_48; // @[Mux.scala 45:41]
  wire [31:0] _GEN_51; // @[Mux.scala 45:41]
  wire  _GEN_52; // @[Mux.scala 45:41]
  wire  _GEN_53; // @[Mux.scala 45:41]
  wire  _T_9; // @[Mux.scala 45:28]
  wire  _GEN_62; // @[Mux.scala 45:41]
  wire  _T_10; // @[Mux.scala 40:46]
  wire [2:0] _T_12; // @[Mux.scala 41:29]
  wire  _T_13; // @[Mux.scala 45:28]
  wire  _GEN_70; // @[Mux.scala 45:41]
  wire  _GEN_71; // @[Mux.scala 45:41]
  wire  _T_14; // @[Mux.scala 45:28]
  wire  _GEN_75; // @[Mux.scala 45:41]
  wire [31:0] _GEN_78; // @[Mux.scala 45:41]
  wire  _GEN_79; // @[Mux.scala 45:41]
  wire  _GEN_80; // @[Mux.scala 45:41]
  wire  _T_15; // @[Mux.scala 45:28]
  wire  _GEN_84; // @[Mux.scala 45:41]
  wire [31:0] _GEN_87; // @[Mux.scala 45:41]
  wire  _GEN_88; // @[Mux.scala 45:41]
  wire  _GEN_89; // @[Mux.scala 45:41]
  wire  _T_16; // @[Mux.scala 45:28]
  wire  _GEN_93; // @[Mux.scala 45:41]
  wire [31:0] _GEN_96; // @[Mux.scala 45:41]
  wire  _GEN_97; // @[Mux.scala 45:41]
  wire  _GEN_98; // @[Mux.scala 45:41]
  wire  _T_17; // @[Mux.scala 45:28]
  wire  _GEN_102; // @[Mux.scala 45:41]
  wire [31:0] _GEN_105; // @[Mux.scala 45:41]
  wire  _GEN_106; // @[Mux.scala 45:41]
  wire  _GEN_107; // @[Mux.scala 45:41]
  wire  _T_18; // @[Mux.scala 45:28]
  wire  _GEN_111; // @[Mux.scala 45:41]
  wire [31:0] _GEN_114; // @[Mux.scala 45:41]
  wire  _GEN_115; // @[Mux.scala 45:41]
  wire  _GEN_116; // @[Mux.scala 45:41]
  wire  _T_19; // @[Mux.scala 45:28]
  wire  _GEN_125; // @[Mux.scala 45:41]
  wire  _T_20; // @[Mux.scala 40:46]
  wire  _T_21; // @[Mux.scala 40:46]
  wire  _T_23; // @[Mux.scala 40:75]
  wire [2:0] _T_24; // @[Mux.scala 41:29]
  wire  _T_25; // @[Mux.scala 45:28]
  wire  _T_26; // @[Mux.scala 45:28]
  wire  _T_27; // @[Mux.scala 45:28]
  wire  _T_28; // @[Mux.scala 45:28]
  wire  _T_29; // @[Mux.scala 45:28]
  wire  _T_30; // @[Mux.scala 45:28]
  wire  _T_31; // @[Mux.scala 45:28]
  wire  _T_33; // @[RegisterRouter.scala 40:39]
  wire  _T_34; // @[RegisterRouter.scala 40:26]
  wire  _T_35; // @[RegisterRouter.scala 42:29]
  wire  _T_78_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 290:17]
  wire [29:0] _T_42; // @[RegisterRouter.scala 48:19]
  wire [1:0] _T_197; // @[Cat.scala 29:58]
  wire  _T_36; // @[RegisterRouter.scala 42:26]
  wire [1:0] _T_45; // @[OneHot.scala 65:12]
  wire [1:0] _T_47; // @[Misc.scala 200:81]
  wire  _T_48; // @[Misc.scala 204:21]
  wire  _T_51; // @[Misc.scala 209:20]
  wire  _T_53; // @[Misc.scala 213:38]
  wire  _T_54; // @[Misc.scala 213:29]
  wire  _T_56; // @[Misc.scala 213:38]
  wire  _T_57; // @[Misc.scala 213:29]
  wire  _T_60; // @[Misc.scala 209:20]
  wire  _T_61; // @[Misc.scala 212:27]
  wire  _T_62; // @[Misc.scala 213:38]
  wire  _T_63; // @[Misc.scala 213:29]
  wire  _T_64; // @[Misc.scala 212:27]
  wire  _T_65; // @[Misc.scala 213:38]
  wire  _T_66; // @[Misc.scala 213:29]
  wire  _T_67; // @[Misc.scala 212:27]
  wire  _T_68; // @[Misc.scala 213:38]
  wire  _T_69; // @[Misc.scala 213:29]
  wire  _T_70; // @[Misc.scala 212:27]
  wire  _T_71; // @[Misc.scala 213:38]
  wire  _T_72; // @[Misc.scala 213:29]
  wire [3:0] _T_75; // @[Cat.scala 29:58]
  wire [3:0] _T_77; // @[RegisterRouter.scala 54:25]
  wire [7:0] _T_98; // @[Bitwise.scala 72:12]
  wire [7:0] _T_100; // @[Bitwise.scala 72:12]
  wire [7:0] _T_102; // @[Bitwise.scala 72:12]
  wire [7:0] _T_104; // @[Bitwise.scala 72:12]
  wire [31:0] _T_107; // @[Cat.scala 29:58]
  wire  _T_126; // @[RegisterRouter.scala 59:16]
  wire  _T_208; // @[RegisterRouter.scala 59:16]
  wire [3:0] _T_198; // @[OneHot.scala 58:35]
  wire  _T_235; // @[RegisterRouter.scala 59:16]
  wire  _T_247; // @[RegisterRouter.scala 59:16]
  wire  _T_133; // @[RegisterRouter.scala 59:16]
  wire  _T_242; // @[RegisterRouter.scala 59:16]
  wire  _T_156; // @[RegisterRouter.scala 59:16]
  wire  _T_237; // @[RegisterRouter.scala 59:16]
  wire  _T_179; // @[RegisterRouter.scala 59:16]
  wire [2:0] _GEN_213; // @[MuxLiteral.scala 48:10]
  wire [2:0] _GEN_214; // @[MuxLiteral.scala 48:10]
  wire [2:0] _GEN_215; // @[MuxLiteral.scala 48:10]
  wire  _T_323_bits_read; // @[Decoupled.scala 308:19 Decoupled.scala 309:14]
  wire  _T_323_valid; // @[Decoupled.scala 308:19 Decoupled.scala 310:15]
  wire  _T_326; // @[RegisterRouter.scala 65:29]
  Queue Queue ( // @[Decoupled.scala 287:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_read(Queue_io_enq_bits_read),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_extra(Queue_io_enq_bits_extra),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_read(Queue_io_deq_bits_read),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_extra(Queue_io_deq_bits_extra)
  );
  assign _T_3 = sels_0 == 3'h0; // @[Mux.scala 45:28]
  assign _GEN_7 = _T_3 & auto_stream_in_0_valid; // @[Mux.scala 45:41]
  assign _GEN_8 = _T_3 & auto_stream_out_0_ready; // @[Mux.scala 45:41]
  assign _T_4 = sels_0 == 3'h1; // @[Mux.scala 45:28]
  assign _GEN_12 = _T_4 ? auto_stream_in_1_bits_last : auto_stream_in_0_bits_last; // @[Mux.scala 45:41]
  assign _GEN_15 = _T_4 ? auto_stream_in_1_bits_data : auto_stream_in_0_bits_data; // @[Mux.scala 45:41]
  assign _GEN_16 = _T_4 ? auto_stream_in_1_valid : _GEN_7; // @[Mux.scala 45:41]
  assign _GEN_17 = _T_4 & auto_stream_out_0_ready; // @[Mux.scala 45:41]
  assign _T_5 = sels_0 == 3'h2; // @[Mux.scala 45:28]
  assign _GEN_21 = _T_5 ? auto_stream_in_2_bits_last : _GEN_12; // @[Mux.scala 45:41]
  assign _GEN_24 = _T_5 ? auto_stream_in_2_bits_data : _GEN_15; // @[Mux.scala 45:41]
  assign _GEN_25 = _T_5 ? auto_stream_in_2_valid : _GEN_16; // @[Mux.scala 45:41]
  assign _GEN_26 = _T_5 & auto_stream_out_0_ready; // @[Mux.scala 45:41]
  assign _T_6 = sels_0 == 3'h3; // @[Mux.scala 45:28]
  assign _GEN_30 = _T_6 ? auto_stream_in_3_bits_last : _GEN_21; // @[Mux.scala 45:41]
  assign _GEN_33 = _T_6 ? auto_stream_in_3_bits_data : _GEN_24; // @[Mux.scala 45:41]
  assign _GEN_34 = _T_6 ? auto_stream_in_3_valid : _GEN_25; // @[Mux.scala 45:41]
  assign _GEN_35 = _T_6 & auto_stream_out_0_ready; // @[Mux.scala 45:41]
  assign _T_7 = sels_0 == 3'h4; // @[Mux.scala 45:28]
  assign _GEN_39 = _T_7 ? auto_stream_in_4_bits_last : _GEN_30; // @[Mux.scala 45:41]
  assign _GEN_42 = _T_7 ? auto_stream_in_4_bits_data : _GEN_33; // @[Mux.scala 45:41]
  assign _GEN_43 = _T_7 ? auto_stream_in_4_valid : _GEN_34; // @[Mux.scala 45:41]
  assign _GEN_44 = _T_7 & auto_stream_out_0_ready; // @[Mux.scala 45:41]
  assign _T_8 = sels_0 == 3'h5; // @[Mux.scala 45:28]
  assign _GEN_48 = _T_8 ? auto_stream_in_5_bits_last : _GEN_39; // @[Mux.scala 45:41]
  assign _GEN_51 = _T_8 ? auto_stream_in_5_bits_data : _GEN_42; // @[Mux.scala 45:41]
  assign _GEN_52 = _T_8 ? auto_stream_in_5_valid : _GEN_43; // @[Mux.scala 45:41]
  assign _GEN_53 = _T_8 & auto_stream_out_0_ready; // @[Mux.scala 45:41]
  assign _T_9 = sels_0 == 3'h6; // @[Mux.scala 45:28]
  assign _GEN_62 = _T_9 & auto_stream_out_0_ready; // @[Mux.scala 45:41]
  assign _T_10 = sels_0 == sels_1; // @[Mux.scala 40:46]
  assign _T_12 = _T_10 ? 3'h7 : sels_1; // @[Mux.scala 41:29]
  assign _T_13 = _T_12 == 3'h0; // @[Mux.scala 45:28]
  assign _GEN_70 = _T_13 & auto_stream_in_0_valid; // @[Mux.scala 45:41]
  assign _GEN_71 = _T_13 ? auto_stream_out_1_ready : _GEN_8; // @[Mux.scala 45:41]
  assign _T_14 = _T_12 == 3'h1; // @[Mux.scala 45:28]
  assign _GEN_75 = _T_14 ? auto_stream_in_1_bits_last : auto_stream_in_0_bits_last; // @[Mux.scala 45:41]
  assign _GEN_78 = _T_14 ? auto_stream_in_1_bits_data : auto_stream_in_0_bits_data; // @[Mux.scala 45:41]
  assign _GEN_79 = _T_14 ? auto_stream_in_1_valid : _GEN_70; // @[Mux.scala 45:41]
  assign _GEN_80 = _T_14 ? auto_stream_out_1_ready : _GEN_17; // @[Mux.scala 45:41]
  assign _T_15 = _T_12 == 3'h2; // @[Mux.scala 45:28]
  assign _GEN_84 = _T_15 ? auto_stream_in_2_bits_last : _GEN_75; // @[Mux.scala 45:41]
  assign _GEN_87 = _T_15 ? auto_stream_in_2_bits_data : _GEN_78; // @[Mux.scala 45:41]
  assign _GEN_88 = _T_15 ? auto_stream_in_2_valid : _GEN_79; // @[Mux.scala 45:41]
  assign _GEN_89 = _T_15 ? auto_stream_out_1_ready : _GEN_26; // @[Mux.scala 45:41]
  assign _T_16 = _T_12 == 3'h3; // @[Mux.scala 45:28]
  assign _GEN_93 = _T_16 ? auto_stream_in_3_bits_last : _GEN_84; // @[Mux.scala 45:41]
  assign _GEN_96 = _T_16 ? auto_stream_in_3_bits_data : _GEN_87; // @[Mux.scala 45:41]
  assign _GEN_97 = _T_16 ? auto_stream_in_3_valid : _GEN_88; // @[Mux.scala 45:41]
  assign _GEN_98 = _T_16 ? auto_stream_out_1_ready : _GEN_35; // @[Mux.scala 45:41]
  assign _T_17 = _T_12 == 3'h4; // @[Mux.scala 45:28]
  assign _GEN_102 = _T_17 ? auto_stream_in_4_bits_last : _GEN_93; // @[Mux.scala 45:41]
  assign _GEN_105 = _T_17 ? auto_stream_in_4_bits_data : _GEN_96; // @[Mux.scala 45:41]
  assign _GEN_106 = _T_17 ? auto_stream_in_4_valid : _GEN_97; // @[Mux.scala 45:41]
  assign _GEN_107 = _T_17 ? auto_stream_out_1_ready : _GEN_44; // @[Mux.scala 45:41]
  assign _T_18 = _T_12 == 3'h5; // @[Mux.scala 45:28]
  assign _GEN_111 = _T_18 ? auto_stream_in_5_bits_last : _GEN_102; // @[Mux.scala 45:41]
  assign _GEN_114 = _T_18 ? auto_stream_in_5_bits_data : _GEN_105; // @[Mux.scala 45:41]
  assign _GEN_115 = _T_18 ? auto_stream_in_5_valid : _GEN_106; // @[Mux.scala 45:41]
  assign _GEN_116 = _T_18 ? auto_stream_out_1_ready : _GEN_53; // @[Mux.scala 45:41]
  assign _T_19 = _T_12 == 3'h6; // @[Mux.scala 45:28]
  assign _GEN_125 = _T_19 ? auto_stream_out_1_ready : _GEN_62; // @[Mux.scala 45:41]
  assign _T_20 = sels_0 == sels_2; // @[Mux.scala 40:46]
  assign _T_21 = sels_1 == sels_2; // @[Mux.scala 40:46]
  assign _T_23 = _T_20 | _T_21; // @[Mux.scala 40:75]
  assign _T_24 = _T_23 ? 3'h7 : sels_2; // @[Mux.scala 41:29]
  assign _T_25 = _T_24 == 3'h0; // @[Mux.scala 45:28]
  assign _T_26 = _T_24 == 3'h1; // @[Mux.scala 45:28]
  assign _T_27 = _T_24 == 3'h2; // @[Mux.scala 45:28]
  assign _T_28 = _T_24 == 3'h3; // @[Mux.scala 45:28]
  assign _T_29 = _T_24 == 3'h4; // @[Mux.scala 45:28]
  assign _T_30 = _T_24 == 3'h5; // @[Mux.scala 45:28]
  assign _T_31 = _T_24 == 3'h6; // @[Mux.scala 45:28]
  assign _T_33 = auto_register_in_aw_valid & auto_register_in_w_valid; // @[RegisterRouter.scala 40:39]
  assign _T_34 = auto_register_in_ar_valid | _T_33; // @[RegisterRouter.scala 40:26]
  assign _T_35 = ~auto_register_in_ar_valid; // @[RegisterRouter.scala 42:29]
  assign _T_78_ready = Queue_io_enq_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 290:17]
  assign _T_42 = auto_register_in_ar_valid ? auto_register_in_ar_bits_addr : auto_register_in_aw_bits_addr; // @[RegisterRouter.scala 48:19]
  assign _T_197 = {_T_42[3],_T_42[2]}; // @[Cat.scala 29:58]
  assign _T_36 = _T_78_ready & _T_35; // @[RegisterRouter.scala 42:26]
  assign _T_45 = 2'h1 << auto_register_in_ar_bits_size[0]; // @[OneHot.scala 65:12]
  assign _T_47 = _T_45 | 2'h1; // @[Misc.scala 200:81]
  assign _T_48 = auto_register_in_ar_bits_size >= 3'h2; // @[Misc.scala 204:21]
  assign _T_51 = ~auto_register_in_ar_bits_addr[1]; // @[Misc.scala 209:20]
  assign _T_53 = _T_47[1] & _T_51; // @[Misc.scala 213:38]
  assign _T_54 = _T_48 | _T_53; // @[Misc.scala 213:29]
  assign _T_56 = _T_47[1] & auto_register_in_ar_bits_addr[1]; // @[Misc.scala 213:38]
  assign _T_57 = _T_48 | _T_56; // @[Misc.scala 213:29]
  assign _T_60 = ~auto_register_in_ar_bits_addr[0]; // @[Misc.scala 209:20]
  assign _T_61 = _T_51 & _T_60; // @[Misc.scala 212:27]
  assign _T_62 = _T_47[0] & _T_61; // @[Misc.scala 213:38]
  assign _T_63 = _T_54 | _T_62; // @[Misc.scala 213:29]
  assign _T_64 = _T_51 & auto_register_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  assign _T_65 = _T_47[0] & _T_64; // @[Misc.scala 213:38]
  assign _T_66 = _T_54 | _T_65; // @[Misc.scala 213:29]
  assign _T_67 = auto_register_in_ar_bits_addr[1] & _T_60; // @[Misc.scala 212:27]
  assign _T_68 = _T_47[0] & _T_67; // @[Misc.scala 213:38]
  assign _T_69 = _T_57 | _T_68; // @[Misc.scala 213:29]
  assign _T_70 = auto_register_in_ar_bits_addr[1] & auto_register_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  assign _T_71 = _T_47[0] & _T_70; // @[Misc.scala 213:38]
  assign _T_72 = _T_57 | _T_71; // @[Misc.scala 213:29]
  assign _T_75 = {_T_72,_T_69,_T_66,_T_63}; // @[Cat.scala 29:58]
  assign _T_77 = auto_register_in_ar_valid ? _T_75 : auto_register_in_w_bits_strb; // @[RegisterRouter.scala 54:25]
  assign _T_98 = _T_77[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_100 = _T_77[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_102 = _T_77[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_104 = _T_77[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_107 = {_T_104,_T_102,_T_100,_T_98}; // @[Cat.scala 29:58]
  assign _T_126 = _T_107[2:0] == 3'h7; // @[RegisterRouter.scala 59:16]
  assign _T_208 = _T_34 & _T_78_ready; // @[RegisterRouter.scala 59:16]
  assign _T_198 = 4'h1 << _T_197; // @[OneHot.scala 58:35]
  assign _T_235 = _T_208 & _T_35; // @[RegisterRouter.scala 59:16]
  assign _T_247 = _T_235 & _T_198[2]; // @[RegisterRouter.scala 59:16]
  assign _T_133 = _T_247 & _T_126; // @[RegisterRouter.scala 59:16]
  assign _T_242 = _T_235 & _T_198[1]; // @[RegisterRouter.scala 59:16]
  assign _T_156 = _T_242 & _T_126; // @[RegisterRouter.scala 59:16]
  assign _T_237 = _T_235 & _T_198[0]; // @[RegisterRouter.scala 59:16]
  assign _T_179 = _T_237 & _T_126; // @[RegisterRouter.scala 59:16]
  assign _GEN_213 = 2'h1 == _T_197 ? sels_1 : sels_0; // @[MuxLiteral.scala 48:10]
  assign _GEN_214 = 2'h2 == _T_197 ? sels_2 : _GEN_213; // @[MuxLiteral.scala 48:10]
  assign _GEN_215 = 2'h3 == _T_197 ? 3'h0 : _GEN_214; // @[MuxLiteral.scala 48:10]
  assign _T_323_bits_read = Queue_io_deq_bits_read; // @[Decoupled.scala 308:19 Decoupled.scala 309:14]
  assign _T_323_valid = Queue_io_deq_valid; // @[Decoupled.scala 308:19 Decoupled.scala 310:15]
  assign _T_326 = ~_T_323_bits_read; // @[RegisterRouter.scala 65:29]
  assign auto_register_in_aw_ready = _T_36 & auto_register_in_w_valid; // @[LazyModule.scala 173:31]
  assign auto_register_in_w_ready = _T_36 & auto_register_in_aw_valid; // @[LazyModule.scala 173:31]
  assign auto_register_in_b_valid = _T_323_valid & _T_326; // @[LazyModule.scala 173:31]
  assign auto_register_in_b_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_register_in_ar_ready = Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_register_in_r_valid = _T_323_valid & _T_323_bits_read; // @[LazyModule.scala 173:31]
  assign auto_register_in_r_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_register_in_r_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 173:31]
  assign auto_stream_in_6_ready = _T_31 | _GEN_125; // @[LazyModule.scala 173:31]
  assign auto_stream_in_5_ready = _T_30 | _GEN_116; // @[LazyModule.scala 173:31]
  assign auto_stream_in_4_ready = _T_29 | _GEN_107; // @[LazyModule.scala 173:31]
  assign auto_stream_in_3_ready = _T_28 | _GEN_98; // @[LazyModule.scala 173:31]
  assign auto_stream_in_2_ready = _T_27 | _GEN_89; // @[LazyModule.scala 173:31]
  assign auto_stream_in_1_ready = _T_26 | _GEN_80; // @[LazyModule.scala 173:31]
  assign auto_stream_in_0_ready = _T_25 | _GEN_71; // @[LazyModule.scala 173:31]
  assign auto_stream_out_1_valid = _T_19 ? auto_stream_in_6_valid : _GEN_115; // @[LazyModule.scala 173:49]
  assign auto_stream_out_1_bits_data = _T_19 ? auto_stream_in_6_bits_data : _GEN_114; // @[LazyModule.scala 173:49]
  assign auto_stream_out_1_bits_last = _T_19 ? auto_stream_in_6_bits_last : _GEN_111; // @[LazyModule.scala 173:49]
  assign auto_stream_out_0_valid = _T_9 ? auto_stream_in_6_valid : _GEN_52; // @[LazyModule.scala 173:49]
  assign auto_stream_out_0_bits_data = _T_9 ? auto_stream_in_6_bits_data : _GEN_51; // @[LazyModule.scala 173:49]
  assign auto_stream_out_0_bits_last = _T_9 ? auto_stream_in_6_bits_last : _GEN_48; // @[LazyModule.scala 173:49]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_register_in_ar_valid | _T_33; // @[Decoupled.scala 288:22]
  assign Queue_io_enq_bits_read = auto_register_in_ar_valid; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_data = {{29'd0}, _GEN_215}; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_extra = auto_register_in_ar_valid ? auto_register_in_ar_bits_id : auto_register_in_aw_bits_id; // @[Decoupled.scala 289:21]
  assign Queue_io_deq_ready = _T_323_bits_read ? auto_register_in_r_ready : auto_register_in_b_ready; // @[Decoupled.scala 311:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  sels_0 = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  sels_1 = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  sels_2 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      sels_0 <= 3'h7;
    end else if (_T_179) begin
      sels_0 <= auto_register_in_w_bits_data[2:0];
    end
    if (reset) begin
      sels_1 <= 3'h7;
    end else if (_T_156) begin
      sels_1 <= auto_register_in_w_bits_data[2:0];
    end
    if (reset) begin
      sels_2 <= 3'h7;
    end else if (_T_133) begin
      sels_2 <= auto_register_in_w_bits_data[2:0];
    end
  end
endmodule
module AXI4Splitter_5(
  input         clock,
  input         reset,
  output        auto_mem_in_aw_ready,
  input         auto_mem_in_aw_valid,
  input         auto_mem_in_aw_bits_id,
  input  [29:0] auto_mem_in_aw_bits_addr,
  output        auto_mem_in_w_ready,
  input         auto_mem_in_w_valid,
  input  [31:0] auto_mem_in_w_bits_data,
  input  [3:0]  auto_mem_in_w_bits_strb,
  input         auto_mem_in_b_ready,
  output        auto_mem_in_b_valid,
  output        auto_mem_in_b_bits_id,
  output        auto_mem_in_ar_ready,
  input         auto_mem_in_ar_valid,
  input         auto_mem_in_ar_bits_id,
  input  [29:0] auto_mem_in_ar_bits_addr,
  input  [2:0]  auto_mem_in_ar_bits_size,
  input         auto_mem_in_r_ready,
  output        auto_mem_in_r_valid,
  output        auto_mem_in_r_bits_id,
  output [31:0] auto_mem_in_r_bits_data,
  output        auto_stream_in_ready,
  input         auto_stream_in_valid,
  input  [31:0] auto_stream_in_bits_data,
  input         auto_stream_in_bits_last,
  input         auto_stream_out_ready,
  output        auto_stream_out_valid,
  output [31:0] auto_stream_out_bits_data,
  output        auto_stream_out_bits_last
);
  wire  Queue_clock; // @[Decoupled.scala 287:21]
  wire  Queue_reset; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_read; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_enq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_extra; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_read; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_deq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_extra; // @[Decoupled.scala 287:21]
  reg [31:0] ctrlReg; // @[Splitter.scala 27:26]
  reg [31:0] _RAND_0;
  reg [31:0] maskReg; // @[Splitter.scala 28:26]
  reg [31:0] _RAND_1;
  wire  _T_3; // @[RegisterRouter.scala 40:39]
  wire  _T_4; // @[RegisterRouter.scala 40:26]
  wire  _T_5; // @[RegisterRouter.scala 42:29]
  wire  _T_48_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 290:17]
  wire [29:0] _T_12; // @[RegisterRouter.scala 48:19]
  wire [1:0] _T_52; // @[RegisterRouter.scala 59:16]
  wire  _T_54; // @[RegisterRouter.scala 59:16]
  wire  _T_6; // @[RegisterRouter.scala 42:26]
  wire [1:0] _T_15; // @[OneHot.scala 65:12]
  wire [1:0] _T_17; // @[Misc.scala 200:81]
  wire  _T_18; // @[Misc.scala 204:21]
  wire  _T_21; // @[Misc.scala 209:20]
  wire  _T_23; // @[Misc.scala 213:38]
  wire  _T_24; // @[Misc.scala 213:29]
  wire  _T_26; // @[Misc.scala 213:38]
  wire  _T_27; // @[Misc.scala 213:29]
  wire  _T_30; // @[Misc.scala 209:20]
  wire  _T_31; // @[Misc.scala 212:27]
  wire  _T_32; // @[Misc.scala 213:38]
  wire  _T_33; // @[Misc.scala 213:29]
  wire  _T_34; // @[Misc.scala 212:27]
  wire  _T_35; // @[Misc.scala 213:38]
  wire  _T_36; // @[Misc.scala 213:29]
  wire  _T_37; // @[Misc.scala 212:27]
  wire  _T_38; // @[Misc.scala 213:38]
  wire  _T_39; // @[Misc.scala 213:29]
  wire  _T_40; // @[Misc.scala 212:27]
  wire  _T_41; // @[Misc.scala 213:38]
  wire  _T_42; // @[Misc.scala 213:29]
  wire [3:0] _T_45; // @[Cat.scala 29:58]
  wire [3:0] _T_47; // @[RegisterRouter.scala 54:25]
  wire [7:0] _T_66; // @[Bitwise.scala 72:12]
  wire [7:0] _T_68; // @[Bitwise.scala 72:12]
  wire [7:0] _T_70; // @[Bitwise.scala 72:12]
  wire [7:0] _T_72; // @[Bitwise.scala 72:12]
  wire [31:0] _T_75; // @[Cat.scala 29:58]
  wire  _T_94; // @[RegisterRouter.scala 59:16]
  wire  _T_147; // @[RegisterRouter.scala 59:16]
  wire [1:0] _T_141; // @[OneHot.scala 58:35]
  wire  _T_164; // @[RegisterRouter.scala 59:16]
  wire  _T_171; // @[RegisterRouter.scala 59:16]
  wire  _T_172; // @[RegisterRouter.scala 59:16]
  wire  _T_101; // @[RegisterRouter.scala 59:16]
  wire  _T_166; // @[RegisterRouter.scala 59:16]
  wire  _T_167; // @[RegisterRouter.scala 59:16]
  wire  _T_124; // @[RegisterRouter.scala 59:16]
  wire  _GEN_11; // @[MuxLiteral.scala 48:10]
  wire [31:0] _GEN_13; // @[MuxLiteral.scala 48:10]
  wire  _T_222_bits_read; // @[Decoupled.scala 308:19 Decoupled.scala 309:14]
  wire  _T_222_valid; // @[Decoupled.scala 308:19 Decoupled.scala 310:15]
  wire  _T_225; // @[RegisterRouter.scala 65:29]
  wire  _T_228; // @[Splitter.scala 49:19]
  wire  _T_229; // @[Splitter.scala 52:24]
  wire  _GEN_14; // @[Splitter.scala 52:33]
  wire  _T_232; // @[Splitter.scala 62:34]
  Queue Queue ( // @[Decoupled.scala 287:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_read(Queue_io_enq_bits_read),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_extra(Queue_io_enq_bits_extra),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_read(Queue_io_deq_bits_read),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_extra(Queue_io_deq_bits_extra)
  );
  assign _T_3 = auto_mem_in_aw_valid & auto_mem_in_w_valid; // @[RegisterRouter.scala 40:39]
  assign _T_4 = auto_mem_in_ar_valid | _T_3; // @[RegisterRouter.scala 40:26]
  assign _T_5 = ~auto_mem_in_ar_valid; // @[RegisterRouter.scala 42:29]
  assign _T_48_ready = Queue_io_enq_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 290:17]
  assign _T_12 = auto_mem_in_ar_valid ? auto_mem_in_ar_bits_addr : auto_mem_in_aw_bits_addr; // @[RegisterRouter.scala 48:19]
  assign _T_52 = _T_12[3:2] & 2'h2; // @[RegisterRouter.scala 59:16]
  assign _T_54 = _T_52 == 2'h0; // @[RegisterRouter.scala 59:16]
  assign _T_6 = _T_48_ready & _T_5; // @[RegisterRouter.scala 42:26]
  assign _T_15 = 2'h1 << auto_mem_in_ar_bits_size[0]; // @[OneHot.scala 65:12]
  assign _T_17 = _T_15 | 2'h1; // @[Misc.scala 200:81]
  assign _T_18 = auto_mem_in_ar_bits_size >= 3'h2; // @[Misc.scala 204:21]
  assign _T_21 = ~auto_mem_in_ar_bits_addr[1]; // @[Misc.scala 209:20]
  assign _T_23 = _T_17[1] & _T_21; // @[Misc.scala 213:38]
  assign _T_24 = _T_18 | _T_23; // @[Misc.scala 213:29]
  assign _T_26 = _T_17[1] & auto_mem_in_ar_bits_addr[1]; // @[Misc.scala 213:38]
  assign _T_27 = _T_18 | _T_26; // @[Misc.scala 213:29]
  assign _T_30 = ~auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 209:20]
  assign _T_31 = _T_21 & _T_30; // @[Misc.scala 212:27]
  assign _T_32 = _T_17[0] & _T_31; // @[Misc.scala 213:38]
  assign _T_33 = _T_24 | _T_32; // @[Misc.scala 213:29]
  assign _T_34 = _T_21 & auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  assign _T_35 = _T_17[0] & _T_34; // @[Misc.scala 213:38]
  assign _T_36 = _T_24 | _T_35; // @[Misc.scala 213:29]
  assign _T_37 = auto_mem_in_ar_bits_addr[1] & _T_30; // @[Misc.scala 212:27]
  assign _T_38 = _T_17[0] & _T_37; // @[Misc.scala 213:38]
  assign _T_39 = _T_27 | _T_38; // @[Misc.scala 213:29]
  assign _T_40 = auto_mem_in_ar_bits_addr[1] & auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  assign _T_41 = _T_17[0] & _T_40; // @[Misc.scala 213:38]
  assign _T_42 = _T_27 | _T_41; // @[Misc.scala 213:29]
  assign _T_45 = {_T_42,_T_39,_T_36,_T_33}; // @[Cat.scala 29:58]
  assign _T_47 = auto_mem_in_ar_valid ? _T_45 : auto_mem_in_w_bits_strb; // @[RegisterRouter.scala 54:25]
  assign _T_66 = _T_47[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_68 = _T_47[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_70 = _T_47[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_72 = _T_47[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_75 = {_T_72,_T_70,_T_68,_T_66}; // @[Cat.scala 29:58]
  assign _T_94 = _T_75 == 32'hffffffff; // @[RegisterRouter.scala 59:16]
  assign _T_147 = _T_4 & _T_48_ready; // @[RegisterRouter.scala 59:16]
  assign _T_141 = 2'h1 << _T_12[2]; // @[OneHot.scala 58:35]
  assign _T_164 = _T_147 & _T_5; // @[RegisterRouter.scala 59:16]
  assign _T_171 = _T_164 & _T_141[1]; // @[RegisterRouter.scala 59:16]
  assign _T_172 = _T_171 & _T_54; // @[RegisterRouter.scala 59:16]
  assign _T_101 = _T_172 & _T_94; // @[RegisterRouter.scala 59:16]
  assign _T_166 = _T_164 & _T_141[0]; // @[RegisterRouter.scala 59:16]
  assign _T_167 = _T_166 & _T_54; // @[RegisterRouter.scala 59:16]
  assign _T_124 = _T_167 & _T_94; // @[RegisterRouter.scala 59:16]
  assign _GEN_11 = _T_12[2] ? _T_54 : _T_54; // @[MuxLiteral.scala 48:10]
  assign _GEN_13 = _T_12[2] ? maskReg : ctrlReg; // @[MuxLiteral.scala 48:10]
  assign _T_222_bits_read = Queue_io_deq_bits_read; // @[Decoupled.scala 308:19 Decoupled.scala 309:14]
  assign _T_222_valid = Queue_io_deq_valid; // @[Decoupled.scala 308:19 Decoupled.scala 310:15]
  assign _T_225 = ~_T_222_bits_read; // @[RegisterRouter.scala 65:29]
  assign _T_228 = ctrlReg == 32'h0; // @[Splitter.scala 49:19]
  assign _T_229 = ctrlReg == 32'h1; // @[Splitter.scala 52:24]
  assign _GEN_14 = _T_229 & auto_stream_out_ready; // @[Splitter.scala 52:33]
  assign _T_232 = ~maskReg[0]; // @[Splitter.scala 62:34]
  assign auto_mem_in_aw_ready = _T_6 & auto_mem_in_w_valid; // @[LazyModule.scala 173:31]
  assign auto_mem_in_w_ready = _T_6 & auto_mem_in_aw_valid; // @[LazyModule.scala 173:31]
  assign auto_mem_in_b_valid = _T_222_valid & _T_225; // @[LazyModule.scala 173:31]
  assign auto_mem_in_b_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_mem_in_ar_ready = Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_valid = _T_222_valid & _T_222_bits_read; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 173:31]
  assign auto_stream_in_ready = _T_228 ? auto_stream_out_ready : _GEN_14; // @[LazyModule.scala 173:31]
  assign auto_stream_out_valid = auto_stream_in_valid & _T_232; // @[LazyModule.scala 173:49]
  assign auto_stream_out_bits_data = auto_stream_in_bits_data; // @[LazyModule.scala 173:49]
  assign auto_stream_out_bits_last = auto_stream_in_bits_last; // @[LazyModule.scala 173:49]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_mem_in_ar_valid | _T_3; // @[Decoupled.scala 288:22]
  assign Queue_io_enq_bits_read = auto_mem_in_ar_valid; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_data = _GEN_11 ? _GEN_13 : 32'h0; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_extra = auto_mem_in_ar_valid ? auto_mem_in_ar_bits_id : auto_mem_in_aw_bits_id; // @[Decoupled.scala 289:21]
  assign Queue_io_deq_ready = _T_222_bits_read ? auto_mem_in_r_ready : auto_mem_in_b_ready; // @[Decoupled.scala 311:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ctrlReg = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  maskReg = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      ctrlReg <= 32'h0;
    end else if (_T_124) begin
      ctrlReg <= auto_mem_in_w_bits_data;
    end
    if (reset) begin
      maskReg <= 32'h0;
    end else if (_T_101) begin
      maskReg <= auto_mem_in_w_bits_data;
    end
  end
endmodule
module Queue_38(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [31:0] io_enq_bits_data,
  input         io_enq_bits_last,
  input         io_deq_ready,
  output        io_deq_valid,
  output [31:0] io_deq_bits_data,
  output        io_deq_bits_last
);
  reg [31:0] _T_data [0:0]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_0;
  wire [31:0] _T_data__T_14_data; // @[Decoupled.scala 209:24]
  wire  _T_data__T_14_addr; // @[Decoupled.scala 209:24]
  wire [31:0] _T_data__T_10_data; // @[Decoupled.scala 209:24]
  wire  _T_data__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T_data__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T_data__T_10_en; // @[Decoupled.scala 209:24]
  reg  _T_last [0:0]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_1;
  wire  _T_last__T_14_data; // @[Decoupled.scala 209:24]
  wire  _T_last__T_14_addr; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_data; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_en; // @[Decoupled.scala 209:24]
  reg  _T_1; // @[Decoupled.scala 212:35]
  reg [31:0] _RAND_2;
  wire  _T_3; // @[Decoupled.scala 215:36]
  wire  _T_6; // @[Decoupled.scala 40:37]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[Decoupled.scala 240:27]
  wire  _GEN_22; // @[Decoupled.scala 237:18]
  wire  _GEN_21; // @[Decoupled.scala 237:18]
  wire  _T_11; // @[Decoupled.scala 227:16]
  wire  _T_12; // @[Decoupled.scala 231:19]
  assign _T_data__T_14_addr = 1'h0;
  assign _T_data__T_14_data = _T_data[_T_data__T_14_addr]; // @[Decoupled.scala 209:24]
  assign _T_data__T_10_data = io_enq_bits_data;
  assign _T_data__T_10_addr = 1'h0;
  assign _T_data__T_10_mask = 1'h1;
  assign _T_data__T_10_en = _T_3 ? _GEN_13 : _T_6;
  assign _T_last__T_14_addr = 1'h0;
  assign _T_last__T_14_data = _T_last[_T_last__T_14_addr]; // @[Decoupled.scala 209:24]
  assign _T_last__T_10_data = io_enq_bits_last;
  assign _T_last__T_10_addr = 1'h0;
  assign _T_last__T_10_mask = 1'h1;
  assign _T_last__T_10_en = _T_3 ? _GEN_13 : _T_6;
  assign _T_3 = ~_T_1; // @[Decoupled.scala 215:36]
  assign _T_6 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  assign _T_8 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = io_deq_ready ? 1'h0 : _T_6; // @[Decoupled.scala 240:27]
  assign _GEN_22 = _T_3 ? _GEN_13 : _T_6; // @[Decoupled.scala 237:18]
  assign _GEN_21 = _T_3 ? 1'h0 : _T_8; // @[Decoupled.scala 237:18]
  assign _T_11 = _GEN_22 != _GEN_21; // @[Decoupled.scala 227:16]
  assign _T_12 = ~_T_3; // @[Decoupled.scala 231:19]
  assign io_enq_ready = io_deq_ready | _T_3; // @[Decoupled.scala 232:16 Decoupled.scala 245:40]
  assign io_deq_valid = io_enq_valid | _T_12; // @[Decoupled.scala 231:16 Decoupled.scala 236:40]
  assign io_deq_bits_data = _T_3 ? io_enq_bits_data : _T_data__T_14_data; // @[Decoupled.scala 233:15 Decoupled.scala 238:19]
  assign io_deq_bits_last = _T_3 ? io_enq_bits_last : _T_last__T_14_data; // @[Decoupled.scala 233:15 Decoupled.scala 238:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_data[initvar] = _RAND_0[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_last[initvar] = _RAND_1[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_1 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T_data__T_10_en & _T_data__T_10_mask) begin
      _T_data[_T_data__T_10_addr] <= _T_data__T_10_data; // @[Decoupled.scala 209:24]
    end
    if(_T_last__T_10_en & _T_last__T_10_mask) begin
      _T_last[_T_last__T_10_addr] <= _T_last__T_10_data; // @[Decoupled.scala 209:24]
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else if (_T_11) begin
      if (_T_3) begin
        if (io_deq_ready) begin
          _T_1 <= 1'h0;
        end else begin
          _T_1 <= _T_6;
        end
      end else begin
        _T_1 <= _T_6;
      end
    end
  end
endmodule
module StreamBuffer_2(
  input         clock,
  input         reset,
  input         auto_out_out_ready,
  output        auto_out_out_valid,
  output [31:0] auto_out_out_bits_data,
  output        auto_out_out_bits_last,
  output        auto_in_in_ready,
  input         auto_in_in_valid,
  input  [31:0] auto_in_in_bits_data,
  input         auto_in_in_bits_last
);
  wire  Queue_clock; // @[Decoupled.scala 287:21]
  wire  Queue_reset; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_enq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_last; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_deq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_last; // @[Decoupled.scala 287:21]
  Queue_38 Queue ( // @[Decoupled.scala 287:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_last(Queue_io_enq_bits_last),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_last(Queue_io_deq_bits_last)
  );
  assign auto_out_out_valid = Queue_io_deq_valid; // @[LazyModule.scala 173:49]
  assign auto_out_out_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_out_bits_last = Queue_io_deq_bits_last; // @[LazyModule.scala 173:49]
  assign auto_in_in_ready = Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_in_in_valid; // @[Decoupled.scala 288:22]
  assign Queue_io_enq_bits_data = auto_in_in_bits_data; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_last = auto_in_in_bits_last; // @[Decoupled.scala 289:21]
  assign Queue_io_deq_ready = auto_out_out_ready; // @[Decoupled.scala 311:15]
endmodule
module AXI4StreamWidthAdapater_1_to_4(
  input         clock,
  input         reset,
  output        auto_in_ready,
  input         auto_in_valid,
  input  [31:0] auto_in_bits_data,
  input         auto_in_bits_last,
  input         auto_out_ready,
  output        auto_out_valid,
  output [7:0]  auto_out_bits_data,
  output        auto_out_bits_last
);
  reg [1:0] _T_5; // @[AXI4StreamWidthAdapter.scala 158:22]
  reg [31:0] _RAND_0;
  wire  _T_6; // @[AXI4StreamWidthAdapter.scala 159:14]
  wire  _T_7; // @[AXI4StreamWidthAdapter.scala 159:38]
  wire [2:0] _T_8; // @[AXI4StreamWidthAdapter.scala 159:60]
  wire [2:0] _T_9; // @[AXI4StreamWidthAdapter.scala 159:33]
  wire [2:0] _GEN_0; // @[AXI4StreamWidthAdapter.scala 159:21]
  wire  ir0; // @[AXI4StreamWidthAdapter.scala 163:34]
  reg [1:0] _T_11; // @[AXI4StreamWidthAdapter.scala 167:22]
  reg [31:0] _RAND_1;
  wire  _T_13; // @[AXI4StreamWidthAdapter.scala 168:38]
  wire [2:0] _T_14; // @[AXI4StreamWidthAdapter.scala 168:60]
  wire [2:0] _T_15; // @[AXI4StreamWidthAdapter.scala 168:33]
  wire [2:0] _GEN_1; // @[AXI4StreamWidthAdapter.scala 168:21]
  wire  ir1; // @[AXI4StreamWidthAdapter.scala 170:60]
  reg [1:0] _T_20; // @[AXI4StreamWidthAdapter.scala 158:22]
  reg [31:0] _RAND_2;
  wire  _T_22; // @[AXI4StreamWidthAdapter.scala 159:38]
  wire [2:0] _T_23; // @[AXI4StreamWidthAdapter.scala 159:60]
  wire [2:0] _T_24; // @[AXI4StreamWidthAdapter.scala 159:33]
  wire [2:0] _GEN_2; // @[AXI4StreamWidthAdapter.scala 159:21]
  wire  ir2; // @[AXI4StreamWidthAdapter.scala 163:34]
  reg [1:0] _T_27; // @[AXI4StreamWidthAdapter.scala 158:22]
  reg [31:0] _RAND_3;
  wire  _T_29; // @[AXI4StreamWidthAdapter.scala 159:38]
  wire [2:0] _T_30; // @[AXI4StreamWidthAdapter.scala 159:60]
  wire [2:0] _T_31; // @[AXI4StreamWidthAdapter.scala 159:33]
  wire [2:0] _GEN_3; // @[AXI4StreamWidthAdapter.scala 159:21]
  wire  ir3; // @[AXI4StreamWidthAdapter.scala 163:34]
  reg [1:0] _T_34; // @[AXI4StreamWidthAdapter.scala 158:22]
  reg [31:0] _RAND_4;
  wire  _T_36; // @[AXI4StreamWidthAdapter.scala 159:38]
  wire [2:0] _T_37; // @[AXI4StreamWidthAdapter.scala 159:60]
  wire [2:0] _T_38; // @[AXI4StreamWidthAdapter.scala 159:33]
  wire [2:0] _GEN_4; // @[AXI4StreamWidthAdapter.scala 159:21]
  wire  ir4; // @[AXI4StreamWidthAdapter.scala 163:34]
  wire  _T_56; // @[AXI4StreamWidthAdapter.scala 46:16]
  wire  _T_58; // @[AXI4StreamWidthAdapter.scala 46:11]
  wire  _T_59; // @[AXI4StreamWidthAdapter.scala 46:11]
  wire  _T_60; // @[AXI4StreamWidthAdapter.scala 47:16]
  wire  _T_62; // @[AXI4StreamWidthAdapter.scala 47:11]
  wire  _T_63; // @[AXI4StreamWidthAdapter.scala 47:11]
  wire  _T_64; // @[AXI4StreamWidthAdapter.scala 48:16]
  wire  _T_66; // @[AXI4StreamWidthAdapter.scala 48:11]
  wire  _T_67; // @[AXI4StreamWidthAdapter.scala 48:11]
  wire  _T_68; // @[AXI4StreamWidthAdapter.scala 49:16]
  wire  _T_70; // @[AXI4StreamWidthAdapter.scala 49:11]
  wire  _T_71; // @[AXI4StreamWidthAdapter.scala 49:11]
  wire [7:0] _GEN_6; // @[AXI4StreamWidthAdapter.scala 54:19]
  wire [7:0] _GEN_7; // @[AXI4StreamWidthAdapter.scala 54:19]
  assign _T_6 = auto_in_valid & auto_out_ready; // @[AXI4StreamWidthAdapter.scala 159:14]
  assign _T_7 = _T_5 == 2'h3; // @[AXI4StreamWidthAdapter.scala 159:38]
  assign _T_8 = _T_5 + 2'h1; // @[AXI4StreamWidthAdapter.scala 159:60]
  assign _T_9 = _T_7 ? 3'h0 : _T_8; // @[AXI4StreamWidthAdapter.scala 159:33]
  assign _GEN_0 = _T_6 ? _T_9 : {{1'd0}, _T_5}; // @[AXI4StreamWidthAdapter.scala 159:21]
  assign ir0 = _T_7 & auto_out_ready; // @[AXI4StreamWidthAdapter.scala 163:34]
  assign _T_13 = _T_11 == 2'h3; // @[AXI4StreamWidthAdapter.scala 168:38]
  assign _T_14 = _T_11 + 2'h1; // @[AXI4StreamWidthAdapter.scala 168:60]
  assign _T_15 = _T_13 ? 3'h0 : _T_14; // @[AXI4StreamWidthAdapter.scala 168:33]
  assign _GEN_1 = _T_6 ? _T_15 : {{1'd0}, _T_11}; // @[AXI4StreamWidthAdapter.scala 168:21]
  assign ir1 = _T_13 & auto_out_ready; // @[AXI4StreamWidthAdapter.scala 170:60]
  assign _T_22 = _T_20 == 2'h3; // @[AXI4StreamWidthAdapter.scala 159:38]
  assign _T_23 = _T_20 + 2'h1; // @[AXI4StreamWidthAdapter.scala 159:60]
  assign _T_24 = _T_22 ? 3'h0 : _T_23; // @[AXI4StreamWidthAdapter.scala 159:33]
  assign _GEN_2 = _T_6 ? _T_24 : {{1'd0}, _T_20}; // @[AXI4StreamWidthAdapter.scala 159:21]
  assign ir2 = _T_22 & auto_out_ready; // @[AXI4StreamWidthAdapter.scala 163:34]
  assign _T_29 = _T_27 == 2'h3; // @[AXI4StreamWidthAdapter.scala 159:38]
  assign _T_30 = _T_27 + 2'h1; // @[AXI4StreamWidthAdapter.scala 159:60]
  assign _T_31 = _T_29 ? 3'h0 : _T_30; // @[AXI4StreamWidthAdapter.scala 159:33]
  assign _GEN_3 = _T_6 ? _T_31 : {{1'd0}, _T_27}; // @[AXI4StreamWidthAdapter.scala 159:21]
  assign ir3 = _T_29 & auto_out_ready; // @[AXI4StreamWidthAdapter.scala 163:34]
  assign _T_36 = _T_34 == 2'h3; // @[AXI4StreamWidthAdapter.scala 159:38]
  assign _T_37 = _T_34 + 2'h1; // @[AXI4StreamWidthAdapter.scala 159:60]
  assign _T_38 = _T_36 ? 3'h0 : _T_37; // @[AXI4StreamWidthAdapter.scala 159:33]
  assign _GEN_4 = _T_6 ? _T_38 : {{1'd0}, _T_34}; // @[AXI4StreamWidthAdapter.scala 159:21]
  assign ir4 = _T_36 & auto_out_ready; // @[AXI4StreamWidthAdapter.scala 163:34]
  assign _T_56 = ir0 == ir1; // @[AXI4StreamWidthAdapter.scala 46:16]
  assign _T_58 = _T_56 | reset; // @[AXI4StreamWidthAdapter.scala 46:11]
  assign _T_59 = ~_T_58; // @[AXI4StreamWidthAdapter.scala 46:11]
  assign _T_60 = ir0 == ir2; // @[AXI4StreamWidthAdapter.scala 47:16]
  assign _T_62 = _T_60 | reset; // @[AXI4StreamWidthAdapter.scala 47:11]
  assign _T_63 = ~_T_62; // @[AXI4StreamWidthAdapter.scala 47:11]
  assign _T_64 = ir0 == ir3; // @[AXI4StreamWidthAdapter.scala 48:16]
  assign _T_66 = _T_64 | reset; // @[AXI4StreamWidthAdapter.scala 48:11]
  assign _T_67 = ~_T_66; // @[AXI4StreamWidthAdapter.scala 48:11]
  assign _T_68 = ir0 == ir4; // @[AXI4StreamWidthAdapter.scala 49:16]
  assign _T_70 = _T_68 | reset; // @[AXI4StreamWidthAdapter.scala 49:11]
  assign _T_71 = ~_T_70; // @[AXI4StreamWidthAdapter.scala 49:11]
  assign _GEN_6 = 2'h1 == _T_5 ? auto_in_bits_data[15:8] : auto_in_bits_data[7:0]; // @[AXI4StreamWidthAdapter.scala 54:19]
  assign _GEN_7 = 2'h2 == _T_5 ? auto_in_bits_data[23:16] : _GEN_6; // @[AXI4StreamWidthAdapter.scala 54:19]
  assign auto_in_ready = _T_7 & auto_out_ready; // @[LazyModule.scala 173:31]
  assign auto_out_valid = auto_in_valid; // @[LazyModule.scala 173:49]
  assign auto_out_bits_data = 2'h3 == _T_5 ? auto_in_bits_data[31:24] : _GEN_7; // @[LazyModule.scala 173:49]
  assign auto_out_bits_last = auto_in_bits_last & _T_13; // @[LazyModule.scala 173:49]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_5 = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_11 = _RAND_1[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_20 = _RAND_2[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_27 = _RAND_3[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_34 = _RAND_4[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      _T_5 <= 2'h0;
    end else begin
      _T_5 <= _GEN_0[1:0];
    end
    if (reset) begin
      _T_11 <= 2'h0;
    end else begin
      _T_11 <= _GEN_1[1:0];
    end
    if (reset) begin
      _T_20 <= 2'h0;
    end else begin
      _T_20 <= _GEN_2[1:0];
    end
    if (reset) begin
      _T_27 <= 2'h0;
    end else begin
      _T_27 <= _GEN_3[1:0];
    end
    if (reset) begin
      _T_34 <= 2'h0;
    end else begin
      _T_34 <= _GEN_4[1:0];
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_59) begin
          $fwrite(32'h80000002,"Assertion failed\n    at AXI4StreamWidthAdapter.scala:46 assert(ir0 === ir1)\n"); // @[AXI4StreamWidthAdapter.scala 46:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_59) begin
          $fatal; // @[AXI4StreamWidthAdapter.scala 46:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_63) begin
          $fwrite(32'h80000002,"Assertion failed\n    at AXI4StreamWidthAdapter.scala:47 assert(ir0 === ir2)\n"); // @[AXI4StreamWidthAdapter.scala 47:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_63) begin
          $fatal; // @[AXI4StreamWidthAdapter.scala 47:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_67) begin
          $fwrite(32'h80000002,"Assertion failed\n    at AXI4StreamWidthAdapter.scala:48 assert(ir0 === ir3)\n"); // @[AXI4StreamWidthAdapter.scala 48:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_67) begin
          $fatal; // @[AXI4StreamWidthAdapter.scala 48:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_71) begin
          $fwrite(32'h80000002,"Assertion failed\n    at AXI4StreamWidthAdapter.scala:49 assert(ir0 === ir4)\n"); // @[AXI4StreamWidthAdapter.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_71) begin
          $fatal; // @[AXI4StreamWidthAdapter.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module Queue_39(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [31:0] io_enq_bits_data,
  input         io_enq_bits_last,
  input         io_deq_ready,
  output        io_deq_valid,
  output [31:0] io_deq_bits_data,
  output        io_deq_bits_last
);
  reg [31:0] _T_data [0:3]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_0;
  wire [31:0] _T_data__T_18_data; // @[Decoupled.scala 209:24]
  wire [1:0] _T_data__T_18_addr; // @[Decoupled.scala 209:24]
  wire [31:0] _T_data__T_10_data; // @[Decoupled.scala 209:24]
  wire [1:0] _T_data__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T_data__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T_data__T_10_en; // @[Decoupled.scala 209:24]
  reg  _T_last [0:3]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_1;
  wire  _T_last__T_18_data; // @[Decoupled.scala 209:24]
  wire [1:0] _T_last__T_18_addr; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_data; // @[Decoupled.scala 209:24]
  wire [1:0] _T_last__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_en; // @[Decoupled.scala 209:24]
  reg [1:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_2;
  reg [1:0] value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_3;
  reg  _T_1; // @[Decoupled.scala 212:35]
  reg [31:0] _RAND_4;
  wire  _T_2; // @[Decoupled.scala 214:41]
  wire  _T_3; // @[Decoupled.scala 215:36]
  wire  _T_4; // @[Decoupled.scala 215:33]
  wire  _T_5; // @[Decoupled.scala 216:32]
  wire  _T_6; // @[Decoupled.scala 40:37]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire [1:0] _T_12; // @[Counter.scala 39:22]
  wire [1:0] _T_14; // @[Counter.scala 39:22]
  wire  _T_15; // @[Decoupled.scala 227:16]
  assign _T_data__T_18_addr = value_1;
  assign _T_data__T_18_data = _T_data[_T_data__T_18_addr]; // @[Decoupled.scala 209:24]
  assign _T_data__T_10_data = io_enq_bits_data;
  assign _T_data__T_10_addr = value;
  assign _T_data__T_10_mask = 1'h1;
  assign _T_data__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_last__T_18_addr = value_1;
  assign _T_last__T_18_data = _T_last[_T_last__T_18_addr]; // @[Decoupled.scala 209:24]
  assign _T_last__T_10_data = io_enq_bits_last;
  assign _T_last__T_10_addr = value;
  assign _T_last__T_10_mask = 1'h1;
  assign _T_last__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_2 = value == value_1; // @[Decoupled.scala 214:41]
  assign _T_3 = ~_T_1; // @[Decoupled.scala 215:36]
  assign _T_4 = _T_2 & _T_3; // @[Decoupled.scala 215:33]
  assign _T_5 = _T_2 & _T_1; // @[Decoupled.scala 216:32]
  assign _T_6 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  assign _T_8 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  assign _T_12 = value + 2'h1; // @[Counter.scala 39:22]
  assign _T_14 = value_1 + 2'h1; // @[Counter.scala 39:22]
  assign _T_15 = _T_6 != _T_8; // @[Decoupled.scala 227:16]
  assign io_enq_ready = ~_T_5; // @[Decoupled.scala 232:16]
  assign io_deq_valid = ~_T_4; // @[Decoupled.scala 231:16]
  assign io_deq_bits_data = _T_data__T_18_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_last = _T_last__T_18_data; // @[Decoupled.scala 233:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    _T_data[initvar] = _RAND_0[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    _T_last[initvar] = _RAND_1[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  value = _RAND_2[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  value_1 = _RAND_3[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T_data__T_10_en & _T_data__T_10_mask) begin
      _T_data[_T_data__T_10_addr] <= _T_data__T_10_data; // @[Decoupled.scala 209:24]
    end
    if(_T_last__T_10_en & _T_last__T_10_mask) begin
      _T_last[_T_last__T_10_addr] <= _T_last__T_10_data; // @[Decoupled.scala 209:24]
    end
    if (reset) begin
      value <= 2'h0;
    end else if (_T_6) begin
      value <= _T_12;
    end
    if (reset) begin
      value_1 <= 2'h0;
    end else if (_T_8) begin
      value_1 <= _T_14;
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else if (_T_15) begin
      _T_1 <= _T_6;
    end
  end
endmodule
module StreamBuffer_3(
  input         clock,
  input         reset,
  input         auto_out_out_ready,
  output        auto_out_out_valid,
  output [31:0] auto_out_out_bits_data,
  output        auto_out_out_bits_last,
  output        auto_in_in_ready,
  input         auto_in_in_valid,
  input  [31:0] auto_in_in_bits_data,
  input         auto_in_in_bits_last
);
  wire  Queue_clock; // @[Decoupled.scala 287:21]
  wire  Queue_reset; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_enq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_last; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_deq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_last; // @[Decoupled.scala 287:21]
  Queue_39 Queue ( // @[Decoupled.scala 287:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_last(Queue_io_enq_bits_last),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_last(Queue_io_deq_bits_last)
  );
  assign auto_out_out_valid = Queue_io_deq_valid; // @[LazyModule.scala 173:49]
  assign auto_out_out_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_out_bits_last = Queue_io_deq_bits_last; // @[LazyModule.scala 173:49]
  assign auto_in_in_ready = Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_in_in_valid; // @[Decoupled.scala 288:22]
  assign Queue_io_enq_bits_data = auto_in_in_bits_data; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_last = auto_in_in_bits_last; // @[Decoupled.scala 289:21]
  assign Queue_io_deq_ready = auto_out_out_ready; // @[Decoupled.scala 311:15]
endmodule
module IntToBundleBridge(
  input   auto_in_0,
  output  auto_out_0
);
  assign auto_out_0 = auto_in_0; // @[LazyModule.scala 173:49]
endmodule
module UARTTx(
  input         clock,
  input         reset,
  input         io_en,
  output        io_in_ready,
  input         io_in_valid,
  input  [7:0]  io_in_bits,
  output        io_out,
  input  [15:0] io_div,
  input         io_nstop
);
  wire [31:0] plusarg_reader_out; // @[PlusArg.scala 44:11]
  reg [15:0] prescaler; // @[UARTTx.scala 21:22]
  reg [31:0] _RAND_0;
  wire  pulse; // @[UARTTx.scala 22:26]
  reg [3:0] counter; // @[UARTTx.scala 25:20]
  reg [31:0] _RAND_1;
  reg [8:0] shifter; // @[UARTTx.scala 26:20]
  reg [31:0] _RAND_2;
  reg  out; // @[UARTTx.scala 27:16]
  reg [31:0] _RAND_3;
  wire  plusarg_tx; // @[UARTTx.scala 30:90]
  wire  busy; // @[UARTTx.scala 32:23]
  wire  _T; // @[UARTTx.scala 33:27]
  wire  _T_2; // @[Decoupled.scala 40:37]
  wire  _T_4; // @[UARTTx.scala 36:11]
  wire  _T_6; // @[UARTTx.scala 38:22]
  wire [9:0] _T_9; // @[Cat.scala 29:58]
  wire  _T_10; // @[UARTTx.scala 55:19]
  wire [3:0] _T_12; // @[Mux.scala 27:72]
  wire [3:0] _T_13; // @[Mux.scala 27:72]
  wire [3:0] _T_14; // @[Mux.scala 27:72]
  wire [3:0] _T_17; // @[UARTTx.scala 55:53]
  wire [9:0] _GEN_0; // @[UARTTx.scala 38:37]
  wire [15:0] _T_20; // @[UARTTx.scala 59:78]
  wire  _T_22; // @[UARTTx.scala 61:15]
  wire [3:0] _T_24; // @[UARTTx.scala 62:24]
  wire [8:0] _T_26; // @[Cat.scala 29:58]
  wire [9:0] _GEN_4; // @[UARTTx.scala 61:24]
  wire  _GEN_5; // @[UARTTx.scala 61:24]
  plusarg_reader #(.FORMAT("uart_tx=%d"), .DEFAULT(1), .WIDTH(32)) plusarg_reader ( // @[PlusArg.scala 44:11]
    .out(plusarg_reader_out)
  );
  assign pulse = prescaler == 16'h0; // @[UARTTx.scala 22:26]
  assign plusarg_tx = plusarg_reader_out != 32'h0; // @[UARTTx.scala 30:90]
  assign busy = counter != 4'h0; // @[UARTTx.scala 32:23]
  assign _T = ~busy; // @[UARTTx.scala 33:27]
  assign _T_2 = io_in_ready & io_in_valid; // @[Decoupled.scala 40:37]
  assign _T_4 = ~reset; // @[UARTTx.scala 36:11]
  assign _T_6 = _T_2 & plusarg_tx; // @[UARTTx.scala 38:22]
  assign _T_9 = {1'h1,io_in_bits,1'h0}; // @[Cat.scala 29:58]
  assign _T_10 = ~io_nstop; // @[UARTTx.scala 55:19]
  assign _T_12 = _T_10 ? 4'ha : 4'h0; // @[Mux.scala 27:72]
  assign _T_13 = io_nstop ? 4'hb : 4'h0; // @[Mux.scala 27:72]
  assign _T_14 = _T_12 | _T_13; // @[Mux.scala 27:72]
  assign _T_17 = _T_14 - 4'h0; // @[UARTTx.scala 55:53]
  assign _GEN_0 = _T_6 ? _T_9 : {{1'd0}, shifter}; // @[UARTTx.scala 38:37]
  assign _T_20 = prescaler - 16'h1; // @[UARTTx.scala 59:78]
  assign _T_22 = pulse & busy; // @[UARTTx.scala 61:15]
  assign _T_24 = counter - 4'h1; // @[UARTTx.scala 62:24]
  assign _T_26 = {1'h1,shifter[8:1]}; // @[Cat.scala 29:58]
  assign _GEN_4 = _T_22 ? {{1'd0}, _T_26} : _GEN_0; // @[UARTTx.scala 61:24]
  assign _GEN_5 = _T_22 ? shifter[0] : out; // @[UARTTx.scala 61:24]
  assign io_in_ready = io_en & _T; // @[UARTTx.scala 33:15]
  assign io_out = out; // @[UARTTx.scala 28:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  prescaler = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  counter = _RAND_1[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  shifter = _RAND_2[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      prescaler <= 16'h0;
    end else if (busy) begin
      if (pulse) begin
        prescaler <= io_div;
      end else begin
        prescaler <= _T_20;
      end
    end
    if (reset) begin
      counter <= 4'h0;
    end else if (_T_22) begin
      counter <= _T_24;
    end else if (_T_6) begin
      counter <= _T_17;
    end
    shifter <= _GEN_4[8:0];
    out <= reset | _GEN_5;
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & _T_4) begin
          $fwrite(32'h80000002,"UART TX (%x): %c\n",io_in_bits,io_in_bits); // @[UARTTx.scala 36:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module QueueCompatibility_6(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input  [7:0] io_enq_bits,
  input        io_deq_ready,
  output       io_deq_valid,
  output [7:0] io_deq_bits,
  output [8:0] io_count
);
  reg [7:0] _T [0:255]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_0;
  wire [7:0] _T__T_18_data; // @[Decoupled.scala 209:24]
  wire [7:0] _T__T_18_addr; // @[Decoupled.scala 209:24]
  wire [7:0] _T__T_10_data; // @[Decoupled.scala 209:24]
  wire [7:0] _T__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T__T_10_en; // @[Decoupled.scala 209:24]
  reg [7:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_1;
  reg [7:0] value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_2;
  reg  _T_1; // @[Decoupled.scala 212:35]
  reg [31:0] _RAND_3;
  wire  _T_2; // @[Decoupled.scala 214:41]
  wire  _T_3; // @[Decoupled.scala 215:36]
  wire  _T_4; // @[Decoupled.scala 215:33]
  wire  _T_5; // @[Decoupled.scala 216:32]
  wire  _T_6; // @[Decoupled.scala 40:37]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire [7:0] _T_12; // @[Counter.scala 39:22]
  wire [7:0] _T_14; // @[Counter.scala 39:22]
  wire  _T_15; // @[Decoupled.scala 227:16]
  wire [7:0] _T_20; // @[Decoupled.scala 248:40]
  wire  _T_21; // @[Decoupled.scala 250:32]
  wire [8:0] _T_22; // @[Decoupled.scala 250:20]
  wire [8:0] _GEN_8; // @[Decoupled.scala 250:62]
  assign _T__T_18_addr = value_1;
  assign _T__T_18_data = _T[_T__T_18_addr]; // @[Decoupled.scala 209:24]
  assign _T__T_10_data = io_enq_bits;
  assign _T__T_10_addr = value;
  assign _T__T_10_mask = 1'h1;
  assign _T__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_2 = value == value_1; // @[Decoupled.scala 214:41]
  assign _T_3 = ~_T_1; // @[Decoupled.scala 215:36]
  assign _T_4 = _T_2 & _T_3; // @[Decoupled.scala 215:33]
  assign _T_5 = _T_2 & _T_1; // @[Decoupled.scala 216:32]
  assign _T_6 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  assign _T_8 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  assign _T_12 = value + 8'h1; // @[Counter.scala 39:22]
  assign _T_14 = value_1 + 8'h1; // @[Counter.scala 39:22]
  assign _T_15 = _T_6 != _T_8; // @[Decoupled.scala 227:16]
  assign _T_20 = value - value_1; // @[Decoupled.scala 248:40]
  assign _T_21 = _T_1 & _T_2; // @[Decoupled.scala 250:32]
  assign _T_22 = _T_21 ? 9'h100 : 9'h0; // @[Decoupled.scala 250:20]
  assign _GEN_8 = {{1'd0}, _T_20}; // @[Decoupled.scala 250:62]
  assign io_enq_ready = ~_T_5; // @[Decoupled.scala 232:16]
  assign io_deq_valid = ~_T_4; // @[Decoupled.scala 231:16]
  assign io_deq_bits = _T__T_18_data; // @[Decoupled.scala 233:15]
  assign io_count = _T_22 | _GEN_8; // @[Decoupled.scala 250:14]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    _T[initvar] = _RAND_0[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  value = _RAND_1[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  value_1 = _RAND_2[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_1 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T__T_10_en & _T__T_10_mask) begin
      _T[_T__T_10_addr] <= _T__T_10_data; // @[Decoupled.scala 209:24]
    end
    if (reset) begin
      value <= 8'h0;
    end else if (_T_6) begin
      value <= _T_12;
    end
    if (reset) begin
      value_1 <= 8'h0;
    end else if (_T_8) begin
      value_1 <= _T_14;
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else if (_T_15) begin
      _T_1 <= _T_6;
    end
  end
endmodule
module UARTRx(
  input         clock,
  input         reset,
  input         io_en,
  input         io_in,
  output        io_out_valid,
  output [7:0]  io_out_bits,
  input  [15:0] io_div
);
  reg [1:0] debounce; // @[UARTRx.scala 22:21]
  reg [31:0] _RAND_0;
  wire  debounce_max; // @[UARTRx.scala 23:32]
  wire  debounce_min; // @[UARTRx.scala 24:32]
  reg [12:0] prescaler; // @[UARTRx.scala 26:22]
  reg [31:0] _RAND_1;
  wire  pulse; // @[UARTRx.scala 28:26]
  reg [3:0] data_count; // @[UARTRx.scala 32:23]
  reg [31:0] _RAND_2;
  wire  data_last; // @[UARTRx.scala 33:31]
  reg [3:0] sample_count; // @[UARTRx.scala 35:25]
  reg [31:0] _RAND_3;
  wire  sample_mid; // @[UARTRx.scala 36:34]
  wire [7:0] _T_1; // @[Cat.scala 29:58]
  wire [7:0] countdown; // @[UARTRx.scala 38:49]
  wire [3:0] remainder; // @[UARTRx.scala 43:25]
  wire  extend; // @[UARTRx.scala 44:30]
  reg  state; // @[UARTRx.scala 59:18]
  reg [31:0] _RAND_4;
  wire  _T_14; // @[Conditional.scala 37:30]
  wire  _T_21; // @[UARTRx.scala 66:13]
  wire  _GEN_8; // @[UARTRx.scala 66:21]
  wire  start; // @[Conditional.scala 40:58]
  wire  restore; // @[UARTRx.scala 45:23]
  wire [12:0] prescaler_in; // @[UARTRx.scala 46:25]
  wire  _T_4; // @[UARTRx.scala 47:51]
  wire  _T_5; // @[UARTRx.scala 47:42]
  wire [12:0] _GEN_41; // @[UARTRx.scala 47:37]
  wire [12:0] prescaler_next; // @[UARTRx.scala 47:37]
  reg [2:0] sample; // @[UARTRx.scala 49:19]
  reg [31:0] _RAND_5;
  wire  _T_10; // @[Misc.scala 165:48]
  wire  _T_11; // @[Misc.scala 165:48]
  wire  _T_12; // @[Misc.scala 166:22]
  wire  _T_13; // @[Misc.scala 165:48]
  wire  voter; // @[Misc.scala 166:22]
  reg [7:0] shifter; // @[UARTRx.scala 51:20]
  reg [31:0] _RAND_6;
  reg  valid; // @[UARTRx.scala 53:18]
  reg [31:0] _RAND_7;
  wire  _T_16; // @[UARTRx.scala 63:13]
  wire  _T_17; // @[UARTRx.scala 63:26]
  wire  _T_18; // @[UARTRx.scala 63:23]
  wire [1:0] _T_20; // @[UARTRx.scala 64:30]
  wire [1:0] _T_23; // @[UARTRx.scala 67:30]
  wire [3:0] _T_27; // @[UARTRx.scala 72:94]
  wire  _GEN_1; // @[UARTRx.scala 68:29]
  wire [3:0] _T_29; // @[Cat.scala 29:58]
  wire [7:0] _T_33; // @[Cat.scala 29:58]
  wire  _GEN_16; // @[UARTRx.scala 85:27]
  wire [3:0] _GEN_18; // @[UARTRx.scala 80:20]
  wire  _GEN_22; // @[UARTRx.scala 80:20]
  wire [3:0] _GEN_25; // @[Conditional.scala 39:67]
  wire  _GEN_29; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_37; // @[Conditional.scala 40:58]
  wire  _T_34; // @[UARTRx.scala 112:9]
  assign debounce_max = debounce == 2'h3; // @[UARTRx.scala 23:32]
  assign debounce_min = debounce == 2'h0; // @[UARTRx.scala 24:32]
  assign pulse = prescaler == 13'h0; // @[UARTRx.scala 28:26]
  assign data_last = data_count == 4'h0; // @[UARTRx.scala 33:31]
  assign sample_mid = sample_count == 4'h7; // @[UARTRx.scala 36:34]
  assign _T_1 = {data_count,sample_count}; // @[Cat.scala 29:58]
  assign countdown = _T_1 - 8'h1; // @[UARTRx.scala 38:49]
  assign remainder = io_div[3:0]; // @[UARTRx.scala 43:25]
  assign extend = sample_count < remainder; // @[UARTRx.scala 44:30]
  assign _T_14 = ~state; // @[Conditional.scala 37:30]
  assign _T_21 = ~io_in; // @[UARTRx.scala 66:13]
  assign _GEN_8 = _T_21 & debounce_max; // @[UARTRx.scala 66:21]
  assign start = _T_14 & _GEN_8; // @[Conditional.scala 40:58]
  assign restore = start | pulse; // @[UARTRx.scala 45:23]
  assign prescaler_in = restore ? {{1'd0}, io_div[15:4]} : prescaler; // @[UARTRx.scala 46:25]
  assign _T_4 = restore & extend; // @[UARTRx.scala 47:51]
  assign _T_5 = _T_4 ? 1'h0 : 1'h1; // @[UARTRx.scala 47:42]
  assign _GEN_41 = {{12'd0}, _T_5}; // @[UARTRx.scala 47:37]
  assign prescaler_next = prescaler_in - _GEN_41; // @[UARTRx.scala 47:37]
  assign _T_10 = sample[0] & sample[1]; // @[Misc.scala 165:48]
  assign _T_11 = sample[0] & sample[2]; // @[Misc.scala 165:48]
  assign _T_12 = _T_10 | _T_11; // @[Misc.scala 166:22]
  assign _T_13 = sample[1] & sample[2]; // @[Misc.scala 165:48]
  assign voter = _T_12 | _T_13; // @[Misc.scala 166:22]
  assign _T_16 = ~_T_21; // @[UARTRx.scala 63:13]
  assign _T_17 = ~debounce_min; // @[UARTRx.scala 63:26]
  assign _T_18 = _T_16 & _T_17; // @[UARTRx.scala 63:23]
  assign _T_20 = debounce - 2'h1; // @[UARTRx.scala 64:30]
  assign _T_23 = debounce + 2'h1; // @[UARTRx.scala 67:30]
  assign _T_27 = 4'h9 - 4'h0; // @[UARTRx.scala 72:94]
  assign _GEN_1 = debounce_max | state; // @[UARTRx.scala 68:29]
  assign _T_29 = {sample,io_in}; // @[Cat.scala 29:58]
  assign _T_33 = {voter,shifter[7:1]}; // @[Cat.scala 29:58]
  assign _GEN_16 = sample_mid & data_last; // @[UARTRx.scala 85:27]
  assign _GEN_18 = pulse ? _T_29 : {{1'd0}, sample}; // @[UARTRx.scala 80:20]
  assign _GEN_22 = pulse & _GEN_16; // @[UARTRx.scala 80:20]
  assign _GEN_25 = state ? _GEN_18 : {{1'd0}, sample}; // @[Conditional.scala 39:67]
  assign _GEN_29 = state & _GEN_22; // @[Conditional.scala 39:67]
  assign _GEN_37 = _T_14 ? {{1'd0}, sample} : _GEN_25; // @[Conditional.scala 40:58]
  assign _T_34 = ~io_en; // @[UARTRx.scala 112:9]
  assign io_out_valid = valid; // @[UARTRx.scala 55:16]
  assign io_out_bits = shifter; // @[UARTRx.scala 56:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  debounce = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  prescaler = _RAND_1[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  data_count = _RAND_2[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  sample_count = _RAND_3[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  state = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  sample = _RAND_5[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  shifter = _RAND_6[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  valid = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      debounce <= 2'h0;
    end else if (_T_34) begin
      debounce <= 2'h0;
    end else if (_T_14) begin
      if (_T_21) begin
        debounce <= _T_23;
      end else if (_T_18) begin
        debounce <= _T_20;
      end
    end
    if (_T_14) begin
      if (_T_21) begin
        if (debounce_max) begin
          prescaler <= prescaler_next;
        end
      end
    end else if (state) begin
      prescaler <= prescaler_next;
    end
    if (_T_14) begin
      if (_T_21) begin
        if (debounce_max) begin
          data_count <= _T_27;
        end
      end
    end else if (state) begin
      if (pulse) begin
        data_count <= countdown[7:4];
      end
    end
    if (_T_14) begin
      if (_T_21) begin
        if (debounce_max) begin
          sample_count <= 4'hf;
        end
      end
    end else if (state) begin
      if (pulse) begin
        sample_count <= countdown[3:0];
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else if (_T_14) begin
      if (_T_21) begin
        state <= _GEN_1;
      end
    end else if (state) begin
      if (pulse) begin
        if (sample_mid) begin
          if (data_last) begin
            state <= 1'h0;
          end
        end
      end
    end
    sample <= _GEN_37[2:0];
    if (!(_T_14)) begin
      if (state) begin
        if (pulse) begin
          if (sample_mid) begin
            if (!(data_last)) begin
              shifter <= _T_33;
            end
          end
        end
      end
    end
    if (reset) begin
      valid <= 1'h0;
    end else if (_T_14) begin
      valid <= 1'h0;
    end else begin
      valid <= _GEN_29;
    end
  end
endmodule
module AXI4UARTBlock(
  input         clock,
  input         reset,
  output        auto_mem_in_aw_ready,
  input         auto_mem_in_aw_valid,
  input         auto_mem_in_aw_bits_id,
  input  [29:0] auto_mem_in_aw_bits_addr,
  output        auto_mem_in_w_ready,
  input         auto_mem_in_w_valid,
  input  [31:0] auto_mem_in_w_bits_data,
  input  [3:0]  auto_mem_in_w_bits_strb,
  input         auto_mem_in_b_ready,
  output        auto_mem_in_b_valid,
  output        auto_mem_in_b_bits_id,
  output        auto_mem_in_ar_ready,
  input         auto_mem_in_ar_valid,
  input         auto_mem_in_ar_bits_id,
  input  [29:0] auto_mem_in_ar_bits_addr,
  input  [2:0]  auto_mem_in_ar_bits_size,
  input         auto_mem_in_r_ready,
  output        auto_mem_in_r_valid,
  output        auto_mem_in_r_bits_id,
  output [31:0] auto_mem_in_r_bits_data,
  output        auto_in_in_ready,
  input         auto_in_in_valid,
  input  [7:0]  auto_in_in_bits_data,
  input         auto_out_out_ready,
  output        auto_out_out_valid,
  output [7:0]  auto_out_out_bits_data,
  output        int_0,
  output        io_txd,
  input         io_rxd
);
  wire  converter_auto_in_0; // @[Nodes.scala 31:31]
  wire  converter_auto_out_0; // @[Nodes.scala 31:31]
  wire  txm_clock; // @[DSPBlockUART.scala 101:21]
  wire  txm_reset; // @[DSPBlockUART.scala 101:21]
  wire  txm_io_en; // @[DSPBlockUART.scala 101:21]
  wire  txm_io_in_ready; // @[DSPBlockUART.scala 101:21]
  wire  txm_io_in_valid; // @[DSPBlockUART.scala 101:21]
  wire [7:0] txm_io_in_bits; // @[DSPBlockUART.scala 101:21]
  wire  txm_io_out; // @[DSPBlockUART.scala 101:21]
  wire [15:0] txm_io_div; // @[DSPBlockUART.scala 101:21]
  wire  txm_io_nstop; // @[DSPBlockUART.scala 101:21]
  wire  txq_clock; // @[DSPBlockUART.scala 102:21]
  wire  txq_reset; // @[DSPBlockUART.scala 102:21]
  wire  txq_io_enq_ready; // @[DSPBlockUART.scala 102:21]
  wire  txq_io_enq_valid; // @[DSPBlockUART.scala 102:21]
  wire [7:0] txq_io_enq_bits; // @[DSPBlockUART.scala 102:21]
  wire  txq_io_deq_ready; // @[DSPBlockUART.scala 102:21]
  wire  txq_io_deq_valid; // @[DSPBlockUART.scala 102:21]
  wire [7:0] txq_io_deq_bits; // @[DSPBlockUART.scala 102:21]
  wire [8:0] txq_io_count; // @[DSPBlockUART.scala 102:21]
  wire  rxm_clock; // @[DSPBlockUART.scala 104:21]
  wire  rxm_reset; // @[DSPBlockUART.scala 104:21]
  wire  rxm_io_en; // @[DSPBlockUART.scala 104:21]
  wire  rxm_io_in; // @[DSPBlockUART.scala 104:21]
  wire  rxm_io_out_valid; // @[DSPBlockUART.scala 104:21]
  wire [7:0] rxm_io_out_bits; // @[DSPBlockUART.scala 104:21]
  wire [15:0] rxm_io_div; // @[DSPBlockUART.scala 104:21]
  wire  rxq_clock; // @[DSPBlockUART.scala 105:21]
  wire  rxq_reset; // @[DSPBlockUART.scala 105:21]
  wire  rxq_io_enq_ready; // @[DSPBlockUART.scala 105:21]
  wire  rxq_io_enq_valid; // @[DSPBlockUART.scala 105:21]
  wire [7:0] rxq_io_enq_bits; // @[DSPBlockUART.scala 105:21]
  wire  rxq_io_deq_ready; // @[DSPBlockUART.scala 105:21]
  wire  rxq_io_deq_valid; // @[DSPBlockUART.scala 105:21]
  wire [7:0] rxq_io_deq_bits; // @[DSPBlockUART.scala 105:21]
  wire [8:0] rxq_io_count; // @[DSPBlockUART.scala 105:21]
  wire  Queue_clock; // @[Decoupled.scala 287:21]
  wire  Queue_reset; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_read; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_enq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_extra; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_read; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_deq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_extra; // @[Decoupled.scala 287:21]
  reg [15:0] div; // @[DSPBlockUART.scala 107:18]
  reg [31:0] _RAND_0;
  reg  txen; // @[DSPBlockUART.scala 113:19]
  reg [31:0] _RAND_1;
  reg  rxen; // @[DSPBlockUART.scala 114:19]
  reg [31:0] _RAND_2;
  reg [8:0] txwm; // @[DSPBlockUART.scala 121:19]
  reg [31:0] _RAND_3;
  reg [8:0] rxwm; // @[DSPBlockUART.scala 122:19]
  reg [31:0] _RAND_4;
  reg  nstop; // @[DSPBlockUART.scala 123:20]
  reg [31:0] _RAND_5;
  reg  ie_rxwm; // @[DSPBlockUART.scala 166:17]
  reg [31:0] _RAND_6;
  reg  ie_txwm; // @[DSPBlockUART.scala 166:17]
  reg [31:0] _RAND_7;
  wire  ip_txwm; // @[DSPBlockUART.scala 169:30]
  wire  ip_rxwm; // @[DSPBlockUART.scala 170:30]
  wire  _T_8; // @[DSPBlockUART.scala 171:31]
  wire  _T_9; // @[DSPBlockUART.scala 171:55]
  reg [31:0] _T_11; // @[DSPBlockUART.scala 175:53]
  reg [31:0] _RAND_8;
  reg [31:0] _T_12; // @[DSPBlockUART.scala 177:53]
  reg [31:0] _RAND_9;
  wire  _T_14; // @[RegisterRouter.scala 40:39]
  wire  _T_15; // @[RegisterRouter.scala 40:26]
  wire  _T_16; // @[RegisterRouter.scala 42:29]
  wire  _T_59_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 290:17]
  wire [29:0] _T_23; // @[RegisterRouter.scala 48:19]
  wire [2:0] _T_413; // @[Cat.scala 29:58]
  wire [5:0] _T_63; // @[RegisterRouter.scala 59:16]
  wire  _T_71; // @[RegisterRouter.scala 59:16]
  wire  _T_17; // @[RegisterRouter.scala 42:26]
  wire [1:0] _T_26; // @[OneHot.scala 65:12]
  wire [1:0] _T_28; // @[Misc.scala 200:81]
  wire  _T_29; // @[Misc.scala 204:21]
  wire  _T_32; // @[Misc.scala 209:20]
  wire  _T_34; // @[Misc.scala 213:38]
  wire  _T_35; // @[Misc.scala 213:29]
  wire  _T_37; // @[Misc.scala 213:38]
  wire  _T_38; // @[Misc.scala 213:29]
  wire  _T_41; // @[Misc.scala 209:20]
  wire  _T_42; // @[Misc.scala 212:27]
  wire  _T_43; // @[Misc.scala 213:38]
  wire  _T_44; // @[Misc.scala 213:29]
  wire  _T_45; // @[Misc.scala 212:27]
  wire  _T_46; // @[Misc.scala 213:38]
  wire  _T_47; // @[Misc.scala 213:29]
  wire  _T_48; // @[Misc.scala 212:27]
  wire  _T_49; // @[Misc.scala 213:38]
  wire  _T_50; // @[Misc.scala 213:29]
  wire  _T_51; // @[Misc.scala 212:27]
  wire  _T_52; // @[Misc.scala 213:38]
  wire  _T_53; // @[Misc.scala 213:29]
  wire [3:0] _T_56; // @[Cat.scala 29:58]
  wire [3:0] _T_58; // @[RegisterRouter.scala 54:25]
  wire [7:0] _T_87; // @[Bitwise.scala 72:12]
  wire [7:0] _T_89; // @[Bitwise.scala 72:12]
  wire [7:0] _T_91; // @[Bitwise.scala 72:12]
  wire [7:0] _T_93; // @[Bitwise.scala 72:12]
  wire [31:0] _T_96; // @[Cat.scala 29:58]
  wire  _T_115; // @[RegisterRouter.scala 59:16]
  wire  _T_432; // @[RegisterRouter.scala 59:16]
  wire [7:0] _T_414; // @[OneHot.scala 58:35]
  wire  _T_479; // @[RegisterRouter.scala 59:16]
  wire  _T_481; // @[RegisterRouter.scala 59:16]
  wire  _T_482; // @[RegisterRouter.scala 59:16]
  wire  _T_122; // @[RegisterRouter.scala 59:16]
  wire [1:0] _T_180; // @[Cat.scala 29:58]
  wire  _T_486; // @[RegisterRouter.scala 59:16]
  wire  _T_487; // @[RegisterRouter.scala 59:16]
  wire  _T_193; // @[RegisterRouter.scala 59:16]
  wire  _T_209; // @[RegisterRouter.scala 59:16]
  wire  _T_511; // @[RegisterRouter.scala 59:16]
  wire  _T_512; // @[RegisterRouter.scala 59:16]
  wire  _T_216; // @[RegisterRouter.scala 59:16]
  wire  _T_491; // @[RegisterRouter.scala 59:16]
  wire  _T_492; // @[RegisterRouter.scala 59:16]
  wire  _T_239; // @[RegisterRouter.scala 59:16]
  wire  _T_262; // @[RegisterRouter.scala 59:16]
  wire [1:0] _T_274; // @[Cat.scala 29:58]
  wire  _T_280; // @[RegisterRouter.scala 59:16]
  wire  _T_287; // @[RegisterRouter.scala 59:16]
  wire [15:0] _T_298; // @[RegisterRouter.scala 59:16]
  wire [24:0] _T_299; // @[Cat.scala 29:58]
  wire  _T_496; // @[RegisterRouter.scala 59:16]
  wire  _T_497; // @[RegisterRouter.scala 59:16]
  wire  _T_312; // @[RegisterRouter.scala 59:16]
  wire  _T_335; // @[RegisterRouter.scala 59:16]
  wire [15:0] _T_346; // @[RegisterRouter.scala 59:16]
  wire [24:0] _T_347; // @[Cat.scala 29:58]
  wire  _T_501; // @[RegisterRouter.scala 59:16]
  wire  _T_502; // @[RegisterRouter.scala 59:16]
  wire  _T_360; // @[RegisterRouter.scala 59:16]
  wire  _T_383; // @[RegisterRouter.scala 59:16]
  wire [1:0] _T_395; // @[Cat.scala 29:58]
  wire  _GEN_43; // @[MuxLiteral.scala 48:10]
  wire  _GEN_44; // @[MuxLiteral.scala 48:10]
  wire  _GEN_45; // @[MuxLiteral.scala 48:10]
  wire  _GEN_46; // @[MuxLiteral.scala 48:10]
  wire  _GEN_47; // @[MuxLiteral.scala 48:10]
  wire  _GEN_48; // @[MuxLiteral.scala 48:10]
  wire  _GEN_58; // @[MuxLiteral.scala 48:10]
  wire  _GEN_49; // @[MuxLiteral.scala 48:10]
  wire [31:0] _GEN_51; // @[MuxLiteral.scala 48:10]
  wire [31:0] _T_624_2; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [31:0] _GEN_52; // @[MuxLiteral.scala 48:10]
  wire [31:0] _T_624_3; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [31:0] _GEN_53; // @[MuxLiteral.scala 48:10]
  wire [31:0] _T_624_4; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [31:0] _GEN_54; // @[MuxLiteral.scala 48:10]
  wire [31:0] _T_624_5; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [31:0] _GEN_55; // @[MuxLiteral.scala 48:10]
  wire [31:0] _T_624_6; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [31:0] _GEN_56; // @[MuxLiteral.scala 48:10]
  wire [31:0] _GEN_57; // @[MuxLiteral.scala 48:10]
  wire  _T_627_bits_read; // @[Decoupled.scala 308:19 Decoupled.scala 309:14]
  wire  _T_627_valid; // @[Decoupled.scala 308:19 Decoupled.scala 310:15]
  wire  _T_630; // @[RegisterRouter.scala 65:29]
  IntToBundleBridge converter ( // @[Nodes.scala 31:31]
    .auto_in_0(converter_auto_in_0),
    .auto_out_0(converter_auto_out_0)
  );
  UARTTx txm ( // @[DSPBlockUART.scala 101:21]
    .clock(txm_clock),
    .reset(txm_reset),
    .io_en(txm_io_en),
    .io_in_ready(txm_io_in_ready),
    .io_in_valid(txm_io_in_valid),
    .io_in_bits(txm_io_in_bits),
    .io_out(txm_io_out),
    .io_div(txm_io_div),
    .io_nstop(txm_io_nstop)
  );
  QueueCompatibility_6 txq ( // @[DSPBlockUART.scala 102:21]
    .clock(txq_clock),
    .reset(txq_reset),
    .io_enq_ready(txq_io_enq_ready),
    .io_enq_valid(txq_io_enq_valid),
    .io_enq_bits(txq_io_enq_bits),
    .io_deq_ready(txq_io_deq_ready),
    .io_deq_valid(txq_io_deq_valid),
    .io_deq_bits(txq_io_deq_bits),
    .io_count(txq_io_count)
  );
  UARTRx rxm ( // @[DSPBlockUART.scala 104:21]
    .clock(rxm_clock),
    .reset(rxm_reset),
    .io_en(rxm_io_en),
    .io_in(rxm_io_in),
    .io_out_valid(rxm_io_out_valid),
    .io_out_bits(rxm_io_out_bits),
    .io_div(rxm_io_div)
  );
  QueueCompatibility_6 rxq ( // @[DSPBlockUART.scala 105:21]
    .clock(rxq_clock),
    .reset(rxq_reset),
    .io_enq_ready(rxq_io_enq_ready),
    .io_enq_valid(rxq_io_enq_valid),
    .io_enq_bits(rxq_io_enq_bits),
    .io_deq_ready(rxq_io_deq_ready),
    .io_deq_valid(rxq_io_deq_valid),
    .io_deq_bits(rxq_io_deq_bits),
    .io_count(rxq_io_count)
  );
  Queue Queue ( // @[Decoupled.scala 287:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_read(Queue_io_enq_bits_read),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_extra(Queue_io_enq_bits_extra),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_read(Queue_io_deq_bits_read),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_extra(Queue_io_deq_bits_extra)
  );
  assign ip_txwm = txq_io_count < txwm; // @[DSPBlockUART.scala 169:30]
  assign ip_rxwm = rxq_io_count > rxwm; // @[DSPBlockUART.scala 170:30]
  assign _T_8 = ip_txwm & ie_txwm; // @[DSPBlockUART.scala 171:31]
  assign _T_9 = ip_rxwm & ie_rxwm; // @[DSPBlockUART.scala 171:55]
  assign _T_14 = auto_mem_in_aw_valid & auto_mem_in_w_valid; // @[RegisterRouter.scala 40:39]
  assign _T_15 = auto_mem_in_ar_valid | _T_14; // @[RegisterRouter.scala 40:26]
  assign _T_16 = ~auto_mem_in_ar_valid; // @[RegisterRouter.scala 42:29]
  assign _T_59_ready = Queue_io_enq_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 290:17]
  assign _T_23 = auto_mem_in_ar_valid ? auto_mem_in_ar_bits_addr : auto_mem_in_aw_bits_addr; // @[RegisterRouter.scala 48:19]
  assign _T_413 = {_T_23[4],_T_23[3],_T_23[2]}; // @[Cat.scala 29:58]
  assign _T_63 = _T_23[7:2] & 6'h38; // @[RegisterRouter.scala 59:16]
  assign _T_71 = _T_63 == 6'h0; // @[RegisterRouter.scala 59:16]
  assign _T_17 = _T_59_ready & _T_16; // @[RegisterRouter.scala 42:26]
  assign _T_26 = 2'h1 << auto_mem_in_ar_bits_size[0]; // @[OneHot.scala 65:12]
  assign _T_28 = _T_26 | 2'h1; // @[Misc.scala 200:81]
  assign _T_29 = auto_mem_in_ar_bits_size >= 3'h2; // @[Misc.scala 204:21]
  assign _T_32 = ~auto_mem_in_ar_bits_addr[1]; // @[Misc.scala 209:20]
  assign _T_34 = _T_28[1] & _T_32; // @[Misc.scala 213:38]
  assign _T_35 = _T_29 | _T_34; // @[Misc.scala 213:29]
  assign _T_37 = _T_28[1] & auto_mem_in_ar_bits_addr[1]; // @[Misc.scala 213:38]
  assign _T_38 = _T_29 | _T_37; // @[Misc.scala 213:29]
  assign _T_41 = ~auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 209:20]
  assign _T_42 = _T_32 & _T_41; // @[Misc.scala 212:27]
  assign _T_43 = _T_28[0] & _T_42; // @[Misc.scala 213:38]
  assign _T_44 = _T_35 | _T_43; // @[Misc.scala 213:29]
  assign _T_45 = _T_32 & auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  assign _T_46 = _T_28[0] & _T_45; // @[Misc.scala 213:38]
  assign _T_47 = _T_35 | _T_46; // @[Misc.scala 213:29]
  assign _T_48 = auto_mem_in_ar_bits_addr[1] & _T_41; // @[Misc.scala 212:27]
  assign _T_49 = _T_28[0] & _T_48; // @[Misc.scala 213:38]
  assign _T_50 = _T_38 | _T_49; // @[Misc.scala 213:29]
  assign _T_51 = auto_mem_in_ar_bits_addr[1] & auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  assign _T_52 = _T_28[0] & _T_51; // @[Misc.scala 213:38]
  assign _T_53 = _T_38 | _T_52; // @[Misc.scala 213:29]
  assign _T_56 = {_T_53,_T_50,_T_47,_T_44}; // @[Cat.scala 29:58]
  assign _T_58 = auto_mem_in_ar_valid ? _T_56 : auto_mem_in_w_bits_strb; // @[RegisterRouter.scala 54:25]
  assign _T_87 = _T_58[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_89 = _T_58[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_91 = _T_58[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_93 = _T_58[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_96 = {_T_93,_T_91,_T_89,_T_87}; // @[Cat.scala 29:58]
  assign _T_115 = _T_96 == 32'hffffffff; // @[RegisterRouter.scala 59:16]
  assign _T_432 = _T_15 & _T_59_ready; // @[RegisterRouter.scala 59:16]
  assign _T_414 = 8'h1 << _T_413; // @[OneHot.scala 58:35]
  assign _T_479 = _T_432 & _T_16; // @[RegisterRouter.scala 59:16]
  assign _T_481 = _T_479 & _T_414[0]; // @[RegisterRouter.scala 59:16]
  assign _T_482 = _T_481 & _T_71; // @[RegisterRouter.scala 59:16]
  assign _T_122 = _T_482 & _T_115; // @[RegisterRouter.scala 59:16]
  assign _T_180 = {ip_rxwm,ip_txwm}; // @[Cat.scala 29:58]
  assign _T_486 = _T_479 & _T_414[1]; // @[RegisterRouter.scala 59:16]
  assign _T_487 = _T_486 & _T_71; // @[RegisterRouter.scala 59:16]
  assign _T_193 = _T_487 & _T_115; // @[RegisterRouter.scala 59:16]
  assign _T_209 = _T_96[15:0] == 16'hffff; // @[RegisterRouter.scala 59:16]
  assign _T_511 = _T_479 & _T_414[6]; // @[RegisterRouter.scala 59:16]
  assign _T_512 = _T_511 & _T_71; // @[RegisterRouter.scala 59:16]
  assign _T_216 = _T_512 & _T_209; // @[RegisterRouter.scala 59:16]
  assign _T_491 = _T_479 & _T_414[2]; // @[RegisterRouter.scala 59:16]
  assign _T_492 = _T_491 & _T_71; // @[RegisterRouter.scala 59:16]
  assign _T_239 = _T_492 & _T_96[0]; // @[RegisterRouter.scala 59:16]
  assign _T_262 = _T_492 & _T_96[1]; // @[RegisterRouter.scala 59:16]
  assign _T_274 = {nstop,txen}; // @[Cat.scala 29:58]
  assign _T_280 = _T_96[24:16] == 9'h1ff; // @[RegisterRouter.scala 59:16]
  assign _T_287 = _T_492 & _T_280; // @[RegisterRouter.scala 59:16]
  assign _T_298 = {{14'd0}, _T_274}; // @[RegisterRouter.scala 59:16]
  assign _T_299 = {txwm,_T_298}; // @[Cat.scala 29:58]
  assign _T_496 = _T_479 & _T_414[3]; // @[RegisterRouter.scala 59:16]
  assign _T_497 = _T_496 & _T_71; // @[RegisterRouter.scala 59:16]
  assign _T_312 = _T_497 & _T_96[0]; // @[RegisterRouter.scala 59:16]
  assign _T_335 = _T_497 & _T_280; // @[RegisterRouter.scala 59:16]
  assign _T_346 = {{15'd0}, rxen}; // @[RegisterRouter.scala 59:16]
  assign _T_347 = {rxwm,_T_346}; // @[Cat.scala 29:58]
  assign _T_501 = _T_479 & _T_414[4]; // @[RegisterRouter.scala 59:16]
  assign _T_502 = _T_501 & _T_71; // @[RegisterRouter.scala 59:16]
  assign _T_360 = _T_502 & _T_96[0]; // @[RegisterRouter.scala 59:16]
  assign _T_383 = _T_502 & _T_96[1]; // @[RegisterRouter.scala 59:16]
  assign _T_395 = {ie_rxwm,ie_txwm}; // @[Cat.scala 29:58]
  assign _GEN_43 = 3'h1 == _T_413 ? _T_71 : _T_71; // @[MuxLiteral.scala 48:10]
  assign _GEN_44 = 3'h2 == _T_413 ? _T_71 : _GEN_43; // @[MuxLiteral.scala 48:10]
  assign _GEN_45 = 3'h3 == _T_413 ? _T_71 : _GEN_44; // @[MuxLiteral.scala 48:10]
  assign _GEN_46 = 3'h4 == _T_413 ? _T_71 : _GEN_45; // @[MuxLiteral.scala 48:10]
  assign _GEN_47 = 3'h5 == _T_413 ? _T_71 : _GEN_46; // @[MuxLiteral.scala 48:10]
  assign _GEN_48 = 3'h6 == _T_413 ? _T_71 : _GEN_47; // @[MuxLiteral.scala 48:10]
  assign _GEN_58 = 3'h7 == _T_413; // @[MuxLiteral.scala 48:10]
  assign _GEN_49 = _GEN_58 | _GEN_48; // @[MuxLiteral.scala 48:10]
  assign _GEN_51 = 3'h1 == _T_413 ? _T_12 : _T_11; // @[MuxLiteral.scala 48:10]
  assign _T_624_2 = {{7'd0}, _T_299}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  assign _GEN_52 = 3'h2 == _T_413 ? _T_624_2 : _GEN_51; // @[MuxLiteral.scala 48:10]
  assign _T_624_3 = {{7'd0}, _T_347}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  assign _GEN_53 = 3'h3 == _T_413 ? _T_624_3 : _GEN_52; // @[MuxLiteral.scala 48:10]
  assign _T_624_4 = {{30'd0}, _T_395}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  assign _GEN_54 = 3'h4 == _T_413 ? _T_624_4 : _GEN_53; // @[MuxLiteral.scala 48:10]
  assign _T_624_5 = {{30'd0}, _T_180}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  assign _GEN_55 = 3'h5 == _T_413 ? _T_624_5 : _GEN_54; // @[MuxLiteral.scala 48:10]
  assign _T_624_6 = {{16'd0}, div}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  assign _GEN_56 = 3'h6 == _T_413 ? _T_624_6 : _GEN_55; // @[MuxLiteral.scala 48:10]
  assign _GEN_57 = 3'h7 == _T_413 ? 32'h0 : _GEN_56; // @[MuxLiteral.scala 48:10]
  assign _T_627_bits_read = Queue_io_deq_bits_read; // @[Decoupled.scala 308:19 Decoupled.scala 309:14]
  assign _T_627_valid = Queue_io_deq_valid; // @[Decoupled.scala 308:19 Decoupled.scala 310:15]
  assign _T_630 = ~_T_627_bits_read; // @[RegisterRouter.scala 65:29]
  assign auto_mem_in_aw_ready = _T_17 & auto_mem_in_w_valid; // @[LazyModule.scala 173:31]
  assign auto_mem_in_w_ready = _T_17 & auto_mem_in_aw_valid; // @[LazyModule.scala 173:31]
  assign auto_mem_in_b_valid = _T_627_valid & _T_630; // @[LazyModule.scala 173:31]
  assign auto_mem_in_b_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_mem_in_ar_ready = Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_valid = _T_627_valid & _T_627_bits_read; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 173:31]
  assign auto_in_in_ready = txq_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_out_out_valid = rxq_io_deq_valid; // @[LazyModule.scala 173:49]
  assign auto_out_out_bits_data = rxq_io_deq_bits; // @[LazyModule.scala 173:49]
  assign int_0 = converter_auto_out_0; // @[SpectrometerTestWithoutLA.scala 119:12]
  assign io_txd = txm_io_out; // @[DSPBlockUART.scala 135:12]
  assign converter_auto_in_0 = _T_8 | _T_9; // @[LazyModule.scala 167:57]
  assign txm_clock = clock;
  assign txm_reset = reset;
  assign txm_io_en = txen; // @[DSPBlockUART.scala 131:19]
  assign txm_io_in_valid = txq_io_deq_valid; // @[DSPBlockUART.scala 132:15]
  assign txm_io_in_bits = txq_io_deq_bits; // @[DSPBlockUART.scala 132:15]
  assign txm_io_div = div; // @[DSPBlockUART.scala 133:16]
  assign txm_io_nstop = nstop; // @[DSPBlockUART.scala 134:18]
  assign txq_clock = clock;
  assign txq_reset = reset;
  assign txq_io_enq_valid = auto_in_in_valid; // @[DSPBlockUART.scala 139:22]
  assign txq_io_enq_bits = auto_in_in_bits_data; // @[DSPBlockUART.scala 138:22]
  assign txq_io_deq_ready = txm_io_in_ready; // @[DSPBlockUART.scala 132:15]
  assign rxm_clock = clock;
  assign rxm_reset = reset;
  assign rxm_io_en = rxen; // @[DSPBlockUART.scala 151:15]
  assign rxm_io_in = io_rxd; // @[DSPBlockUART.scala 152:15]
  assign rxm_io_div = div; // @[DSPBlockUART.scala 154:16]
  assign rxq_clock = clock;
  assign rxq_reset = reset;
  assign rxq_io_enq_valid = rxm_io_out_valid; // @[DSPBlockUART.scala 153:16]
  assign rxq_io_enq_bits = rxm_io_out_bits; // @[DSPBlockUART.scala 153:16]
  assign rxq_io_deq_ready = auto_out_out_ready; // @[DSPBlockUART.scala 144:22]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_mem_in_ar_valid | _T_14; // @[Decoupled.scala 288:22]
  assign Queue_io_enq_bits_read = auto_mem_in_ar_valid; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_data = _GEN_49 ? _GEN_57 : 32'h0; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_extra = auto_mem_in_ar_valid ? auto_mem_in_ar_bits_id : auto_mem_in_aw_bits_id; // @[Decoupled.scala 289:21]
  assign Queue_io_deq_ready = _T_627_bits_read ? auto_mem_in_r_ready : auto_mem_in_b_ready; // @[Decoupled.scala 311:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  div = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  txen = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  rxen = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  txwm = _RAND_3[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  rxwm = _RAND_4[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  nstop = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  ie_rxwm = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  ie_txwm = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_11 = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_12 = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      div <= 16'h365;
    end else if (_T_216) begin
      div <= auto_mem_in_w_bits_data[15:0];
    end
    if (reset) begin
      txen <= 1'h0;
    end else if (_T_239) begin
      txen <= auto_mem_in_w_bits_data[0];
    end
    if (reset) begin
      rxen <= 1'h0;
    end else if (_T_312) begin
      rxen <= auto_mem_in_w_bits_data[0];
    end
    if (reset) begin
      txwm <= 9'h0;
    end else if (_T_287) begin
      txwm <= auto_mem_in_w_bits_data[24:16];
    end
    if (reset) begin
      rxwm <= 9'h0;
    end else if (_T_335) begin
      rxwm <= auto_mem_in_w_bits_data[24:16];
    end
    if (reset) begin
      nstop <= 1'h0;
    end else if (_T_262) begin
      nstop <= auto_mem_in_w_bits_data[1];
    end
    if (reset) begin
      ie_rxwm <= 1'h0;
    end else if (_T_383) begin
      ie_rxwm <= auto_mem_in_w_bits_data[1];
    end
    if (reset) begin
      ie_txwm <= 1'h0;
    end else if (_T_360) begin
      ie_txwm <= auto_mem_in_w_bits_data[0];
    end
    if (reset) begin
      _T_11 <= 32'h0;
    end else if (_T_122) begin
      _T_11 <= auto_mem_in_w_bits_data;
    end
    if (reset) begin
      _T_12 <= 32'h0;
    end else if (_T_193) begin
      _T_12 <= auto_mem_in_w_bits_data;
    end
  end
endmodule
module QueueCompatibility_8(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [21:0] io_enq_bits,
  input         io_deq_ready,
  output        io_deq_valid,
  output [21:0] io_deq_bits
);
  reg [21:0] _T [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_0;
  wire [21:0] _T__T_18_data; // @[Decoupled.scala 209:24]
  wire  _T__T_18_addr; // @[Decoupled.scala 209:24]
  wire [21:0] _T__T_10_data; // @[Decoupled.scala 209:24]
  wire  _T__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T__T_10_en; // @[Decoupled.scala 209:24]
  reg  value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_1;
  reg  value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_2;
  reg  _T_1; // @[Decoupled.scala 212:35]
  reg [31:0] _RAND_3;
  wire  _T_2; // @[Decoupled.scala 214:41]
  wire  _T_3; // @[Decoupled.scala 215:36]
  wire  _T_4; // @[Decoupled.scala 215:33]
  wire  _T_5; // @[Decoupled.scala 216:32]
  wire  _T_6; // @[Decoupled.scala 40:37]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _T_12; // @[Counter.scala 39:22]
  wire  _GEN_9; // @[Decoupled.scala 240:27]
  wire  _GEN_12; // @[Decoupled.scala 237:18]
  wire  _T_14; // @[Counter.scala 39:22]
  wire  _GEN_11; // @[Decoupled.scala 237:18]
  wire  _T_15; // @[Decoupled.scala 227:16]
  wire  _T_16; // @[Decoupled.scala 231:19]
  assign _T__T_18_addr = value_1;
  assign _T__T_18_data = _T[_T__T_18_addr]; // @[Decoupled.scala 209:24]
  assign _T__T_10_data = io_enq_bits;
  assign _T__T_10_addr = value;
  assign _T__T_10_mask = 1'h1;
  assign _T__T_10_en = _T_4 ? _GEN_9 : _T_6;
  assign _T_2 = value == value_1; // @[Decoupled.scala 214:41]
  assign _T_3 = ~_T_1; // @[Decoupled.scala 215:36]
  assign _T_4 = _T_2 & _T_3; // @[Decoupled.scala 215:33]
  assign _T_5 = _T_2 & _T_1; // @[Decoupled.scala 216:32]
  assign _T_6 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  assign _T_8 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  assign _T_12 = value + 1'h1; // @[Counter.scala 39:22]
  assign _GEN_9 = io_deq_ready ? 1'h0 : _T_6; // @[Decoupled.scala 240:27]
  assign _GEN_12 = _T_4 ? _GEN_9 : _T_6; // @[Decoupled.scala 237:18]
  assign _T_14 = value_1 + 1'h1; // @[Counter.scala 39:22]
  assign _GEN_11 = _T_4 ? 1'h0 : _T_8; // @[Decoupled.scala 237:18]
  assign _T_15 = _GEN_12 != _GEN_11; // @[Decoupled.scala 227:16]
  assign _T_16 = ~_T_4; // @[Decoupled.scala 231:19]
  assign io_enq_ready = ~_T_5; // @[Decoupled.scala 232:16]
  assign io_deq_valid = io_enq_valid | _T_16; // @[Decoupled.scala 231:16 Decoupled.scala 236:40]
  assign io_deq_bits = _T_4 ? io_enq_bits : _T__T_18_data; // @[Decoupled.scala 233:15 Decoupled.scala 238:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T[initvar] = _RAND_0[21:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  value = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  value_1 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_1 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T__T_10_en & _T__T_10_mask) begin
      _T[_T__T_10_addr] <= _T__T_10_data; // @[Decoupled.scala 209:24]
    end
    if (reset) begin
      value <= 1'h0;
    end else if (_GEN_12) begin
      value <= _T_12;
    end
    if (reset) begin
      value_1 <= 1'h0;
    end else if (_GEN_11) begin
      value_1 <= _T_14;
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else if (_T_15) begin
      if (_T_4) begin
        if (io_deq_ready) begin
          _T_1 <= 1'h0;
        end else begin
          _T_1 <= _T_6;
        end
      end else begin
        _T_1 <= _T_6;
      end
    end
  end
endmodule
module AXI4Xbar_2(
  input         clock,
  input         reset,
  output        auto_in_aw_ready,
  input         auto_in_aw_valid,
  input         auto_in_aw_bits_id,
  input  [29:0] auto_in_aw_bits_addr,
  input  [2:0]  auto_in_aw_bits_size,
  output        auto_in_w_ready,
  input         auto_in_w_valid,
  input  [31:0] auto_in_w_bits_data,
  input  [3:0]  auto_in_w_bits_strb,
  input         auto_in_w_bits_last,
  input         auto_in_b_ready,
  output        auto_in_b_valid,
  output [1:0]  auto_in_b_bits_resp,
  output        auto_in_ar_ready,
  input         auto_in_ar_valid,
  input         auto_in_ar_bits_id,
  input  [29:0] auto_in_ar_bits_addr,
  input  [2:0]  auto_in_ar_bits_size,
  input         auto_in_r_ready,
  output        auto_in_r_valid,
  output [31:0] auto_in_r_bits_data,
  output [1:0]  auto_in_r_bits_resp,
  output        auto_in_r_bits_last,
  input         auto_out_21_aw_ready,
  output        auto_out_21_aw_valid,
  output        auto_out_21_aw_bits_id,
  output [29:0] auto_out_21_aw_bits_addr,
  output [2:0]  auto_out_21_aw_bits_size,
  input         auto_out_21_w_ready,
  output        auto_out_21_w_valid,
  output [31:0] auto_out_21_w_bits_data,
  output [3:0]  auto_out_21_w_bits_strb,
  output        auto_out_21_w_bits_last,
  output        auto_out_21_b_ready,
  input         auto_out_21_b_valid,
  input  [1:0]  auto_out_21_b_bits_resp,
  input         auto_out_21_ar_ready,
  output        auto_out_21_ar_valid,
  output        auto_out_21_ar_bits_id,
  output [29:0] auto_out_21_ar_bits_addr,
  output [2:0]  auto_out_21_ar_bits_size,
  output        auto_out_21_r_ready,
  input         auto_out_21_r_valid,
  input  [31:0] auto_out_21_r_bits_data,
  input  [1:0]  auto_out_21_r_bits_resp,
  input         auto_out_21_r_bits_last,
  input         auto_out_20_aw_ready,
  output        auto_out_20_aw_valid,
  output        auto_out_20_aw_bits_id,
  output [29:0] auto_out_20_aw_bits_addr,
  output [2:0]  auto_out_20_aw_bits_size,
  input         auto_out_20_w_ready,
  output        auto_out_20_w_valid,
  output [31:0] auto_out_20_w_bits_data,
  output [3:0]  auto_out_20_w_bits_strb,
  output        auto_out_20_w_bits_last,
  output        auto_out_20_b_ready,
  input         auto_out_20_b_valid,
  input         auto_out_20_b_bits_id,
  input  [1:0]  auto_out_20_b_bits_resp,
  input         auto_out_20_ar_ready,
  output        auto_out_20_ar_valid,
  output        auto_out_20_ar_bits_id,
  output [29:0] auto_out_20_ar_bits_addr,
  output [2:0]  auto_out_20_ar_bits_size,
  output        auto_out_20_r_ready,
  input         auto_out_20_r_valid,
  input         auto_out_20_r_bits_id,
  input  [31:0] auto_out_20_r_bits_data,
  input  [1:0]  auto_out_20_r_bits_resp,
  input         auto_out_20_r_bits_last,
  input         auto_out_19_aw_ready,
  output        auto_out_19_aw_valid,
  output        auto_out_19_aw_bits_id,
  output [29:0] auto_out_19_aw_bits_addr,
  output [2:0]  auto_out_19_aw_bits_size,
  input         auto_out_19_w_ready,
  output        auto_out_19_w_valid,
  output [31:0] auto_out_19_w_bits_data,
  output [3:0]  auto_out_19_w_bits_strb,
  output        auto_out_19_w_bits_last,
  output        auto_out_19_b_ready,
  input         auto_out_19_b_valid,
  input         auto_out_19_b_bits_id,
  input  [1:0]  auto_out_19_b_bits_resp,
  input         auto_out_19_ar_ready,
  output        auto_out_19_ar_valid,
  output        auto_out_19_ar_bits_id,
  output [29:0] auto_out_19_ar_bits_addr,
  output [2:0]  auto_out_19_ar_bits_size,
  output        auto_out_19_r_ready,
  input         auto_out_19_r_valid,
  input         auto_out_19_r_bits_id,
  input  [31:0] auto_out_19_r_bits_data,
  input  [1:0]  auto_out_19_r_bits_resp,
  input         auto_out_19_r_bits_last,
  input         auto_out_18_aw_ready,
  output        auto_out_18_aw_valid,
  output        auto_out_18_aw_bits_id,
  output [29:0] auto_out_18_aw_bits_addr,
  output [2:0]  auto_out_18_aw_bits_size,
  input         auto_out_18_w_ready,
  output        auto_out_18_w_valid,
  output [31:0] auto_out_18_w_bits_data,
  output [3:0]  auto_out_18_w_bits_strb,
  output        auto_out_18_w_bits_last,
  output        auto_out_18_b_ready,
  input         auto_out_18_b_valid,
  input         auto_out_18_b_bits_id,
  input  [1:0]  auto_out_18_b_bits_resp,
  input         auto_out_18_ar_ready,
  output        auto_out_18_ar_valid,
  output        auto_out_18_ar_bits_id,
  output [29:0] auto_out_18_ar_bits_addr,
  output [2:0]  auto_out_18_ar_bits_size,
  output        auto_out_18_r_ready,
  input         auto_out_18_r_valid,
  input         auto_out_18_r_bits_id,
  input  [31:0] auto_out_18_r_bits_data,
  input  [1:0]  auto_out_18_r_bits_resp,
  input         auto_out_18_r_bits_last,
  input         auto_out_17_aw_ready,
  output        auto_out_17_aw_valid,
  output        auto_out_17_aw_bits_id,
  output [29:0] auto_out_17_aw_bits_addr,
  output [2:0]  auto_out_17_aw_bits_size,
  input         auto_out_17_w_ready,
  output        auto_out_17_w_valid,
  output [31:0] auto_out_17_w_bits_data,
  output [3:0]  auto_out_17_w_bits_strb,
  output        auto_out_17_w_bits_last,
  output        auto_out_17_b_ready,
  input         auto_out_17_b_valid,
  input         auto_out_17_b_bits_id,
  input  [1:0]  auto_out_17_b_bits_resp,
  input         auto_out_17_ar_ready,
  output        auto_out_17_ar_valid,
  output        auto_out_17_ar_bits_id,
  output [29:0] auto_out_17_ar_bits_addr,
  output [2:0]  auto_out_17_ar_bits_size,
  output        auto_out_17_r_ready,
  input         auto_out_17_r_valid,
  input         auto_out_17_r_bits_id,
  input  [31:0] auto_out_17_r_bits_data,
  input  [1:0]  auto_out_17_r_bits_resp,
  input         auto_out_17_r_bits_last,
  input         auto_out_16_aw_ready,
  output        auto_out_16_aw_valid,
  output        auto_out_16_aw_bits_id,
  output [29:0] auto_out_16_aw_bits_addr,
  output [2:0]  auto_out_16_aw_bits_size,
  input         auto_out_16_w_ready,
  output        auto_out_16_w_valid,
  output [31:0] auto_out_16_w_bits_data,
  output [3:0]  auto_out_16_w_bits_strb,
  output        auto_out_16_w_bits_last,
  output        auto_out_16_b_ready,
  input         auto_out_16_b_valid,
  input         auto_out_16_b_bits_id,
  input  [1:0]  auto_out_16_b_bits_resp,
  input         auto_out_16_ar_ready,
  output        auto_out_16_ar_valid,
  output        auto_out_16_ar_bits_id,
  output [29:0] auto_out_16_ar_bits_addr,
  output [2:0]  auto_out_16_ar_bits_size,
  output        auto_out_16_r_ready,
  input         auto_out_16_r_valid,
  input         auto_out_16_r_bits_id,
  input  [31:0] auto_out_16_r_bits_data,
  input  [1:0]  auto_out_16_r_bits_resp,
  input         auto_out_16_r_bits_last,
  input         auto_out_15_aw_ready,
  output        auto_out_15_aw_valid,
  output        auto_out_15_aw_bits_id,
  output [29:0] auto_out_15_aw_bits_addr,
  output [2:0]  auto_out_15_aw_bits_size,
  input         auto_out_15_w_ready,
  output        auto_out_15_w_valid,
  output [31:0] auto_out_15_w_bits_data,
  output [3:0]  auto_out_15_w_bits_strb,
  output        auto_out_15_w_bits_last,
  output        auto_out_15_b_ready,
  input         auto_out_15_b_valid,
  input         auto_out_15_b_bits_id,
  input  [1:0]  auto_out_15_b_bits_resp,
  input         auto_out_15_ar_ready,
  output        auto_out_15_ar_valid,
  output        auto_out_15_ar_bits_id,
  output [29:0] auto_out_15_ar_bits_addr,
  output [2:0]  auto_out_15_ar_bits_size,
  output        auto_out_15_r_ready,
  input         auto_out_15_r_valid,
  input         auto_out_15_r_bits_id,
  input  [31:0] auto_out_15_r_bits_data,
  input  [1:0]  auto_out_15_r_bits_resp,
  input         auto_out_15_r_bits_last,
  input         auto_out_14_aw_ready,
  output        auto_out_14_aw_valid,
  output        auto_out_14_aw_bits_id,
  output [29:0] auto_out_14_aw_bits_addr,
  output [2:0]  auto_out_14_aw_bits_size,
  input         auto_out_14_w_ready,
  output        auto_out_14_w_valid,
  output [31:0] auto_out_14_w_bits_data,
  output [3:0]  auto_out_14_w_bits_strb,
  output        auto_out_14_w_bits_last,
  output        auto_out_14_b_ready,
  input         auto_out_14_b_valid,
  input         auto_out_14_b_bits_id,
  input  [1:0]  auto_out_14_b_bits_resp,
  input         auto_out_14_ar_ready,
  output        auto_out_14_ar_valid,
  output        auto_out_14_ar_bits_id,
  output [29:0] auto_out_14_ar_bits_addr,
  output [2:0]  auto_out_14_ar_bits_size,
  output        auto_out_14_r_ready,
  input         auto_out_14_r_valid,
  input         auto_out_14_r_bits_id,
  input  [31:0] auto_out_14_r_bits_data,
  input  [1:0]  auto_out_14_r_bits_resp,
  input         auto_out_14_r_bits_last,
  input         auto_out_13_aw_ready,
  output        auto_out_13_aw_valid,
  output        auto_out_13_aw_bits_id,
  output [29:0] auto_out_13_aw_bits_addr,
  output [2:0]  auto_out_13_aw_bits_size,
  input         auto_out_13_w_ready,
  output        auto_out_13_w_valid,
  output [31:0] auto_out_13_w_bits_data,
  output [3:0]  auto_out_13_w_bits_strb,
  output        auto_out_13_w_bits_last,
  output        auto_out_13_b_ready,
  input         auto_out_13_b_valid,
  input         auto_out_13_b_bits_id,
  input  [1:0]  auto_out_13_b_bits_resp,
  input         auto_out_13_ar_ready,
  output        auto_out_13_ar_valid,
  output        auto_out_13_ar_bits_id,
  output [29:0] auto_out_13_ar_bits_addr,
  output [2:0]  auto_out_13_ar_bits_size,
  output        auto_out_13_r_ready,
  input         auto_out_13_r_valid,
  input         auto_out_13_r_bits_id,
  input  [31:0] auto_out_13_r_bits_data,
  input  [1:0]  auto_out_13_r_bits_resp,
  input         auto_out_13_r_bits_last,
  input         auto_out_12_aw_ready,
  output        auto_out_12_aw_valid,
  output        auto_out_12_aw_bits_id,
  output [29:0] auto_out_12_aw_bits_addr,
  output [2:0]  auto_out_12_aw_bits_size,
  input         auto_out_12_w_ready,
  output        auto_out_12_w_valid,
  output [31:0] auto_out_12_w_bits_data,
  output [3:0]  auto_out_12_w_bits_strb,
  output        auto_out_12_w_bits_last,
  output        auto_out_12_b_ready,
  input         auto_out_12_b_valid,
  input         auto_out_12_b_bits_id,
  input  [1:0]  auto_out_12_b_bits_resp,
  input         auto_out_12_ar_ready,
  output        auto_out_12_ar_valid,
  output        auto_out_12_ar_bits_id,
  output [29:0] auto_out_12_ar_bits_addr,
  output [2:0]  auto_out_12_ar_bits_size,
  output        auto_out_12_r_ready,
  input         auto_out_12_r_valid,
  input         auto_out_12_r_bits_id,
  input  [31:0] auto_out_12_r_bits_data,
  input  [1:0]  auto_out_12_r_bits_resp,
  input         auto_out_12_r_bits_last,
  input         auto_out_11_aw_ready,
  output        auto_out_11_aw_valid,
  output        auto_out_11_aw_bits_id,
  output [29:0] auto_out_11_aw_bits_addr,
  output [2:0]  auto_out_11_aw_bits_size,
  input         auto_out_11_w_ready,
  output        auto_out_11_w_valid,
  output [31:0] auto_out_11_w_bits_data,
  output [3:0]  auto_out_11_w_bits_strb,
  output        auto_out_11_w_bits_last,
  output        auto_out_11_b_ready,
  input         auto_out_11_b_valid,
  input         auto_out_11_b_bits_id,
  input  [1:0]  auto_out_11_b_bits_resp,
  input         auto_out_11_ar_ready,
  output        auto_out_11_ar_valid,
  output        auto_out_11_ar_bits_id,
  output [29:0] auto_out_11_ar_bits_addr,
  output [2:0]  auto_out_11_ar_bits_size,
  output        auto_out_11_r_ready,
  input         auto_out_11_r_valid,
  input         auto_out_11_r_bits_id,
  input  [31:0] auto_out_11_r_bits_data,
  input  [1:0]  auto_out_11_r_bits_resp,
  input         auto_out_11_r_bits_last,
  input         auto_out_10_aw_ready,
  output        auto_out_10_aw_valid,
  output        auto_out_10_aw_bits_id,
  output [29:0] auto_out_10_aw_bits_addr,
  output [2:0]  auto_out_10_aw_bits_size,
  input         auto_out_10_w_ready,
  output        auto_out_10_w_valid,
  output [31:0] auto_out_10_w_bits_data,
  output [3:0]  auto_out_10_w_bits_strb,
  output        auto_out_10_w_bits_last,
  output        auto_out_10_b_ready,
  input         auto_out_10_b_valid,
  input         auto_out_10_b_bits_id,
  input  [1:0]  auto_out_10_b_bits_resp,
  input         auto_out_10_ar_ready,
  output        auto_out_10_ar_valid,
  output        auto_out_10_ar_bits_id,
  output [29:0] auto_out_10_ar_bits_addr,
  output [2:0]  auto_out_10_ar_bits_size,
  output        auto_out_10_r_ready,
  input         auto_out_10_r_valid,
  input         auto_out_10_r_bits_id,
  input  [31:0] auto_out_10_r_bits_data,
  input  [1:0]  auto_out_10_r_bits_resp,
  input         auto_out_10_r_bits_last,
  input         auto_out_9_aw_ready,
  output        auto_out_9_aw_valid,
  output        auto_out_9_aw_bits_id,
  output [29:0] auto_out_9_aw_bits_addr,
  output [2:0]  auto_out_9_aw_bits_size,
  input         auto_out_9_w_ready,
  output        auto_out_9_w_valid,
  output [31:0] auto_out_9_w_bits_data,
  output [3:0]  auto_out_9_w_bits_strb,
  output        auto_out_9_w_bits_last,
  output        auto_out_9_b_ready,
  input         auto_out_9_b_valid,
  input         auto_out_9_b_bits_id,
  input  [1:0]  auto_out_9_b_bits_resp,
  input         auto_out_9_ar_ready,
  output        auto_out_9_ar_valid,
  output        auto_out_9_ar_bits_id,
  output [29:0] auto_out_9_ar_bits_addr,
  output [2:0]  auto_out_9_ar_bits_size,
  output        auto_out_9_r_ready,
  input         auto_out_9_r_valid,
  input         auto_out_9_r_bits_id,
  input  [31:0] auto_out_9_r_bits_data,
  input  [1:0]  auto_out_9_r_bits_resp,
  input         auto_out_9_r_bits_last,
  input         auto_out_8_aw_ready,
  output        auto_out_8_aw_valid,
  output        auto_out_8_aw_bits_id,
  output [29:0] auto_out_8_aw_bits_addr,
  output [2:0]  auto_out_8_aw_bits_size,
  input         auto_out_8_w_ready,
  output        auto_out_8_w_valid,
  output [31:0] auto_out_8_w_bits_data,
  output [3:0]  auto_out_8_w_bits_strb,
  output        auto_out_8_w_bits_last,
  output        auto_out_8_b_ready,
  input         auto_out_8_b_valid,
  input         auto_out_8_b_bits_id,
  input  [1:0]  auto_out_8_b_bits_resp,
  input         auto_out_8_ar_ready,
  output        auto_out_8_ar_valid,
  output        auto_out_8_ar_bits_id,
  output [29:0] auto_out_8_ar_bits_addr,
  output [2:0]  auto_out_8_ar_bits_size,
  output        auto_out_8_r_ready,
  input         auto_out_8_r_valid,
  input         auto_out_8_r_bits_id,
  input  [31:0] auto_out_8_r_bits_data,
  input  [1:0]  auto_out_8_r_bits_resp,
  input         auto_out_8_r_bits_last,
  input         auto_out_7_aw_ready,
  output        auto_out_7_aw_valid,
  output        auto_out_7_aw_bits_id,
  output [29:0] auto_out_7_aw_bits_addr,
  output [2:0]  auto_out_7_aw_bits_size,
  input         auto_out_7_w_ready,
  output        auto_out_7_w_valid,
  output [31:0] auto_out_7_w_bits_data,
  output [3:0]  auto_out_7_w_bits_strb,
  output        auto_out_7_w_bits_last,
  output        auto_out_7_b_ready,
  input         auto_out_7_b_valid,
  input         auto_out_7_b_bits_id,
  input  [1:0]  auto_out_7_b_bits_resp,
  input         auto_out_7_ar_ready,
  output        auto_out_7_ar_valid,
  output        auto_out_7_ar_bits_id,
  output [29:0] auto_out_7_ar_bits_addr,
  output [2:0]  auto_out_7_ar_bits_size,
  output        auto_out_7_r_ready,
  input         auto_out_7_r_valid,
  input         auto_out_7_r_bits_id,
  input  [31:0] auto_out_7_r_bits_data,
  input  [1:0]  auto_out_7_r_bits_resp,
  input         auto_out_7_r_bits_last,
  input         auto_out_6_aw_ready,
  output        auto_out_6_aw_valid,
  output        auto_out_6_aw_bits_id,
  output [29:0] auto_out_6_aw_bits_addr,
  output [2:0]  auto_out_6_aw_bits_size,
  input         auto_out_6_w_ready,
  output        auto_out_6_w_valid,
  output [31:0] auto_out_6_w_bits_data,
  output [3:0]  auto_out_6_w_bits_strb,
  output        auto_out_6_w_bits_last,
  output        auto_out_6_b_ready,
  input         auto_out_6_b_valid,
  input         auto_out_6_b_bits_id,
  input  [1:0]  auto_out_6_b_bits_resp,
  input         auto_out_6_ar_ready,
  output        auto_out_6_ar_valid,
  output        auto_out_6_ar_bits_id,
  output [29:0] auto_out_6_ar_bits_addr,
  output [2:0]  auto_out_6_ar_bits_size,
  output        auto_out_6_r_ready,
  input         auto_out_6_r_valid,
  input         auto_out_6_r_bits_id,
  input  [31:0] auto_out_6_r_bits_data,
  input  [1:0]  auto_out_6_r_bits_resp,
  input         auto_out_6_r_bits_last,
  input         auto_out_5_aw_ready,
  output        auto_out_5_aw_valid,
  output        auto_out_5_aw_bits_id,
  output [29:0] auto_out_5_aw_bits_addr,
  output [2:0]  auto_out_5_aw_bits_size,
  input         auto_out_5_w_ready,
  output        auto_out_5_w_valid,
  output [31:0] auto_out_5_w_bits_data,
  output [3:0]  auto_out_5_w_bits_strb,
  output        auto_out_5_w_bits_last,
  output        auto_out_5_b_ready,
  input         auto_out_5_b_valid,
  input         auto_out_5_b_bits_id,
  input  [1:0]  auto_out_5_b_bits_resp,
  input         auto_out_5_ar_ready,
  output        auto_out_5_ar_valid,
  output        auto_out_5_ar_bits_id,
  output [29:0] auto_out_5_ar_bits_addr,
  output [2:0]  auto_out_5_ar_bits_size,
  output        auto_out_5_r_ready,
  input         auto_out_5_r_valid,
  input         auto_out_5_r_bits_id,
  input  [31:0] auto_out_5_r_bits_data,
  input  [1:0]  auto_out_5_r_bits_resp,
  input         auto_out_5_r_bits_last,
  input         auto_out_4_aw_ready,
  output        auto_out_4_aw_valid,
  output        auto_out_4_aw_bits_id,
  output [29:0] auto_out_4_aw_bits_addr,
  output [2:0]  auto_out_4_aw_bits_size,
  input         auto_out_4_w_ready,
  output        auto_out_4_w_valid,
  output [31:0] auto_out_4_w_bits_data,
  output [3:0]  auto_out_4_w_bits_strb,
  output        auto_out_4_w_bits_last,
  output        auto_out_4_b_ready,
  input         auto_out_4_b_valid,
  input         auto_out_4_b_bits_id,
  input  [1:0]  auto_out_4_b_bits_resp,
  input         auto_out_4_ar_ready,
  output        auto_out_4_ar_valid,
  output        auto_out_4_ar_bits_id,
  output [29:0] auto_out_4_ar_bits_addr,
  output [2:0]  auto_out_4_ar_bits_size,
  output        auto_out_4_r_ready,
  input         auto_out_4_r_valid,
  input         auto_out_4_r_bits_id,
  input  [31:0] auto_out_4_r_bits_data,
  input  [1:0]  auto_out_4_r_bits_resp,
  input         auto_out_4_r_bits_last,
  input         auto_out_3_aw_ready,
  output        auto_out_3_aw_valid,
  output        auto_out_3_aw_bits_id,
  output [29:0] auto_out_3_aw_bits_addr,
  output [2:0]  auto_out_3_aw_bits_size,
  input         auto_out_3_w_ready,
  output        auto_out_3_w_valid,
  output [31:0] auto_out_3_w_bits_data,
  output [3:0]  auto_out_3_w_bits_strb,
  output        auto_out_3_w_bits_last,
  output        auto_out_3_b_ready,
  input         auto_out_3_b_valid,
  input         auto_out_3_b_bits_id,
  input  [1:0]  auto_out_3_b_bits_resp,
  input         auto_out_3_ar_ready,
  output        auto_out_3_ar_valid,
  output        auto_out_3_ar_bits_id,
  output [29:0] auto_out_3_ar_bits_addr,
  output [2:0]  auto_out_3_ar_bits_size,
  output        auto_out_3_r_ready,
  input         auto_out_3_r_valid,
  input         auto_out_3_r_bits_id,
  input  [31:0] auto_out_3_r_bits_data,
  input  [1:0]  auto_out_3_r_bits_resp,
  input         auto_out_3_r_bits_last,
  input         auto_out_2_aw_ready,
  output        auto_out_2_aw_valid,
  output        auto_out_2_aw_bits_id,
  output [29:0] auto_out_2_aw_bits_addr,
  output [2:0]  auto_out_2_aw_bits_size,
  input         auto_out_2_w_ready,
  output        auto_out_2_w_valid,
  output [31:0] auto_out_2_w_bits_data,
  output [3:0]  auto_out_2_w_bits_strb,
  output        auto_out_2_w_bits_last,
  output        auto_out_2_b_ready,
  input         auto_out_2_b_valid,
  input         auto_out_2_b_bits_id,
  input  [1:0]  auto_out_2_b_bits_resp,
  input         auto_out_2_ar_ready,
  output        auto_out_2_ar_valid,
  output        auto_out_2_ar_bits_id,
  output [29:0] auto_out_2_ar_bits_addr,
  output [2:0]  auto_out_2_ar_bits_size,
  output        auto_out_2_r_ready,
  input         auto_out_2_r_valid,
  input         auto_out_2_r_bits_id,
  input  [31:0] auto_out_2_r_bits_data,
  input  [1:0]  auto_out_2_r_bits_resp,
  input         auto_out_2_r_bits_last,
  input         auto_out_1_aw_ready,
  output        auto_out_1_aw_valid,
  output        auto_out_1_aw_bits_id,
  output [29:0] auto_out_1_aw_bits_addr,
  output [2:0]  auto_out_1_aw_bits_size,
  input         auto_out_1_w_ready,
  output        auto_out_1_w_valid,
  output [31:0] auto_out_1_w_bits_data,
  output [3:0]  auto_out_1_w_bits_strb,
  output        auto_out_1_w_bits_last,
  output        auto_out_1_b_ready,
  input         auto_out_1_b_valid,
  input         auto_out_1_b_bits_id,
  input  [1:0]  auto_out_1_b_bits_resp,
  input         auto_out_1_ar_ready,
  output        auto_out_1_ar_valid,
  output        auto_out_1_ar_bits_id,
  output [29:0] auto_out_1_ar_bits_addr,
  output [2:0]  auto_out_1_ar_bits_size,
  output        auto_out_1_r_ready,
  input         auto_out_1_r_valid,
  input         auto_out_1_r_bits_id,
  input  [31:0] auto_out_1_r_bits_data,
  input  [1:0]  auto_out_1_r_bits_resp,
  input         auto_out_1_r_bits_last,
  input         auto_out_0_aw_ready,
  output        auto_out_0_aw_valid,
  output        auto_out_0_aw_bits_id,
  output [29:0] auto_out_0_aw_bits_addr,
  output [2:0]  auto_out_0_aw_bits_size,
  input         auto_out_0_w_ready,
  output        auto_out_0_w_valid,
  output [31:0] auto_out_0_w_bits_data,
  output [3:0]  auto_out_0_w_bits_strb,
  output        auto_out_0_w_bits_last,
  output        auto_out_0_b_ready,
  input         auto_out_0_b_valid,
  input         auto_out_0_b_bits_id,
  input  [1:0]  auto_out_0_b_bits_resp,
  input         auto_out_0_ar_ready,
  output        auto_out_0_ar_valid,
  output        auto_out_0_ar_bits_id,
  output [29:0] auto_out_0_ar_bits_addr,
  output [2:0]  auto_out_0_ar_bits_size,
  output        auto_out_0_r_ready,
  input         auto_out_0_r_valid,
  input         auto_out_0_r_bits_id,
  input  [31:0] auto_out_0_r_bits_data,
  input  [1:0]  auto_out_0_r_bits_resp,
  input         auto_out_0_r_bits_last
);
  wire  awIn_0_clock; // @[Xbar.scala 55:47]
  wire  awIn_0_reset; // @[Xbar.scala 55:47]
  wire  awIn_0_io_enq_ready; // @[Xbar.scala 55:47]
  wire  awIn_0_io_enq_valid; // @[Xbar.scala 55:47]
  wire [21:0] awIn_0_io_enq_bits; // @[Xbar.scala 55:47]
  wire  awIn_0_io_deq_ready; // @[Xbar.scala 55:47]
  wire  awIn_0_io_deq_valid; // @[Xbar.scala 55:47]
  wire [21:0] awIn_0_io_deq_bits; // @[Xbar.scala 55:47]
  wire [30:0] _T_1; // @[Parameters.scala 137:49]
  wire [30:0] _T_3; // @[Parameters.scala 137:52]
  wire  requestARIO_0_0; // @[Parameters.scala 137:67]
  wire [29:0] _T_5; // @[Parameters.scala 137:31]
  wire [30:0] _T_6; // @[Parameters.scala 137:49]
  wire [30:0] _T_8; // @[Parameters.scala 137:52]
  wire  _T_9; // @[Parameters.scala 137:67]
  wire [29:0] _T_10; // @[Parameters.scala 137:31]
  wire [30:0] _T_11; // @[Parameters.scala 137:49]
  wire [30:0] _T_13; // @[Parameters.scala 137:52]
  wire  _T_14; // @[Parameters.scala 137:67]
  wire  requestARIO_0_1; // @[Xbar.scala 52:97]
  wire [29:0] _T_16; // @[Parameters.scala 137:31]
  wire [30:0] _T_17; // @[Parameters.scala 137:49]
  wire [30:0] _T_19; // @[Parameters.scala 137:52]
  wire  requestARIO_0_2; // @[Parameters.scala 137:67]
  wire [29:0] _T_21; // @[Parameters.scala 137:31]
  wire [30:0] _T_22; // @[Parameters.scala 137:49]
  wire [30:0] _T_24; // @[Parameters.scala 137:52]
  wire  requestARIO_0_3; // @[Parameters.scala 137:67]
  wire [29:0] _T_26; // @[Parameters.scala 137:31]
  wire [30:0] _T_27; // @[Parameters.scala 137:49]
  wire [30:0] _T_29; // @[Parameters.scala 137:52]
  wire  requestARIO_0_4; // @[Parameters.scala 137:67]
  wire [29:0] _T_31; // @[Parameters.scala 137:31]
  wire [30:0] _T_32; // @[Parameters.scala 137:49]
  wire [30:0] _T_34; // @[Parameters.scala 137:52]
  wire  requestARIO_0_5; // @[Parameters.scala 137:67]
  wire [29:0] _T_36; // @[Parameters.scala 137:31]
  wire [30:0] _T_37; // @[Parameters.scala 137:49]
  wire [30:0] _T_39; // @[Parameters.scala 137:52]
  wire  requestARIO_0_6; // @[Parameters.scala 137:67]
  wire [29:0] _T_41; // @[Parameters.scala 137:31]
  wire [30:0] _T_42; // @[Parameters.scala 137:49]
  wire [30:0] _T_44; // @[Parameters.scala 137:52]
  wire  requestARIO_0_7; // @[Parameters.scala 137:67]
  wire [29:0] _T_46; // @[Parameters.scala 137:31]
  wire [30:0] _T_47; // @[Parameters.scala 137:49]
  wire [30:0] _T_49; // @[Parameters.scala 137:52]
  wire  requestARIO_0_8; // @[Parameters.scala 137:67]
  wire [29:0] _T_51; // @[Parameters.scala 137:31]
  wire [30:0] _T_52; // @[Parameters.scala 137:49]
  wire [30:0] _T_54; // @[Parameters.scala 137:52]
  wire  requestARIO_0_9; // @[Parameters.scala 137:67]
  wire [29:0] _T_56; // @[Parameters.scala 137:31]
  wire [30:0] _T_57; // @[Parameters.scala 137:49]
  wire [30:0] _T_59; // @[Parameters.scala 137:52]
  wire  requestARIO_0_10; // @[Parameters.scala 137:67]
  wire [29:0] _T_61; // @[Parameters.scala 137:31]
  wire [30:0] _T_62; // @[Parameters.scala 137:49]
  wire [30:0] _T_64; // @[Parameters.scala 137:52]
  wire  requestARIO_0_11; // @[Parameters.scala 137:67]
  wire [29:0] _T_66; // @[Parameters.scala 137:31]
  wire [30:0] _T_67; // @[Parameters.scala 137:49]
  wire [30:0] _T_69; // @[Parameters.scala 137:52]
  wire  requestARIO_0_12; // @[Parameters.scala 137:67]
  wire [29:0] _T_71; // @[Parameters.scala 137:31]
  wire [30:0] _T_72; // @[Parameters.scala 137:49]
  wire [30:0] _T_74; // @[Parameters.scala 137:52]
  wire  requestARIO_0_13; // @[Parameters.scala 137:67]
  wire [29:0] _T_76; // @[Parameters.scala 137:31]
  wire [30:0] _T_77; // @[Parameters.scala 137:49]
  wire [30:0] _T_79; // @[Parameters.scala 137:52]
  wire  requestARIO_0_14; // @[Parameters.scala 137:67]
  wire [29:0] _T_81; // @[Parameters.scala 137:31]
  wire [30:0] _T_82; // @[Parameters.scala 137:49]
  wire [30:0] _T_84; // @[Parameters.scala 137:52]
  wire  requestARIO_0_15; // @[Parameters.scala 137:67]
  wire [29:0] _T_86; // @[Parameters.scala 137:31]
  wire [30:0] _T_87; // @[Parameters.scala 137:49]
  wire [30:0] _T_89; // @[Parameters.scala 137:52]
  wire  requestARIO_0_16; // @[Parameters.scala 137:67]
  wire [29:0] _T_91; // @[Parameters.scala 137:31]
  wire [30:0] _T_92; // @[Parameters.scala 137:49]
  wire [30:0] _T_94; // @[Parameters.scala 137:52]
  wire  requestARIO_0_17; // @[Parameters.scala 137:67]
  wire [29:0] _T_96; // @[Parameters.scala 137:31]
  wire [30:0] _T_97; // @[Parameters.scala 137:49]
  wire [30:0] _T_99; // @[Parameters.scala 137:52]
  wire  requestARIO_0_18; // @[Parameters.scala 137:67]
  wire [29:0] _T_101; // @[Parameters.scala 137:31]
  wire [30:0] _T_102; // @[Parameters.scala 137:49]
  wire [30:0] _T_104; // @[Parameters.scala 137:52]
  wire  requestARIO_0_19; // @[Parameters.scala 137:67]
  wire [29:0] _T_106; // @[Parameters.scala 137:31]
  wire [30:0] _T_107; // @[Parameters.scala 137:49]
  wire [30:0] _T_109; // @[Parameters.scala 137:52]
  wire  requestARIO_0_20; // @[Parameters.scala 137:67]
  wire [29:0] _T_111; // @[Parameters.scala 137:31]
  wire [30:0] _T_112; // @[Parameters.scala 137:49]
  wire [30:0] _T_114; // @[Parameters.scala 137:52]
  wire  _T_115; // @[Parameters.scala 137:67]
  wire [29:0] _T_116; // @[Parameters.scala 137:31]
  wire [30:0] _T_117; // @[Parameters.scala 137:49]
  wire [30:0] _T_119; // @[Parameters.scala 137:52]
  wire  _T_120; // @[Parameters.scala 137:67]
  wire  requestARIO_0_21; // @[Xbar.scala 52:97]
  wire [30:0] _T_123; // @[Parameters.scala 137:49]
  wire [30:0] _T_125; // @[Parameters.scala 137:52]
  wire  requestAWIO_0_0; // @[Parameters.scala 137:67]
  wire [29:0] _T_127; // @[Parameters.scala 137:31]
  wire [30:0] _T_128; // @[Parameters.scala 137:49]
  wire [30:0] _T_130; // @[Parameters.scala 137:52]
  wire  _T_131; // @[Parameters.scala 137:67]
  wire [29:0] _T_132; // @[Parameters.scala 137:31]
  wire [30:0] _T_133; // @[Parameters.scala 137:49]
  wire [30:0] _T_135; // @[Parameters.scala 137:52]
  wire  _T_136; // @[Parameters.scala 137:67]
  wire  requestAWIO_0_1; // @[Xbar.scala 52:97]
  wire [29:0] _T_138; // @[Parameters.scala 137:31]
  wire [30:0] _T_139; // @[Parameters.scala 137:49]
  wire [30:0] _T_141; // @[Parameters.scala 137:52]
  wire  requestAWIO_0_2; // @[Parameters.scala 137:67]
  wire [29:0] _T_143; // @[Parameters.scala 137:31]
  wire [30:0] _T_144; // @[Parameters.scala 137:49]
  wire [30:0] _T_146; // @[Parameters.scala 137:52]
  wire  requestAWIO_0_3; // @[Parameters.scala 137:67]
  wire [29:0] _T_148; // @[Parameters.scala 137:31]
  wire [30:0] _T_149; // @[Parameters.scala 137:49]
  wire [30:0] _T_151; // @[Parameters.scala 137:52]
  wire  requestAWIO_0_4; // @[Parameters.scala 137:67]
  wire [29:0] _T_153; // @[Parameters.scala 137:31]
  wire [30:0] _T_154; // @[Parameters.scala 137:49]
  wire [30:0] _T_156; // @[Parameters.scala 137:52]
  wire  requestAWIO_0_5; // @[Parameters.scala 137:67]
  wire [29:0] _T_158; // @[Parameters.scala 137:31]
  wire [30:0] _T_159; // @[Parameters.scala 137:49]
  wire [30:0] _T_161; // @[Parameters.scala 137:52]
  wire  requestAWIO_0_6; // @[Parameters.scala 137:67]
  wire [29:0] _T_163; // @[Parameters.scala 137:31]
  wire [30:0] _T_164; // @[Parameters.scala 137:49]
  wire [30:0] _T_166; // @[Parameters.scala 137:52]
  wire  requestAWIO_0_7; // @[Parameters.scala 137:67]
  wire [29:0] _T_168; // @[Parameters.scala 137:31]
  wire [30:0] _T_169; // @[Parameters.scala 137:49]
  wire [30:0] _T_171; // @[Parameters.scala 137:52]
  wire  requestAWIO_0_8; // @[Parameters.scala 137:67]
  wire [29:0] _T_173; // @[Parameters.scala 137:31]
  wire [30:0] _T_174; // @[Parameters.scala 137:49]
  wire [30:0] _T_176; // @[Parameters.scala 137:52]
  wire  requestAWIO_0_9; // @[Parameters.scala 137:67]
  wire [29:0] _T_178; // @[Parameters.scala 137:31]
  wire [30:0] _T_179; // @[Parameters.scala 137:49]
  wire [30:0] _T_181; // @[Parameters.scala 137:52]
  wire  requestAWIO_0_10; // @[Parameters.scala 137:67]
  wire [29:0] _T_183; // @[Parameters.scala 137:31]
  wire [30:0] _T_184; // @[Parameters.scala 137:49]
  wire [30:0] _T_186; // @[Parameters.scala 137:52]
  wire  requestAWIO_0_11; // @[Parameters.scala 137:67]
  wire [29:0] _T_188; // @[Parameters.scala 137:31]
  wire [30:0] _T_189; // @[Parameters.scala 137:49]
  wire [30:0] _T_191; // @[Parameters.scala 137:52]
  wire  requestAWIO_0_12; // @[Parameters.scala 137:67]
  wire [29:0] _T_193; // @[Parameters.scala 137:31]
  wire [30:0] _T_194; // @[Parameters.scala 137:49]
  wire [30:0] _T_196; // @[Parameters.scala 137:52]
  wire  requestAWIO_0_13; // @[Parameters.scala 137:67]
  wire [29:0] _T_198; // @[Parameters.scala 137:31]
  wire [30:0] _T_199; // @[Parameters.scala 137:49]
  wire [30:0] _T_201; // @[Parameters.scala 137:52]
  wire  requestAWIO_0_14; // @[Parameters.scala 137:67]
  wire [29:0] _T_203; // @[Parameters.scala 137:31]
  wire [30:0] _T_204; // @[Parameters.scala 137:49]
  wire [30:0] _T_206; // @[Parameters.scala 137:52]
  wire  requestAWIO_0_15; // @[Parameters.scala 137:67]
  wire [29:0] _T_208; // @[Parameters.scala 137:31]
  wire [30:0] _T_209; // @[Parameters.scala 137:49]
  wire [30:0] _T_211; // @[Parameters.scala 137:52]
  wire  requestAWIO_0_16; // @[Parameters.scala 137:67]
  wire [29:0] _T_213; // @[Parameters.scala 137:31]
  wire [30:0] _T_214; // @[Parameters.scala 137:49]
  wire [30:0] _T_216; // @[Parameters.scala 137:52]
  wire  requestAWIO_0_17; // @[Parameters.scala 137:67]
  wire [29:0] _T_218; // @[Parameters.scala 137:31]
  wire [30:0] _T_219; // @[Parameters.scala 137:49]
  wire [30:0] _T_221; // @[Parameters.scala 137:52]
  wire  requestAWIO_0_18; // @[Parameters.scala 137:67]
  wire [29:0] _T_223; // @[Parameters.scala 137:31]
  wire [30:0] _T_224; // @[Parameters.scala 137:49]
  wire [30:0] _T_226; // @[Parameters.scala 137:52]
  wire  requestAWIO_0_19; // @[Parameters.scala 137:67]
  wire [29:0] _T_228; // @[Parameters.scala 137:31]
  wire [30:0] _T_229; // @[Parameters.scala 137:49]
  wire [30:0] _T_231; // @[Parameters.scala 137:52]
  wire  requestAWIO_0_20; // @[Parameters.scala 137:67]
  wire [29:0] _T_233; // @[Parameters.scala 137:31]
  wire [30:0] _T_234; // @[Parameters.scala 137:49]
  wire [30:0] _T_236; // @[Parameters.scala 137:52]
  wire  _T_237; // @[Parameters.scala 137:67]
  wire [29:0] _T_238; // @[Parameters.scala 137:31]
  wire [30:0] _T_239; // @[Parameters.scala 137:49]
  wire [30:0] _T_241; // @[Parameters.scala 137:52]
  wire  _T_242; // @[Parameters.scala 137:67]
  wire  requestAWIO_0_21; // @[Xbar.scala 52:97]
  wire  requestROI_0_0; // @[Parameters.scala 47:9]
  wire  requestROI_1_0; // @[Parameters.scala 47:9]
  wire  requestROI_2_0; // @[Parameters.scala 47:9]
  wire  requestROI_3_0; // @[Parameters.scala 47:9]
  wire  requestROI_4_0; // @[Parameters.scala 47:9]
  wire  requestROI_5_0; // @[Parameters.scala 47:9]
  wire  requestROI_6_0; // @[Parameters.scala 47:9]
  wire  requestROI_7_0; // @[Parameters.scala 47:9]
  wire  requestROI_8_0; // @[Parameters.scala 47:9]
  wire  requestROI_9_0; // @[Parameters.scala 47:9]
  wire  requestROI_10_0; // @[Parameters.scala 47:9]
  wire  requestROI_11_0; // @[Parameters.scala 47:9]
  wire  requestROI_12_0; // @[Parameters.scala 47:9]
  wire  requestROI_13_0; // @[Parameters.scala 47:9]
  wire  requestROI_14_0; // @[Parameters.scala 47:9]
  wire  requestROI_15_0; // @[Parameters.scala 47:9]
  wire  requestROI_16_0; // @[Parameters.scala 47:9]
  wire  requestROI_17_0; // @[Parameters.scala 47:9]
  wire  requestROI_18_0; // @[Parameters.scala 47:9]
  wire  requestROI_19_0; // @[Parameters.scala 47:9]
  wire  requestROI_20_0; // @[Parameters.scala 47:9]
  wire  requestBOI_0_0; // @[Parameters.scala 47:9]
  wire  requestBOI_1_0; // @[Parameters.scala 47:9]
  wire  requestBOI_2_0; // @[Parameters.scala 47:9]
  wire  requestBOI_3_0; // @[Parameters.scala 47:9]
  wire  requestBOI_4_0; // @[Parameters.scala 47:9]
  wire  requestBOI_5_0; // @[Parameters.scala 47:9]
  wire  requestBOI_6_0; // @[Parameters.scala 47:9]
  wire  requestBOI_7_0; // @[Parameters.scala 47:9]
  wire  requestBOI_8_0; // @[Parameters.scala 47:9]
  wire  requestBOI_9_0; // @[Parameters.scala 47:9]
  wire  requestBOI_10_0; // @[Parameters.scala 47:9]
  wire  requestBOI_11_0; // @[Parameters.scala 47:9]
  wire  requestBOI_12_0; // @[Parameters.scala 47:9]
  wire  requestBOI_13_0; // @[Parameters.scala 47:9]
  wire  requestBOI_14_0; // @[Parameters.scala 47:9]
  wire  requestBOI_15_0; // @[Parameters.scala 47:9]
  wire  requestBOI_16_0; // @[Parameters.scala 47:9]
  wire  requestBOI_17_0; // @[Parameters.scala 47:9]
  wire  requestBOI_18_0; // @[Parameters.scala 47:9]
  wire  requestBOI_19_0; // @[Parameters.scala 47:9]
  wire  requestBOI_20_0; // @[Parameters.scala 47:9]
  wire [4:0] _T_247; // @[Xbar.scala 64:75]
  wire [10:0] _T_253; // @[Xbar.scala 64:75]
  wire [4:0] _T_257; // @[Xbar.scala 64:75]
  wire [10:0] _T_263; // @[Xbar.scala 64:75]
  wire [21:0] _T_264; // @[Xbar.scala 64:75]
  wire  requestWIO_0_0; // @[Xbar.scala 65:73]
  wire  requestWIO_0_1; // @[Xbar.scala 65:73]
  wire  requestWIO_0_2; // @[Xbar.scala 65:73]
  wire  requestWIO_0_3; // @[Xbar.scala 65:73]
  wire  requestWIO_0_4; // @[Xbar.scala 65:73]
  wire  requestWIO_0_5; // @[Xbar.scala 65:73]
  wire  requestWIO_0_6; // @[Xbar.scala 65:73]
  wire  requestWIO_0_7; // @[Xbar.scala 65:73]
  wire  requestWIO_0_8; // @[Xbar.scala 65:73]
  wire  requestWIO_0_9; // @[Xbar.scala 65:73]
  wire  requestWIO_0_10; // @[Xbar.scala 65:73]
  wire  requestWIO_0_11; // @[Xbar.scala 65:73]
  wire  requestWIO_0_12; // @[Xbar.scala 65:73]
  wire  requestWIO_0_13; // @[Xbar.scala 65:73]
  wire  requestWIO_0_14; // @[Xbar.scala 65:73]
  wire  requestWIO_0_15; // @[Xbar.scala 65:73]
  wire  requestWIO_0_16; // @[Xbar.scala 65:73]
  wire  requestWIO_0_17; // @[Xbar.scala 65:73]
  wire  requestWIO_0_18; // @[Xbar.scala 65:73]
  wire  requestWIO_0_19; // @[Xbar.scala 65:73]
  wire  requestWIO_0_20; // @[Xbar.scala 65:73]
  wire  requestWIO_0_21; // @[Xbar.scala 65:73]
  wire [4:0] _T_274; // @[Xbar.scala 93:45]
  wire [10:0] _T_280; // @[Xbar.scala 93:45]
  wire [4:0] _T_284; // @[Xbar.scala 93:45]
  wire [21:0] _T_291; // @[Xbar.scala 93:45]
  wire  _T_294; // @[OneHot.scala 32:14]
  wire [15:0] _GEN_98; // @[OneHot.scala 32:28]
  wire [15:0] _T_295; // @[OneHot.scala 32:28]
  wire  _T_298; // @[OneHot.scala 32:14]
  wire [7:0] _T_299; // @[OneHot.scala 32:28]
  wire  _T_302; // @[OneHot.scala 32:14]
  wire [3:0] _T_303; // @[OneHot.scala 32:28]
  wire  _T_306; // @[OneHot.scala 32:14]
  wire [1:0] _T_307; // @[OneHot.scala 32:28]
  wire [4:0] _T_312; // @[Cat.scala 29:58]
  wire  _T_336; // @[OneHot.scala 32:14]
  wire [15:0] _GEN_99; // @[OneHot.scala 32:28]
  wire [15:0] _T_337; // @[OneHot.scala 32:28]
  wire  _T_340; // @[OneHot.scala 32:14]
  wire [7:0] _T_341; // @[OneHot.scala 32:28]
  wire  _T_344; // @[OneHot.scala 32:14]
  wire [3:0] _T_345; // @[OneHot.scala 32:28]
  wire  _T_348; // @[OneHot.scala 32:14]
  wire [1:0] _T_349; // @[OneHot.scala 32:28]
  wire [4:0] _T_354; // @[Cat.scala 29:58]
  wire  _T_452; // @[Mux.scala 27:72]
  wire  _T_453; // @[Mux.scala 27:72]
  wire  _T_474; // @[Mux.scala 27:72]
  wire  _T_454; // @[Mux.scala 27:72]
  wire  _T_475; // @[Mux.scala 27:72]
  wire  _T_455; // @[Mux.scala 27:72]
  wire  _T_476; // @[Mux.scala 27:72]
  wire  _T_456; // @[Mux.scala 27:72]
  wire  _T_477; // @[Mux.scala 27:72]
  wire  _T_457; // @[Mux.scala 27:72]
  wire  _T_478; // @[Mux.scala 27:72]
  wire  _T_458; // @[Mux.scala 27:72]
  wire  _T_479; // @[Mux.scala 27:72]
  wire  _T_459; // @[Mux.scala 27:72]
  wire  _T_480; // @[Mux.scala 27:72]
  wire  _T_460; // @[Mux.scala 27:72]
  wire  _T_481; // @[Mux.scala 27:72]
  wire  _T_461; // @[Mux.scala 27:72]
  wire  _T_482; // @[Mux.scala 27:72]
  wire  _T_462; // @[Mux.scala 27:72]
  wire  _T_483; // @[Mux.scala 27:72]
  wire  _T_463; // @[Mux.scala 27:72]
  wire  _T_484; // @[Mux.scala 27:72]
  wire  _T_464; // @[Mux.scala 27:72]
  wire  _T_485; // @[Mux.scala 27:72]
  wire  _T_465; // @[Mux.scala 27:72]
  wire  _T_486; // @[Mux.scala 27:72]
  wire  _T_466; // @[Mux.scala 27:72]
  wire  _T_487; // @[Mux.scala 27:72]
  wire  _T_467; // @[Mux.scala 27:72]
  wire  _T_488; // @[Mux.scala 27:72]
  wire  _T_468; // @[Mux.scala 27:72]
  wire  _T_489; // @[Mux.scala 27:72]
  wire  _T_469; // @[Mux.scala 27:72]
  wire  _T_490; // @[Mux.scala 27:72]
  wire  _T_470; // @[Mux.scala 27:72]
  wire  _T_491; // @[Mux.scala 27:72]
  wire  _T_471; // @[Mux.scala 27:72]
  wire  _T_492; // @[Mux.scala 27:72]
  wire  _T_472; // @[Mux.scala 27:72]
  wire  _T_493; // @[Mux.scala 27:72]
  wire  _T_473; // @[Mux.scala 27:72]
  wire  in_0_ar_ready; // @[Mux.scala 27:72]
  reg [2:0] _T_360; // @[Xbar.scala 104:34]
  reg [31:0] _RAND_0;
  wire  _T_379; // @[Xbar.scala 112:22]
  reg [4:0] _T_361; // @[Xbar.scala 105:29]
  reg [31:0] _RAND_1;
  wire  _T_378; // @[Xbar.scala 111:75]
  wire  _T_380; // @[Xbar.scala 112:34]
  wire  _T_381; // @[Xbar.scala 112:80]
  wire  _T_383; // @[Xbar.scala 112:48]
  wire  io_in_0_ar_ready; // @[Xbar.scala 130:45]
  wire  _T_355; // @[Decoupled.scala 40:37]
  reg  _T_1686; // @[Xbar.scala 242:23]
  reg [31:0] _RAND_2;
  wire  _T_631; // @[Xbar.scala 222:40]
  wire  _T_633; // @[Xbar.scala 222:40]
  wire  _T_1687; // @[Xbar.scala 246:36]
  wire  _T_635; // @[Xbar.scala 222:40]
  wire  _T_1688; // @[Xbar.scala 246:36]
  wire  _T_637; // @[Xbar.scala 222:40]
  wire  _T_1689; // @[Xbar.scala 246:36]
  wire  _T_639; // @[Xbar.scala 222:40]
  wire  _T_1690; // @[Xbar.scala 246:36]
  wire  _T_641; // @[Xbar.scala 222:40]
  wire  _T_1691; // @[Xbar.scala 246:36]
  wire  _T_643; // @[Xbar.scala 222:40]
  wire  _T_1692; // @[Xbar.scala 246:36]
  wire  _T_645; // @[Xbar.scala 222:40]
  wire  _T_1693; // @[Xbar.scala 246:36]
  wire  _T_647; // @[Xbar.scala 222:40]
  wire  _T_1694; // @[Xbar.scala 246:36]
  wire  _T_649; // @[Xbar.scala 222:40]
  wire  _T_1695; // @[Xbar.scala 246:36]
  wire  _T_651; // @[Xbar.scala 222:40]
  wire  _T_1696; // @[Xbar.scala 246:36]
  wire  _T_653; // @[Xbar.scala 222:40]
  wire  _T_1697; // @[Xbar.scala 246:36]
  wire  _T_655; // @[Xbar.scala 222:40]
  wire  _T_1698; // @[Xbar.scala 246:36]
  wire  _T_657; // @[Xbar.scala 222:40]
  wire  _T_1699; // @[Xbar.scala 246:36]
  wire  _T_659; // @[Xbar.scala 222:40]
  wire  _T_1700; // @[Xbar.scala 246:36]
  wire  _T_661; // @[Xbar.scala 222:40]
  wire  _T_1701; // @[Xbar.scala 246:36]
  wire  _T_663; // @[Xbar.scala 222:40]
  wire  _T_1702; // @[Xbar.scala 246:36]
  wire  _T_665; // @[Xbar.scala 222:40]
  wire  _T_1703; // @[Xbar.scala 246:36]
  wire  _T_667; // @[Xbar.scala 222:40]
  wire  _T_1704; // @[Xbar.scala 246:36]
  wire  _T_669; // @[Xbar.scala 222:40]
  wire  _T_1705; // @[Xbar.scala 246:36]
  wire  _T_671; // @[Xbar.scala 222:40]
  wire  _T_1706; // @[Xbar.scala 246:36]
  wire  _T_1707; // @[Xbar.scala 246:36]
  reg  _T_1962_0; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_3;
  wire  _T_1988; // @[Mux.scala 27:72]
  reg  _T_1962_1; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_4;
  wire  _T_1989; // @[Mux.scala 27:72]
  wire  _T_2010; // @[Mux.scala 27:72]
  reg  _T_1962_2; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_5;
  wire  _T_1990; // @[Mux.scala 27:72]
  wire  _T_2011; // @[Mux.scala 27:72]
  reg  _T_1962_3; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_6;
  wire  _T_1991; // @[Mux.scala 27:72]
  wire  _T_2012; // @[Mux.scala 27:72]
  reg  _T_1962_4; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_7;
  wire  _T_1992; // @[Mux.scala 27:72]
  wire  _T_2013; // @[Mux.scala 27:72]
  reg  _T_1962_5; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_8;
  wire  _T_1993; // @[Mux.scala 27:72]
  wire  _T_2014; // @[Mux.scala 27:72]
  reg  _T_1962_6; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_9;
  wire  _T_1994; // @[Mux.scala 27:72]
  wire  _T_2015; // @[Mux.scala 27:72]
  reg  _T_1962_7; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_10;
  wire  _T_1995; // @[Mux.scala 27:72]
  wire  _T_2016; // @[Mux.scala 27:72]
  reg  _T_1962_8; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_11;
  wire  _T_1996; // @[Mux.scala 27:72]
  wire  _T_2017; // @[Mux.scala 27:72]
  reg  _T_1962_9; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_12;
  wire  _T_1997; // @[Mux.scala 27:72]
  wire  _T_2018; // @[Mux.scala 27:72]
  reg  _T_1962_10; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_13;
  wire  _T_1998; // @[Mux.scala 27:72]
  wire  _T_2019; // @[Mux.scala 27:72]
  reg  _T_1962_11; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_14;
  wire  _T_1999; // @[Mux.scala 27:72]
  wire  _T_2020; // @[Mux.scala 27:72]
  reg  _T_1962_12; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_15;
  wire  _T_2000; // @[Mux.scala 27:72]
  wire  _T_2021; // @[Mux.scala 27:72]
  reg  _T_1962_13; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_16;
  wire  _T_2001; // @[Mux.scala 27:72]
  wire  _T_2022; // @[Mux.scala 27:72]
  reg  _T_1962_14; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_17;
  wire  _T_2002; // @[Mux.scala 27:72]
  wire  _T_2023; // @[Mux.scala 27:72]
  reg  _T_1962_15; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_18;
  wire  _T_2003; // @[Mux.scala 27:72]
  wire  _T_2024; // @[Mux.scala 27:72]
  reg  _T_1962_16; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_19;
  wire  _T_2004; // @[Mux.scala 27:72]
  wire  _T_2025; // @[Mux.scala 27:72]
  reg  _T_1962_17; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_20;
  wire  _T_2005; // @[Mux.scala 27:72]
  wire  _T_2026; // @[Mux.scala 27:72]
  reg  _T_1962_18; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_21;
  wire  _T_2006; // @[Mux.scala 27:72]
  wire  _T_2027; // @[Mux.scala 27:72]
  reg  _T_1962_19; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_22;
  wire  _T_2007; // @[Mux.scala 27:72]
  wire  _T_2028; // @[Mux.scala 27:72]
  reg  _T_1962_20; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_23;
  wire  _T_2008; // @[Mux.scala 27:72]
  wire  _T_2029; // @[Mux.scala 27:72]
  reg  _T_1962_21; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_24;
  wire  _T_2009; // @[Mux.scala 27:72]
  wire  _T_2030; // @[Mux.scala 27:72]
  wire  in_0_r_valid; // @[Xbar.scala 278:22]
  wire  _T_357; // @[Decoupled.scala 40:37]
  wire [4:0] _T_1721; // @[Cat.scala 29:58]
  wire [4:0] _T_1711; // @[Cat.scala 29:58]
  wire [10:0] _T_1717; // @[Cat.scala 29:58]
  wire [21:0] _T_1728; // @[Cat.scala 29:58]
  reg [21:0] _T_1735; // @[Arbiter.scala 20:23]
  reg [31:0] _RAND_25;
  wire [21:0] _T_1736; // @[Arbiter.scala 21:30]
  wire [21:0] _T_1737; // @[Arbiter.scala 21:28]
  wire [43:0] _T_1738; // @[Cat.scala 29:58]
  wire [43:0] _GEN_100; // @[package.scala 208:43]
  wire [43:0] _T_1740; // @[package.scala 208:43]
  wire [43:0] _GEN_101; // @[package.scala 208:43]
  wire [43:0] _T_1742; // @[package.scala 208:43]
  wire [43:0] _GEN_102; // @[package.scala 208:43]
  wire [43:0] _T_1744; // @[package.scala 208:43]
  wire [43:0] _GEN_103; // @[package.scala 208:43]
  wire [43:0] _T_1746; // @[package.scala 208:43]
  wire [43:0] _GEN_104; // @[package.scala 208:43]
  wire [43:0] _T_1748; // @[package.scala 208:43]
  wire [43:0] _T_1751; // @[Arbiter.scala 22:66]
  wire [43:0] _GEN_105; // @[Arbiter.scala 22:58]
  wire [43:0] _T_1752; // @[Arbiter.scala 22:58]
  wire [21:0] _T_1755; // @[Arbiter.scala 23:39]
  wire [21:0] _T_1756; // @[Arbiter.scala 23:18]
  wire  _T_1800; // @[Xbar.scala 250:63]
  wire  _T_1963_0; // @[Xbar.scala 262:23]
  wire [35:0] _T_2035; // @[Mux.scala 27:72]
  wire [35:0] _T_2036; // @[Mux.scala 27:72]
  wire  _T_1801; // @[Xbar.scala 250:63]
  wire  _T_1963_1; // @[Xbar.scala 262:23]
  wire [35:0] _T_2039; // @[Mux.scala 27:72]
  wire [35:0] _T_2040; // @[Mux.scala 27:72]
  wire [35:0] _T_2121; // @[Mux.scala 27:72]
  wire  _T_1802; // @[Xbar.scala 250:63]
  wire  _T_1963_2; // @[Xbar.scala 262:23]
  wire [35:0] _T_2043; // @[Mux.scala 27:72]
  wire [35:0] _T_2044; // @[Mux.scala 27:72]
  wire [35:0] _T_2122; // @[Mux.scala 27:72]
  wire  _T_1803; // @[Xbar.scala 250:63]
  wire  _T_1963_3; // @[Xbar.scala 262:23]
  wire [35:0] _T_2047; // @[Mux.scala 27:72]
  wire [35:0] _T_2048; // @[Mux.scala 27:72]
  wire [35:0] _T_2123; // @[Mux.scala 27:72]
  wire  _T_1804; // @[Xbar.scala 250:63]
  wire  _T_1963_4; // @[Xbar.scala 262:23]
  wire [35:0] _T_2051; // @[Mux.scala 27:72]
  wire [35:0] _T_2052; // @[Mux.scala 27:72]
  wire [35:0] _T_2124; // @[Mux.scala 27:72]
  wire  _T_1805; // @[Xbar.scala 250:63]
  wire  _T_1963_5; // @[Xbar.scala 262:23]
  wire [35:0] _T_2055; // @[Mux.scala 27:72]
  wire [35:0] _T_2056; // @[Mux.scala 27:72]
  wire [35:0] _T_2125; // @[Mux.scala 27:72]
  wire  _T_1806; // @[Xbar.scala 250:63]
  wire  _T_1963_6; // @[Xbar.scala 262:23]
  wire [35:0] _T_2059; // @[Mux.scala 27:72]
  wire [35:0] _T_2060; // @[Mux.scala 27:72]
  wire [35:0] _T_2126; // @[Mux.scala 27:72]
  wire  _T_1807; // @[Xbar.scala 250:63]
  wire  _T_1963_7; // @[Xbar.scala 262:23]
  wire [35:0] _T_2063; // @[Mux.scala 27:72]
  wire [35:0] _T_2064; // @[Mux.scala 27:72]
  wire [35:0] _T_2127; // @[Mux.scala 27:72]
  wire  _T_1808; // @[Xbar.scala 250:63]
  wire  _T_1963_8; // @[Xbar.scala 262:23]
  wire [35:0] _T_2067; // @[Mux.scala 27:72]
  wire [35:0] _T_2068; // @[Mux.scala 27:72]
  wire [35:0] _T_2128; // @[Mux.scala 27:72]
  wire  _T_1809; // @[Xbar.scala 250:63]
  wire  _T_1963_9; // @[Xbar.scala 262:23]
  wire [35:0] _T_2071; // @[Mux.scala 27:72]
  wire [35:0] _T_2072; // @[Mux.scala 27:72]
  wire [35:0] _T_2129; // @[Mux.scala 27:72]
  wire  _T_1810; // @[Xbar.scala 250:63]
  wire  _T_1963_10; // @[Xbar.scala 262:23]
  wire [35:0] _T_2075; // @[Mux.scala 27:72]
  wire [35:0] _T_2076; // @[Mux.scala 27:72]
  wire [35:0] _T_2130; // @[Mux.scala 27:72]
  wire  _T_1811; // @[Xbar.scala 250:63]
  wire  _T_1963_11; // @[Xbar.scala 262:23]
  wire [35:0] _T_2079; // @[Mux.scala 27:72]
  wire [35:0] _T_2080; // @[Mux.scala 27:72]
  wire [35:0] _T_2131; // @[Mux.scala 27:72]
  wire  _T_1812; // @[Xbar.scala 250:63]
  wire  _T_1963_12; // @[Xbar.scala 262:23]
  wire [35:0] _T_2083; // @[Mux.scala 27:72]
  wire [35:0] _T_2084; // @[Mux.scala 27:72]
  wire [35:0] _T_2132; // @[Mux.scala 27:72]
  wire  _T_1813; // @[Xbar.scala 250:63]
  wire  _T_1963_13; // @[Xbar.scala 262:23]
  wire [35:0] _T_2087; // @[Mux.scala 27:72]
  wire [35:0] _T_2088; // @[Mux.scala 27:72]
  wire [35:0] _T_2133; // @[Mux.scala 27:72]
  wire  _T_1814; // @[Xbar.scala 250:63]
  wire  _T_1963_14; // @[Xbar.scala 262:23]
  wire [35:0] _T_2091; // @[Mux.scala 27:72]
  wire [35:0] _T_2092; // @[Mux.scala 27:72]
  wire [35:0] _T_2134; // @[Mux.scala 27:72]
  wire  _T_1815; // @[Xbar.scala 250:63]
  wire  _T_1963_15; // @[Xbar.scala 262:23]
  wire [35:0] _T_2095; // @[Mux.scala 27:72]
  wire [35:0] _T_2096; // @[Mux.scala 27:72]
  wire [35:0] _T_2135; // @[Mux.scala 27:72]
  wire  _T_1816; // @[Xbar.scala 250:63]
  wire  _T_1963_16; // @[Xbar.scala 262:23]
  wire [35:0] _T_2099; // @[Mux.scala 27:72]
  wire [35:0] _T_2100; // @[Mux.scala 27:72]
  wire [35:0] _T_2136; // @[Mux.scala 27:72]
  wire  _T_1817; // @[Xbar.scala 250:63]
  wire  _T_1963_17; // @[Xbar.scala 262:23]
  wire [35:0] _T_2103; // @[Mux.scala 27:72]
  wire [35:0] _T_2104; // @[Mux.scala 27:72]
  wire [35:0] _T_2137; // @[Mux.scala 27:72]
  wire  _T_1818; // @[Xbar.scala 250:63]
  wire  _T_1963_18; // @[Xbar.scala 262:23]
  wire [35:0] _T_2107; // @[Mux.scala 27:72]
  wire [35:0] _T_2108; // @[Mux.scala 27:72]
  wire [35:0] _T_2138; // @[Mux.scala 27:72]
  wire  _T_1819; // @[Xbar.scala 250:63]
  wire  _T_1963_19; // @[Xbar.scala 262:23]
  wire [35:0] _T_2111; // @[Mux.scala 27:72]
  wire [35:0] _T_2112; // @[Mux.scala 27:72]
  wire [35:0] _T_2139; // @[Mux.scala 27:72]
  wire  _T_1820; // @[Xbar.scala 250:63]
  wire  _T_1963_20; // @[Xbar.scala 262:23]
  wire [35:0] _T_2115; // @[Mux.scala 27:72]
  wire [35:0] _T_2116; // @[Mux.scala 27:72]
  wire [35:0] _T_2140; // @[Mux.scala 27:72]
  wire  _T_1821; // @[Xbar.scala 250:63]
  wire  _T_1963_21; // @[Xbar.scala 262:23]
  wire [35:0] _T_2119; // @[Mux.scala 27:72]
  wire [35:0] _T_2120; // @[Mux.scala 27:72]
  wire [35:0] _T_2141; // @[Mux.scala 27:72]
  wire  in_0_r_bits_last; // @[Mux.scala 27:72]
  wire  _T_359; // @[Xbar.scala 120:45]
  wire [2:0] _GEN_106; // @[Xbar.scala 106:30]
  wire [2:0] _T_363; // @[Xbar.scala 106:30]
  wire [2:0] _GEN_107; // @[Xbar.scala 106:48]
  wire [2:0] _T_365; // @[Xbar.scala 106:48]
  wire  _T_366; // @[Xbar.scala 107:23]
  wire  _T_367; // @[Xbar.scala 107:43]
  wire  _T_368; // @[Xbar.scala 107:34]
  wire  _T_370; // @[Xbar.scala 107:22]
  wire  _T_371; // @[Xbar.scala 107:22]
  wire  _T_372; // @[Xbar.scala 108:23]
  wire  _T_374; // @[Xbar.scala 108:34]
  wire  _T_376; // @[Xbar.scala 108:22]
  wire  _T_377; // @[Xbar.scala 108:22]
  wire  _T_519; // @[Mux.scala 27:72]
  wire  _T_520; // @[Mux.scala 27:72]
  wire  _T_541; // @[Mux.scala 27:72]
  wire  _T_521; // @[Mux.scala 27:72]
  wire  _T_542; // @[Mux.scala 27:72]
  wire  _T_522; // @[Mux.scala 27:72]
  wire  _T_543; // @[Mux.scala 27:72]
  wire  _T_523; // @[Mux.scala 27:72]
  wire  _T_544; // @[Mux.scala 27:72]
  wire  _T_524; // @[Mux.scala 27:72]
  wire  _T_545; // @[Mux.scala 27:72]
  wire  _T_525; // @[Mux.scala 27:72]
  wire  _T_546; // @[Mux.scala 27:72]
  wire  _T_526; // @[Mux.scala 27:72]
  wire  _T_547; // @[Mux.scala 27:72]
  wire  _T_527; // @[Mux.scala 27:72]
  wire  _T_548; // @[Mux.scala 27:72]
  wire  _T_528; // @[Mux.scala 27:72]
  wire  _T_549; // @[Mux.scala 27:72]
  wire  _T_529; // @[Mux.scala 27:72]
  wire  _T_550; // @[Mux.scala 27:72]
  wire  _T_530; // @[Mux.scala 27:72]
  wire  _T_551; // @[Mux.scala 27:72]
  wire  _T_531; // @[Mux.scala 27:72]
  wire  _T_552; // @[Mux.scala 27:72]
  wire  _T_532; // @[Mux.scala 27:72]
  wire  _T_553; // @[Mux.scala 27:72]
  wire  _T_533; // @[Mux.scala 27:72]
  wire  _T_554; // @[Mux.scala 27:72]
  wire  _T_534; // @[Mux.scala 27:72]
  wire  _T_555; // @[Mux.scala 27:72]
  wire  _T_535; // @[Mux.scala 27:72]
  wire  _T_556; // @[Mux.scala 27:72]
  wire  _T_536; // @[Mux.scala 27:72]
  wire  _T_557; // @[Mux.scala 27:72]
  wire  _T_537; // @[Mux.scala 27:72]
  wire  _T_558; // @[Mux.scala 27:72]
  wire  _T_538; // @[Mux.scala 27:72]
  wire  _T_559; // @[Mux.scala 27:72]
  wire  _T_539; // @[Mux.scala 27:72]
  wire  _T_560; // @[Mux.scala 27:72]
  wire  _T_540; // @[Mux.scala 27:72]
  wire  in_0_aw_ready; // @[Mux.scala 27:72]
  reg  _T_414; // @[Xbar.scala 137:30]
  reg [31:0] _RAND_26;
  wire  _T_418; // @[Xbar.scala 139:57]
  wire  _T_419; // @[Xbar.scala 139:45]
  reg [2:0] _T_388; // @[Xbar.scala 104:34]
  reg [31:0] _RAND_27;
  wire  _T_407; // @[Xbar.scala 112:22]
  reg [4:0] _T_389; // @[Xbar.scala 105:29]
  reg [31:0] _RAND_28;
  wire  _T_406; // @[Xbar.scala 111:75]
  wire  _T_408; // @[Xbar.scala 112:34]
  wire  _T_409; // @[Xbar.scala 112:80]
  wire  _T_411; // @[Xbar.scala 112:48]
  wire  io_in_0_aw_ready; // @[Xbar.scala 139:82]
  wire  _T_384; // @[Decoupled.scala 40:37]
  reg  _T_2148; // @[Xbar.scala 242:23]
  reg [31:0] _RAND_29;
  wire  _T_675; // @[Xbar.scala 222:40]
  wire  _T_677; // @[Xbar.scala 222:40]
  wire  _T_2149; // @[Xbar.scala 246:36]
  wire  _T_679; // @[Xbar.scala 222:40]
  wire  _T_2150; // @[Xbar.scala 246:36]
  wire  _T_681; // @[Xbar.scala 222:40]
  wire  _T_2151; // @[Xbar.scala 246:36]
  wire  _T_683; // @[Xbar.scala 222:40]
  wire  _T_2152; // @[Xbar.scala 246:36]
  wire  _T_685; // @[Xbar.scala 222:40]
  wire  _T_2153; // @[Xbar.scala 246:36]
  wire  _T_687; // @[Xbar.scala 222:40]
  wire  _T_2154; // @[Xbar.scala 246:36]
  wire  _T_689; // @[Xbar.scala 222:40]
  wire  _T_2155; // @[Xbar.scala 246:36]
  wire  _T_691; // @[Xbar.scala 222:40]
  wire  _T_2156; // @[Xbar.scala 246:36]
  wire  _T_693; // @[Xbar.scala 222:40]
  wire  _T_2157; // @[Xbar.scala 246:36]
  wire  _T_695; // @[Xbar.scala 222:40]
  wire  _T_2158; // @[Xbar.scala 246:36]
  wire  _T_697; // @[Xbar.scala 222:40]
  wire  _T_2159; // @[Xbar.scala 246:36]
  wire  _T_699; // @[Xbar.scala 222:40]
  wire  _T_2160; // @[Xbar.scala 246:36]
  wire  _T_701; // @[Xbar.scala 222:40]
  wire  _T_2161; // @[Xbar.scala 246:36]
  wire  _T_703; // @[Xbar.scala 222:40]
  wire  _T_2162; // @[Xbar.scala 246:36]
  wire  _T_705; // @[Xbar.scala 222:40]
  wire  _T_2163; // @[Xbar.scala 246:36]
  wire  _T_707; // @[Xbar.scala 222:40]
  wire  _T_2164; // @[Xbar.scala 246:36]
  wire  _T_709; // @[Xbar.scala 222:40]
  wire  _T_2165; // @[Xbar.scala 246:36]
  wire  _T_711; // @[Xbar.scala 222:40]
  wire  _T_2166; // @[Xbar.scala 246:36]
  wire  _T_713; // @[Xbar.scala 222:40]
  wire  _T_2167; // @[Xbar.scala 246:36]
  wire  _T_715; // @[Xbar.scala 222:40]
  wire  _T_2168; // @[Xbar.scala 246:36]
  wire  _T_2169; // @[Xbar.scala 246:36]
  reg  _T_2424_0; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_30;
  wire  _T_2450; // @[Mux.scala 27:72]
  reg  _T_2424_1; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_31;
  wire  _T_2451; // @[Mux.scala 27:72]
  wire  _T_2472; // @[Mux.scala 27:72]
  reg  _T_2424_2; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_32;
  wire  _T_2452; // @[Mux.scala 27:72]
  wire  _T_2473; // @[Mux.scala 27:72]
  reg  _T_2424_3; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_33;
  wire  _T_2453; // @[Mux.scala 27:72]
  wire  _T_2474; // @[Mux.scala 27:72]
  reg  _T_2424_4; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_34;
  wire  _T_2454; // @[Mux.scala 27:72]
  wire  _T_2475; // @[Mux.scala 27:72]
  reg  _T_2424_5; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_35;
  wire  _T_2455; // @[Mux.scala 27:72]
  wire  _T_2476; // @[Mux.scala 27:72]
  reg  _T_2424_6; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_36;
  wire  _T_2456; // @[Mux.scala 27:72]
  wire  _T_2477; // @[Mux.scala 27:72]
  reg  _T_2424_7; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_37;
  wire  _T_2457; // @[Mux.scala 27:72]
  wire  _T_2478; // @[Mux.scala 27:72]
  reg  _T_2424_8; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_38;
  wire  _T_2458; // @[Mux.scala 27:72]
  wire  _T_2479; // @[Mux.scala 27:72]
  reg  _T_2424_9; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_39;
  wire  _T_2459; // @[Mux.scala 27:72]
  wire  _T_2480; // @[Mux.scala 27:72]
  reg  _T_2424_10; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_40;
  wire  _T_2460; // @[Mux.scala 27:72]
  wire  _T_2481; // @[Mux.scala 27:72]
  reg  _T_2424_11; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_41;
  wire  _T_2461; // @[Mux.scala 27:72]
  wire  _T_2482; // @[Mux.scala 27:72]
  reg  _T_2424_12; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_42;
  wire  _T_2462; // @[Mux.scala 27:72]
  wire  _T_2483; // @[Mux.scala 27:72]
  reg  _T_2424_13; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_43;
  wire  _T_2463; // @[Mux.scala 27:72]
  wire  _T_2484; // @[Mux.scala 27:72]
  reg  _T_2424_14; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_44;
  wire  _T_2464; // @[Mux.scala 27:72]
  wire  _T_2485; // @[Mux.scala 27:72]
  reg  _T_2424_15; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_45;
  wire  _T_2465; // @[Mux.scala 27:72]
  wire  _T_2486; // @[Mux.scala 27:72]
  reg  _T_2424_16; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_46;
  wire  _T_2466; // @[Mux.scala 27:72]
  wire  _T_2487; // @[Mux.scala 27:72]
  reg  _T_2424_17; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_47;
  wire  _T_2467; // @[Mux.scala 27:72]
  wire  _T_2488; // @[Mux.scala 27:72]
  reg  _T_2424_18; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_48;
  wire  _T_2468; // @[Mux.scala 27:72]
  wire  _T_2489; // @[Mux.scala 27:72]
  reg  _T_2424_19; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_49;
  wire  _T_2469; // @[Mux.scala 27:72]
  wire  _T_2490; // @[Mux.scala 27:72]
  reg  _T_2424_20; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_50;
  wire  _T_2470; // @[Mux.scala 27:72]
  wire  _T_2491; // @[Mux.scala 27:72]
  reg  _T_2424_21; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_51;
  wire  _T_2471; // @[Mux.scala 27:72]
  wire  _T_2492; // @[Mux.scala 27:72]
  wire  in_0_b_valid; // @[Xbar.scala 278:22]
  wire  _T_386; // @[Decoupled.scala 40:37]
  wire [2:0] _GEN_108; // @[Xbar.scala 106:30]
  wire [2:0] _T_391; // @[Xbar.scala 106:30]
  wire [2:0] _GEN_109; // @[Xbar.scala 106:48]
  wire [2:0] _T_393; // @[Xbar.scala 106:48]
  wire  _T_394; // @[Xbar.scala 107:23]
  wire  _T_395; // @[Xbar.scala 107:43]
  wire  _T_396; // @[Xbar.scala 107:34]
  wire  _T_398; // @[Xbar.scala 107:22]
  wire  _T_399; // @[Xbar.scala 107:22]
  wire  _T_400; // @[Xbar.scala 108:23]
  wire  _T_402; // @[Xbar.scala 108:34]
  wire  _T_404; // @[Xbar.scala 108:22]
  wire  _T_405; // @[Xbar.scala 108:22]
  wire  in_0_ar_valid; // @[Xbar.scala 129:45]
  wire  _T_416; // @[Xbar.scala 138:45]
  wire  in_0_aw_valid; // @[Xbar.scala 138:82]
  wire  _T_421; // @[Xbar.scala 140:54]
  wire  _T_423; // @[Decoupled.scala 40:37]
  wire  _GEN_2; // @[Xbar.scala 141:38]
  wire  _T_424; // @[Decoupled.scala 40:37]
  wire  in_0_w_valid; // @[Xbar.scala 145:43]
  wire  _T_586; // @[Mux.scala 27:72]
  wire  _T_587; // @[Mux.scala 27:72]
  wire  _T_608; // @[Mux.scala 27:72]
  wire  _T_588; // @[Mux.scala 27:72]
  wire  _T_609; // @[Mux.scala 27:72]
  wire  _T_589; // @[Mux.scala 27:72]
  wire  _T_610; // @[Mux.scala 27:72]
  wire  _T_590; // @[Mux.scala 27:72]
  wire  _T_611; // @[Mux.scala 27:72]
  wire  _T_591; // @[Mux.scala 27:72]
  wire  _T_612; // @[Mux.scala 27:72]
  wire  _T_592; // @[Mux.scala 27:72]
  wire  _T_613; // @[Mux.scala 27:72]
  wire  _T_593; // @[Mux.scala 27:72]
  wire  _T_614; // @[Mux.scala 27:72]
  wire  _T_594; // @[Mux.scala 27:72]
  wire  _T_615; // @[Mux.scala 27:72]
  wire  _T_595; // @[Mux.scala 27:72]
  wire  _T_616; // @[Mux.scala 27:72]
  wire  _T_596; // @[Mux.scala 27:72]
  wire  _T_617; // @[Mux.scala 27:72]
  wire  _T_597; // @[Mux.scala 27:72]
  wire  _T_618; // @[Mux.scala 27:72]
  wire  _T_598; // @[Mux.scala 27:72]
  wire  _T_619; // @[Mux.scala 27:72]
  wire  _T_599; // @[Mux.scala 27:72]
  wire  _T_620; // @[Mux.scala 27:72]
  wire  _T_600; // @[Mux.scala 27:72]
  wire  _T_621; // @[Mux.scala 27:72]
  wire  _T_601; // @[Mux.scala 27:72]
  wire  _T_622; // @[Mux.scala 27:72]
  wire  _T_602; // @[Mux.scala 27:72]
  wire  _T_623; // @[Mux.scala 27:72]
  wire  _T_603; // @[Mux.scala 27:72]
  wire  _T_624; // @[Mux.scala 27:72]
  wire  _T_604; // @[Mux.scala 27:72]
  wire  _T_625; // @[Mux.scala 27:72]
  wire  _T_605; // @[Mux.scala 27:72]
  wire  _T_626; // @[Mux.scala 27:72]
  wire  _T_606; // @[Mux.scala 27:72]
  wire  _T_627; // @[Mux.scala 27:72]
  wire  _T_607; // @[Mux.scala 27:72]
  wire  in_0_w_ready; // @[Mux.scala 27:72]
  wire  _T_427; // @[Xbar.scala 147:50]
  wire  out_0_ar_valid; // @[Xbar.scala 222:40]
  wire  out_1_ar_valid; // @[Xbar.scala 222:40]
  wire  out_2_ar_valid; // @[Xbar.scala 222:40]
  wire  out_3_ar_valid; // @[Xbar.scala 222:40]
  wire  out_4_ar_valid; // @[Xbar.scala 222:40]
  wire  out_5_ar_valid; // @[Xbar.scala 222:40]
  wire  out_6_ar_valid; // @[Xbar.scala 222:40]
  wire  out_7_ar_valid; // @[Xbar.scala 222:40]
  wire  out_8_ar_valid; // @[Xbar.scala 222:40]
  wire  out_9_ar_valid; // @[Xbar.scala 222:40]
  wire  out_10_ar_valid; // @[Xbar.scala 222:40]
  wire  out_11_ar_valid; // @[Xbar.scala 222:40]
  wire  out_12_ar_valid; // @[Xbar.scala 222:40]
  wire  out_13_ar_valid; // @[Xbar.scala 222:40]
  wire  out_14_ar_valid; // @[Xbar.scala 222:40]
  wire  out_15_ar_valid; // @[Xbar.scala 222:40]
  wire  out_16_ar_valid; // @[Xbar.scala 222:40]
  wire  out_17_ar_valid; // @[Xbar.scala 222:40]
  wire  out_18_ar_valid; // @[Xbar.scala 222:40]
  wire  out_19_ar_valid; // @[Xbar.scala 222:40]
  wire  out_20_ar_valid; // @[Xbar.scala 222:40]
  wire  out_21_ar_valid; // @[Xbar.scala 222:40]
  wire  out_0_aw_valid; // @[Xbar.scala 222:40]
  wire  out_1_aw_valid; // @[Xbar.scala 222:40]
  wire  out_2_aw_valid; // @[Xbar.scala 222:40]
  wire  out_3_aw_valid; // @[Xbar.scala 222:40]
  wire  out_4_aw_valid; // @[Xbar.scala 222:40]
  wire  out_5_aw_valid; // @[Xbar.scala 222:40]
  wire  out_6_aw_valid; // @[Xbar.scala 222:40]
  wire  out_7_aw_valid; // @[Xbar.scala 222:40]
  wire  out_8_aw_valid; // @[Xbar.scala 222:40]
  wire  out_9_aw_valid; // @[Xbar.scala 222:40]
  wire  out_10_aw_valid; // @[Xbar.scala 222:40]
  wire  out_11_aw_valid; // @[Xbar.scala 222:40]
  wire  out_12_aw_valid; // @[Xbar.scala 222:40]
  wire  out_13_aw_valid; // @[Xbar.scala 222:40]
  wire  out_14_aw_valid; // @[Xbar.scala 222:40]
  wire  out_15_aw_valid; // @[Xbar.scala 222:40]
  wire  out_16_aw_valid; // @[Xbar.scala 222:40]
  wire  out_17_aw_valid; // @[Xbar.scala 222:40]
  wire  out_18_aw_valid; // @[Xbar.scala 222:40]
  wire  out_19_aw_valid; // @[Xbar.scala 222:40]
  wire  out_20_aw_valid; // @[Xbar.scala 222:40]
  wire  out_21_aw_valid; // @[Xbar.scala 222:40]
  wire  _T_724; // @[Xbar.scala 256:60]
  wire  _T_730; // @[Xbar.scala 258:23]
  wire  _T_732; // @[Xbar.scala 258:12]
  wire  _T_733; // @[Xbar.scala 258:12]
  wire  _T_745; // @[Xbar.scala 256:60]
  wire  _T_751; // @[Xbar.scala 258:23]
  wire  _T_753; // @[Xbar.scala 258:12]
  wire  _T_754; // @[Xbar.scala 258:12]
  wire  _T_768; // @[Xbar.scala 256:60]
  wire  _T_774; // @[Xbar.scala 258:23]
  wire  _T_776; // @[Xbar.scala 258:12]
  wire  _T_777; // @[Xbar.scala 258:12]
  wire  _T_789; // @[Xbar.scala 256:60]
  wire  _T_795; // @[Xbar.scala 258:23]
  wire  _T_797; // @[Xbar.scala 258:12]
  wire  _T_798; // @[Xbar.scala 258:12]
  wire  _T_812; // @[Xbar.scala 256:60]
  wire  _T_818; // @[Xbar.scala 258:23]
  wire  _T_820; // @[Xbar.scala 258:12]
  wire  _T_821; // @[Xbar.scala 258:12]
  wire  _T_833; // @[Xbar.scala 256:60]
  wire  _T_839; // @[Xbar.scala 258:23]
  wire  _T_841; // @[Xbar.scala 258:12]
  wire  _T_842; // @[Xbar.scala 258:12]
  wire  _T_856; // @[Xbar.scala 256:60]
  wire  _T_862; // @[Xbar.scala 258:23]
  wire  _T_864; // @[Xbar.scala 258:12]
  wire  _T_865; // @[Xbar.scala 258:12]
  wire  _T_877; // @[Xbar.scala 256:60]
  wire  _T_883; // @[Xbar.scala 258:23]
  wire  _T_885; // @[Xbar.scala 258:12]
  wire  _T_886; // @[Xbar.scala 258:12]
  wire  _T_900; // @[Xbar.scala 256:60]
  wire  _T_906; // @[Xbar.scala 258:23]
  wire  _T_908; // @[Xbar.scala 258:12]
  wire  _T_909; // @[Xbar.scala 258:12]
  wire  _T_921; // @[Xbar.scala 256:60]
  wire  _T_927; // @[Xbar.scala 258:23]
  wire  _T_929; // @[Xbar.scala 258:12]
  wire  _T_930; // @[Xbar.scala 258:12]
  wire  _T_944; // @[Xbar.scala 256:60]
  wire  _T_950; // @[Xbar.scala 258:23]
  wire  _T_952; // @[Xbar.scala 258:12]
  wire  _T_953; // @[Xbar.scala 258:12]
  wire  _T_965; // @[Xbar.scala 256:60]
  wire  _T_971; // @[Xbar.scala 258:23]
  wire  _T_973; // @[Xbar.scala 258:12]
  wire  _T_974; // @[Xbar.scala 258:12]
  wire  _T_988; // @[Xbar.scala 256:60]
  wire  _T_994; // @[Xbar.scala 258:23]
  wire  _T_996; // @[Xbar.scala 258:12]
  wire  _T_997; // @[Xbar.scala 258:12]
  wire  _T_1009; // @[Xbar.scala 256:60]
  wire  _T_1015; // @[Xbar.scala 258:23]
  wire  _T_1017; // @[Xbar.scala 258:12]
  wire  _T_1018; // @[Xbar.scala 258:12]
  wire  _T_1032; // @[Xbar.scala 256:60]
  wire  _T_1038; // @[Xbar.scala 258:23]
  wire  _T_1040; // @[Xbar.scala 258:12]
  wire  _T_1041; // @[Xbar.scala 258:12]
  wire  _T_1053; // @[Xbar.scala 256:60]
  wire  _T_1059; // @[Xbar.scala 258:23]
  wire  _T_1061; // @[Xbar.scala 258:12]
  wire  _T_1062; // @[Xbar.scala 258:12]
  wire  _T_1076; // @[Xbar.scala 256:60]
  wire  _T_1082; // @[Xbar.scala 258:23]
  wire  _T_1084; // @[Xbar.scala 258:12]
  wire  _T_1085; // @[Xbar.scala 258:12]
  wire  _T_1097; // @[Xbar.scala 256:60]
  wire  _T_1103; // @[Xbar.scala 258:23]
  wire  _T_1105; // @[Xbar.scala 258:12]
  wire  _T_1106; // @[Xbar.scala 258:12]
  wire  _T_1120; // @[Xbar.scala 256:60]
  wire  _T_1126; // @[Xbar.scala 258:23]
  wire  _T_1128; // @[Xbar.scala 258:12]
  wire  _T_1129; // @[Xbar.scala 258:12]
  wire  _T_1141; // @[Xbar.scala 256:60]
  wire  _T_1147; // @[Xbar.scala 258:23]
  wire  _T_1149; // @[Xbar.scala 258:12]
  wire  _T_1150; // @[Xbar.scala 258:12]
  wire  _T_1164; // @[Xbar.scala 256:60]
  wire  _T_1170; // @[Xbar.scala 258:23]
  wire  _T_1172; // @[Xbar.scala 258:12]
  wire  _T_1173; // @[Xbar.scala 258:12]
  wire  _T_1185; // @[Xbar.scala 256:60]
  wire  _T_1191; // @[Xbar.scala 258:23]
  wire  _T_1193; // @[Xbar.scala 258:12]
  wire  _T_1194; // @[Xbar.scala 258:12]
  wire  _T_1208; // @[Xbar.scala 256:60]
  wire  _T_1214; // @[Xbar.scala 258:23]
  wire  _T_1216; // @[Xbar.scala 258:12]
  wire  _T_1217; // @[Xbar.scala 258:12]
  wire  _T_1229; // @[Xbar.scala 256:60]
  wire  _T_1235; // @[Xbar.scala 258:23]
  wire  _T_1237; // @[Xbar.scala 258:12]
  wire  _T_1238; // @[Xbar.scala 258:12]
  wire  _T_1252; // @[Xbar.scala 256:60]
  wire  _T_1258; // @[Xbar.scala 258:23]
  wire  _T_1260; // @[Xbar.scala 258:12]
  wire  _T_1261; // @[Xbar.scala 258:12]
  wire  _T_1273; // @[Xbar.scala 256:60]
  wire  _T_1279; // @[Xbar.scala 258:23]
  wire  _T_1281; // @[Xbar.scala 258:12]
  wire  _T_1282; // @[Xbar.scala 258:12]
  wire  _T_1296; // @[Xbar.scala 256:60]
  wire  _T_1302; // @[Xbar.scala 258:23]
  wire  _T_1304; // @[Xbar.scala 258:12]
  wire  _T_1305; // @[Xbar.scala 258:12]
  wire  _T_1317; // @[Xbar.scala 256:60]
  wire  _T_1323; // @[Xbar.scala 258:23]
  wire  _T_1325; // @[Xbar.scala 258:12]
  wire  _T_1326; // @[Xbar.scala 258:12]
  wire  _T_1340; // @[Xbar.scala 256:60]
  wire  _T_1346; // @[Xbar.scala 258:23]
  wire  _T_1348; // @[Xbar.scala 258:12]
  wire  _T_1349; // @[Xbar.scala 258:12]
  wire  _T_1361; // @[Xbar.scala 256:60]
  wire  _T_1367; // @[Xbar.scala 258:23]
  wire  _T_1369; // @[Xbar.scala 258:12]
  wire  _T_1370; // @[Xbar.scala 258:12]
  wire  _T_1384; // @[Xbar.scala 256:60]
  wire  _T_1390; // @[Xbar.scala 258:23]
  wire  _T_1392; // @[Xbar.scala 258:12]
  wire  _T_1393; // @[Xbar.scala 258:12]
  wire  _T_1405; // @[Xbar.scala 256:60]
  wire  _T_1411; // @[Xbar.scala 258:23]
  wire  _T_1413; // @[Xbar.scala 258:12]
  wire  _T_1414; // @[Xbar.scala 258:12]
  wire  _T_1428; // @[Xbar.scala 256:60]
  wire  _T_1434; // @[Xbar.scala 258:23]
  wire  _T_1436; // @[Xbar.scala 258:12]
  wire  _T_1437; // @[Xbar.scala 258:12]
  wire  _T_1449; // @[Xbar.scala 256:60]
  wire  _T_1455; // @[Xbar.scala 258:23]
  wire  _T_1457; // @[Xbar.scala 258:12]
  wire  _T_1458; // @[Xbar.scala 258:12]
  wire  _T_1472; // @[Xbar.scala 256:60]
  wire  _T_1478; // @[Xbar.scala 258:23]
  wire  _T_1480; // @[Xbar.scala 258:12]
  wire  _T_1481; // @[Xbar.scala 258:12]
  wire  _T_1493; // @[Xbar.scala 256:60]
  wire  _T_1499; // @[Xbar.scala 258:23]
  wire  _T_1501; // @[Xbar.scala 258:12]
  wire  _T_1502; // @[Xbar.scala 258:12]
  wire  _T_1516; // @[Xbar.scala 256:60]
  wire  _T_1522; // @[Xbar.scala 258:23]
  wire  _T_1524; // @[Xbar.scala 258:12]
  wire  _T_1525; // @[Xbar.scala 258:12]
  wire  _T_1537; // @[Xbar.scala 256:60]
  wire  _T_1543; // @[Xbar.scala 258:23]
  wire  _T_1545; // @[Xbar.scala 258:12]
  wire  _T_1546; // @[Xbar.scala 258:12]
  wire  _T_1560; // @[Xbar.scala 256:60]
  wire  _T_1566; // @[Xbar.scala 258:23]
  wire  _T_1568; // @[Xbar.scala 258:12]
  wire  _T_1569; // @[Xbar.scala 258:12]
  wire  _T_1581; // @[Xbar.scala 256:60]
  wire  _T_1587; // @[Xbar.scala 258:23]
  wire  _T_1589; // @[Xbar.scala 258:12]
  wire  _T_1590; // @[Xbar.scala 258:12]
  wire  _T_1604; // @[Xbar.scala 256:60]
  wire  _T_1610; // @[Xbar.scala 258:23]
  wire  _T_1612; // @[Xbar.scala 258:12]
  wire  _T_1613; // @[Xbar.scala 258:12]
  wire  _T_1625; // @[Xbar.scala 256:60]
  wire  _T_1631; // @[Xbar.scala 258:23]
  wire  _T_1633; // @[Xbar.scala 258:12]
  wire  _T_1634; // @[Xbar.scala 258:12]
  wire  _T_1648; // @[Xbar.scala 256:60]
  wire  _T_1654; // @[Xbar.scala 258:23]
  wire  _T_1656; // @[Xbar.scala 258:12]
  wire  _T_1657; // @[Xbar.scala 258:12]
  wire  _T_1669; // @[Xbar.scala 256:60]
  wire  _T_1675; // @[Xbar.scala 258:23]
  wire  _T_1677; // @[Xbar.scala 258:12]
  wire  _T_1678; // @[Xbar.scala 258:12]
  wire  _T_1757; // @[Arbiter.scala 24:27]
  wire  _T_1758; // @[Arbiter.scala 24:18]
  wire [21:0] _T_1759; // @[Arbiter.scala 25:29]
  wire [22:0] _T_1760; // @[package.scala 199:48]
  wire [21:0] _T_1762; // @[package.scala 199:43]
  wire [23:0] _T_1763; // @[package.scala 199:48]
  wire [21:0] _T_1765; // @[package.scala 199:43]
  wire [25:0] _T_1766; // @[package.scala 199:48]
  wire [21:0] _T_1768; // @[package.scala 199:43]
  wire [29:0] _T_1769; // @[package.scala 199:48]
  wire [21:0] _T_1771; // @[package.scala 199:43]
  wire [37:0] _T_1772; // @[package.scala 199:48]
  wire [21:0] _T_1774; // @[package.scala 199:43]
  wire  _T_1824; // @[Xbar.scala 255:50]
  wire  _T_1825; // @[Xbar.scala 255:50]
  wire  _T_1826; // @[Xbar.scala 255:50]
  wire  _T_1827; // @[Xbar.scala 255:50]
  wire  _T_1828; // @[Xbar.scala 255:50]
  wire  _T_1829; // @[Xbar.scala 255:50]
  wire  _T_1830; // @[Xbar.scala 255:50]
  wire  _T_1831; // @[Xbar.scala 255:50]
  wire  _T_1832; // @[Xbar.scala 255:50]
  wire  _T_1833; // @[Xbar.scala 255:50]
  wire  _T_1834; // @[Xbar.scala 255:50]
  wire  _T_1835; // @[Xbar.scala 255:50]
  wire  _T_1836; // @[Xbar.scala 255:50]
  wire  _T_1837; // @[Xbar.scala 255:50]
  wire  _T_1838; // @[Xbar.scala 255:50]
  wire  _T_1839; // @[Xbar.scala 255:50]
  wire  _T_1840; // @[Xbar.scala 255:50]
  wire  _T_1841; // @[Xbar.scala 255:50]
  wire  _T_1842; // @[Xbar.scala 255:50]
  wire  _T_1843; // @[Xbar.scala 255:50]
  wire  _T_1844; // @[Xbar.scala 255:50]
  wire  _T_1846; // @[Xbar.scala 256:60]
  wire  _T_1849; // @[Xbar.scala 256:60]
  wire  _T_1850; // @[Xbar.scala 256:57]
  wire  _T_1851; // @[Xbar.scala 256:54]
  wire  _T_1852; // @[Xbar.scala 256:60]
  wire  _T_1853; // @[Xbar.scala 256:57]
  wire  _T_1854; // @[Xbar.scala 256:54]
  wire  _T_1855; // @[Xbar.scala 256:60]
  wire  _T_1856; // @[Xbar.scala 256:57]
  wire  _T_1857; // @[Xbar.scala 256:54]
  wire  _T_1858; // @[Xbar.scala 256:60]
  wire  _T_1859; // @[Xbar.scala 256:57]
  wire  _T_1860; // @[Xbar.scala 256:54]
  wire  _T_1861; // @[Xbar.scala 256:60]
  wire  _T_1862; // @[Xbar.scala 256:57]
  wire  _T_1863; // @[Xbar.scala 256:54]
  wire  _T_1864; // @[Xbar.scala 256:60]
  wire  _T_1865; // @[Xbar.scala 256:57]
  wire  _T_1866; // @[Xbar.scala 256:54]
  wire  _T_1867; // @[Xbar.scala 256:60]
  wire  _T_1868; // @[Xbar.scala 256:57]
  wire  _T_1869; // @[Xbar.scala 256:54]
  wire  _T_1870; // @[Xbar.scala 256:60]
  wire  _T_1871; // @[Xbar.scala 256:57]
  wire  _T_1872; // @[Xbar.scala 256:54]
  wire  _T_1873; // @[Xbar.scala 256:60]
  wire  _T_1874; // @[Xbar.scala 256:57]
  wire  _T_1875; // @[Xbar.scala 256:54]
  wire  _T_1876; // @[Xbar.scala 256:60]
  wire  _T_1877; // @[Xbar.scala 256:57]
  wire  _T_1878; // @[Xbar.scala 256:54]
  wire  _T_1879; // @[Xbar.scala 256:60]
  wire  _T_1880; // @[Xbar.scala 256:57]
  wire  _T_1881; // @[Xbar.scala 256:54]
  wire  _T_1882; // @[Xbar.scala 256:60]
  wire  _T_1883; // @[Xbar.scala 256:57]
  wire  _T_1884; // @[Xbar.scala 256:54]
  wire  _T_1885; // @[Xbar.scala 256:60]
  wire  _T_1886; // @[Xbar.scala 256:57]
  wire  _T_1887; // @[Xbar.scala 256:54]
  wire  _T_1888; // @[Xbar.scala 256:60]
  wire  _T_1889; // @[Xbar.scala 256:57]
  wire  _T_1890; // @[Xbar.scala 256:54]
  wire  _T_1891; // @[Xbar.scala 256:60]
  wire  _T_1892; // @[Xbar.scala 256:57]
  wire  _T_1893; // @[Xbar.scala 256:54]
  wire  _T_1894; // @[Xbar.scala 256:60]
  wire  _T_1895; // @[Xbar.scala 256:57]
  wire  _T_1896; // @[Xbar.scala 256:54]
  wire  _T_1897; // @[Xbar.scala 256:60]
  wire  _T_1898; // @[Xbar.scala 256:57]
  wire  _T_1899; // @[Xbar.scala 256:54]
  wire  _T_1900; // @[Xbar.scala 256:60]
  wire  _T_1901; // @[Xbar.scala 256:57]
  wire  _T_1902; // @[Xbar.scala 256:54]
  wire  _T_1903; // @[Xbar.scala 256:60]
  wire  _T_1904; // @[Xbar.scala 256:57]
  wire  _T_1905; // @[Xbar.scala 256:54]
  wire  _T_1906; // @[Xbar.scala 256:60]
  wire  _T_1907; // @[Xbar.scala 256:57]
  wire  _T_1908; // @[Xbar.scala 256:54]
  wire  _T_1909; // @[Xbar.scala 256:60]
  wire  _T_1910; // @[Xbar.scala 256:57]
  wire  _T_1912; // @[Xbar.scala 256:75]
  wire  _T_1913; // @[Xbar.scala 256:75]
  wire  _T_1914; // @[Xbar.scala 256:75]
  wire  _T_1915; // @[Xbar.scala 256:75]
  wire  _T_1916; // @[Xbar.scala 256:75]
  wire  _T_1917; // @[Xbar.scala 256:75]
  wire  _T_1918; // @[Xbar.scala 256:75]
  wire  _T_1919; // @[Xbar.scala 256:75]
  wire  _T_1920; // @[Xbar.scala 256:75]
  wire  _T_1921; // @[Xbar.scala 256:75]
  wire  _T_1922; // @[Xbar.scala 256:75]
  wire  _T_1923; // @[Xbar.scala 256:75]
  wire  _T_1924; // @[Xbar.scala 256:75]
  wire  _T_1925; // @[Xbar.scala 256:75]
  wire  _T_1926; // @[Xbar.scala 256:75]
  wire  _T_1927; // @[Xbar.scala 256:75]
  wire  _T_1928; // @[Xbar.scala 256:75]
  wire  _T_1929; // @[Xbar.scala 256:75]
  wire  _T_1930; // @[Xbar.scala 256:75]
  wire  _T_1931; // @[Xbar.scala 256:75]
  wire  _T_1933; // @[Xbar.scala 256:11]
  wire  _T_1934; // @[Xbar.scala 256:11]
  wire  _T_1935; // @[Xbar.scala 258:13]
  wire  _T_1957; // @[Xbar.scala 258:23]
  wire  _T_1959; // @[Xbar.scala 258:12]
  wire  _T_1960; // @[Xbar.scala 258:12]
  wire  _GEN_93; // @[Xbar.scala 266:21]
  wire  _GEN_94; // @[Xbar.scala 267:24]
  wire  _T_1965_0; // @[Xbar.scala 270:24]
  wire  _T_1965_1; // @[Xbar.scala 270:24]
  wire  _T_1965_2; // @[Xbar.scala 270:24]
  wire  _T_1965_3; // @[Xbar.scala 270:24]
  wire  _T_1965_4; // @[Xbar.scala 270:24]
  wire  _T_1965_5; // @[Xbar.scala 270:24]
  wire  _T_1965_6; // @[Xbar.scala 270:24]
  wire  _T_1965_7; // @[Xbar.scala 270:24]
  wire  _T_1965_8; // @[Xbar.scala 270:24]
  wire  _T_1965_9; // @[Xbar.scala 270:24]
  wire  _T_1965_10; // @[Xbar.scala 270:24]
  wire  _T_1965_11; // @[Xbar.scala 270:24]
  wire  _T_1965_12; // @[Xbar.scala 270:24]
  wire  _T_1965_13; // @[Xbar.scala 270:24]
  wire  _T_1965_14; // @[Xbar.scala 270:24]
  wire  _T_1965_15; // @[Xbar.scala 270:24]
  wire  _T_1965_16; // @[Xbar.scala 270:24]
  wire  _T_1965_17; // @[Xbar.scala 270:24]
  wire  _T_1965_18; // @[Xbar.scala 270:24]
  wire  _T_1965_19; // @[Xbar.scala 270:24]
  wire  _T_1965_20; // @[Xbar.scala 270:24]
  wire  _T_1965_21; // @[Xbar.scala 270:24]
  wire [4:0] _T_2173; // @[Cat.scala 29:58]
  wire [10:0] _T_2179; // @[Cat.scala 29:58]
  wire [4:0] _T_2183; // @[Cat.scala 29:58]
  wire [21:0] _T_2190; // @[Cat.scala 29:58]
  reg [21:0] _T_2197; // @[Arbiter.scala 20:23]
  reg [31:0] _RAND_52;
  wire [21:0] _T_2198; // @[Arbiter.scala 21:30]
  wire [21:0] _T_2199; // @[Arbiter.scala 21:28]
  wire [43:0] _T_2200; // @[Cat.scala 29:58]
  wire [43:0] _GEN_110; // @[package.scala 208:43]
  wire [43:0] _T_2202; // @[package.scala 208:43]
  wire [43:0] _GEN_111; // @[package.scala 208:43]
  wire [43:0] _T_2204; // @[package.scala 208:43]
  wire [43:0] _GEN_112; // @[package.scala 208:43]
  wire [43:0] _T_2206; // @[package.scala 208:43]
  wire [43:0] _GEN_113; // @[package.scala 208:43]
  wire [43:0] _T_2208; // @[package.scala 208:43]
  wire [43:0] _GEN_114; // @[package.scala 208:43]
  wire [43:0] _T_2210; // @[package.scala 208:43]
  wire [43:0] _T_2213; // @[Arbiter.scala 22:66]
  wire [43:0] _GEN_115; // @[Arbiter.scala 22:58]
  wire [43:0] _T_2214; // @[Arbiter.scala 22:58]
  wire [21:0] _T_2217; // @[Arbiter.scala 23:39]
  wire [21:0] _T_2218; // @[Arbiter.scala 23:18]
  wire  _T_2219; // @[Arbiter.scala 24:27]
  wire  _T_2220; // @[Arbiter.scala 24:18]
  wire [21:0] _T_2221; // @[Arbiter.scala 25:29]
  wire [22:0] _T_2222; // @[package.scala 199:48]
  wire [21:0] _T_2224; // @[package.scala 199:43]
  wire [23:0] _T_2225; // @[package.scala 199:48]
  wire [21:0] _T_2227; // @[package.scala 199:43]
  wire [25:0] _T_2228; // @[package.scala 199:48]
  wire [21:0] _T_2230; // @[package.scala 199:43]
  wire [29:0] _T_2231; // @[package.scala 199:48]
  wire [21:0] _T_2233; // @[package.scala 199:43]
  wire [37:0] _T_2234; // @[package.scala 199:48]
  wire [21:0] _T_2236; // @[package.scala 199:43]
  wire  _T_2262; // @[Xbar.scala 250:63]
  wire  _T_2263; // @[Xbar.scala 250:63]
  wire  _T_2264; // @[Xbar.scala 250:63]
  wire  _T_2265; // @[Xbar.scala 250:63]
  wire  _T_2266; // @[Xbar.scala 250:63]
  wire  _T_2267; // @[Xbar.scala 250:63]
  wire  _T_2268; // @[Xbar.scala 250:63]
  wire  _T_2269; // @[Xbar.scala 250:63]
  wire  _T_2270; // @[Xbar.scala 250:63]
  wire  _T_2271; // @[Xbar.scala 250:63]
  wire  _T_2272; // @[Xbar.scala 250:63]
  wire  _T_2273; // @[Xbar.scala 250:63]
  wire  _T_2274; // @[Xbar.scala 250:63]
  wire  _T_2275; // @[Xbar.scala 250:63]
  wire  _T_2276; // @[Xbar.scala 250:63]
  wire  _T_2277; // @[Xbar.scala 250:63]
  wire  _T_2278; // @[Xbar.scala 250:63]
  wire  _T_2279; // @[Xbar.scala 250:63]
  wire  _T_2280; // @[Xbar.scala 250:63]
  wire  _T_2281; // @[Xbar.scala 250:63]
  wire  _T_2282; // @[Xbar.scala 250:63]
  wire  _T_2283; // @[Xbar.scala 250:63]
  wire  _T_2286; // @[Xbar.scala 255:50]
  wire  _T_2287; // @[Xbar.scala 255:50]
  wire  _T_2288; // @[Xbar.scala 255:50]
  wire  _T_2289; // @[Xbar.scala 255:50]
  wire  _T_2290; // @[Xbar.scala 255:50]
  wire  _T_2291; // @[Xbar.scala 255:50]
  wire  _T_2292; // @[Xbar.scala 255:50]
  wire  _T_2293; // @[Xbar.scala 255:50]
  wire  _T_2294; // @[Xbar.scala 255:50]
  wire  _T_2295; // @[Xbar.scala 255:50]
  wire  _T_2296; // @[Xbar.scala 255:50]
  wire  _T_2297; // @[Xbar.scala 255:50]
  wire  _T_2298; // @[Xbar.scala 255:50]
  wire  _T_2299; // @[Xbar.scala 255:50]
  wire  _T_2300; // @[Xbar.scala 255:50]
  wire  _T_2301; // @[Xbar.scala 255:50]
  wire  _T_2302; // @[Xbar.scala 255:50]
  wire  _T_2303; // @[Xbar.scala 255:50]
  wire  _T_2304; // @[Xbar.scala 255:50]
  wire  _T_2305; // @[Xbar.scala 255:50]
  wire  _T_2306; // @[Xbar.scala 255:50]
  wire  _T_2308; // @[Xbar.scala 256:60]
  wire  _T_2311; // @[Xbar.scala 256:60]
  wire  _T_2312; // @[Xbar.scala 256:57]
  wire  _T_2313; // @[Xbar.scala 256:54]
  wire  _T_2314; // @[Xbar.scala 256:60]
  wire  _T_2315; // @[Xbar.scala 256:57]
  wire  _T_2316; // @[Xbar.scala 256:54]
  wire  _T_2317; // @[Xbar.scala 256:60]
  wire  _T_2318; // @[Xbar.scala 256:57]
  wire  _T_2319; // @[Xbar.scala 256:54]
  wire  _T_2320; // @[Xbar.scala 256:60]
  wire  _T_2321; // @[Xbar.scala 256:57]
  wire  _T_2322; // @[Xbar.scala 256:54]
  wire  _T_2323; // @[Xbar.scala 256:60]
  wire  _T_2324; // @[Xbar.scala 256:57]
  wire  _T_2325; // @[Xbar.scala 256:54]
  wire  _T_2326; // @[Xbar.scala 256:60]
  wire  _T_2327; // @[Xbar.scala 256:57]
  wire  _T_2328; // @[Xbar.scala 256:54]
  wire  _T_2329; // @[Xbar.scala 256:60]
  wire  _T_2330; // @[Xbar.scala 256:57]
  wire  _T_2331; // @[Xbar.scala 256:54]
  wire  _T_2332; // @[Xbar.scala 256:60]
  wire  _T_2333; // @[Xbar.scala 256:57]
  wire  _T_2334; // @[Xbar.scala 256:54]
  wire  _T_2335; // @[Xbar.scala 256:60]
  wire  _T_2336; // @[Xbar.scala 256:57]
  wire  _T_2337; // @[Xbar.scala 256:54]
  wire  _T_2338; // @[Xbar.scala 256:60]
  wire  _T_2339; // @[Xbar.scala 256:57]
  wire  _T_2340; // @[Xbar.scala 256:54]
  wire  _T_2341; // @[Xbar.scala 256:60]
  wire  _T_2342; // @[Xbar.scala 256:57]
  wire  _T_2343; // @[Xbar.scala 256:54]
  wire  _T_2344; // @[Xbar.scala 256:60]
  wire  _T_2345; // @[Xbar.scala 256:57]
  wire  _T_2346; // @[Xbar.scala 256:54]
  wire  _T_2347; // @[Xbar.scala 256:60]
  wire  _T_2348; // @[Xbar.scala 256:57]
  wire  _T_2349; // @[Xbar.scala 256:54]
  wire  _T_2350; // @[Xbar.scala 256:60]
  wire  _T_2351; // @[Xbar.scala 256:57]
  wire  _T_2352; // @[Xbar.scala 256:54]
  wire  _T_2353; // @[Xbar.scala 256:60]
  wire  _T_2354; // @[Xbar.scala 256:57]
  wire  _T_2355; // @[Xbar.scala 256:54]
  wire  _T_2356; // @[Xbar.scala 256:60]
  wire  _T_2357; // @[Xbar.scala 256:57]
  wire  _T_2358; // @[Xbar.scala 256:54]
  wire  _T_2359; // @[Xbar.scala 256:60]
  wire  _T_2360; // @[Xbar.scala 256:57]
  wire  _T_2361; // @[Xbar.scala 256:54]
  wire  _T_2362; // @[Xbar.scala 256:60]
  wire  _T_2363; // @[Xbar.scala 256:57]
  wire  _T_2364; // @[Xbar.scala 256:54]
  wire  _T_2365; // @[Xbar.scala 256:60]
  wire  _T_2366; // @[Xbar.scala 256:57]
  wire  _T_2367; // @[Xbar.scala 256:54]
  wire  _T_2368; // @[Xbar.scala 256:60]
  wire  _T_2369; // @[Xbar.scala 256:57]
  wire  _T_2370; // @[Xbar.scala 256:54]
  wire  _T_2371; // @[Xbar.scala 256:60]
  wire  _T_2372; // @[Xbar.scala 256:57]
  wire  _T_2374; // @[Xbar.scala 256:75]
  wire  _T_2375; // @[Xbar.scala 256:75]
  wire  _T_2376; // @[Xbar.scala 256:75]
  wire  _T_2377; // @[Xbar.scala 256:75]
  wire  _T_2378; // @[Xbar.scala 256:75]
  wire  _T_2379; // @[Xbar.scala 256:75]
  wire  _T_2380; // @[Xbar.scala 256:75]
  wire  _T_2381; // @[Xbar.scala 256:75]
  wire  _T_2382; // @[Xbar.scala 256:75]
  wire  _T_2383; // @[Xbar.scala 256:75]
  wire  _T_2384; // @[Xbar.scala 256:75]
  wire  _T_2385; // @[Xbar.scala 256:75]
  wire  _T_2386; // @[Xbar.scala 256:75]
  wire  _T_2387; // @[Xbar.scala 256:75]
  wire  _T_2388; // @[Xbar.scala 256:75]
  wire  _T_2389; // @[Xbar.scala 256:75]
  wire  _T_2390; // @[Xbar.scala 256:75]
  wire  _T_2391; // @[Xbar.scala 256:75]
  wire  _T_2392; // @[Xbar.scala 256:75]
  wire  _T_2393; // @[Xbar.scala 256:75]
  wire  _T_2395; // @[Xbar.scala 256:11]
  wire  _T_2396; // @[Xbar.scala 256:11]
  wire  _T_2397; // @[Xbar.scala 258:13]
  wire  _T_2419; // @[Xbar.scala 258:23]
  wire  _T_2421; // @[Xbar.scala 258:12]
  wire  _T_2422; // @[Xbar.scala 258:12]
  wire  _T_2425_0; // @[Xbar.scala 262:23]
  wire  _T_2425_1; // @[Xbar.scala 262:23]
  wire  _T_2425_2; // @[Xbar.scala 262:23]
  wire  _T_2425_3; // @[Xbar.scala 262:23]
  wire  _T_2425_4; // @[Xbar.scala 262:23]
  wire  _T_2425_5; // @[Xbar.scala 262:23]
  wire  _T_2425_6; // @[Xbar.scala 262:23]
  wire  _T_2425_7; // @[Xbar.scala 262:23]
  wire  _T_2425_8; // @[Xbar.scala 262:23]
  wire  _T_2425_9; // @[Xbar.scala 262:23]
  wire  _T_2425_10; // @[Xbar.scala 262:23]
  wire  _T_2425_11; // @[Xbar.scala 262:23]
  wire  _T_2425_12; // @[Xbar.scala 262:23]
  wire  _T_2425_13; // @[Xbar.scala 262:23]
  wire  _T_2425_14; // @[Xbar.scala 262:23]
  wire  _T_2425_15; // @[Xbar.scala 262:23]
  wire  _T_2425_16; // @[Xbar.scala 262:23]
  wire  _T_2425_17; // @[Xbar.scala 262:23]
  wire  _T_2425_18; // @[Xbar.scala 262:23]
  wire  _T_2425_19; // @[Xbar.scala 262:23]
  wire  _T_2425_20; // @[Xbar.scala 262:23]
  wire  _T_2425_21; // @[Xbar.scala 262:23]
  wire  _GEN_96; // @[Xbar.scala 266:21]
  wire  _GEN_97; // @[Xbar.scala 267:24]
  wire  _T_2427_0; // @[Xbar.scala 270:24]
  wire  _T_2427_1; // @[Xbar.scala 270:24]
  wire  _T_2427_2; // @[Xbar.scala 270:24]
  wire  _T_2427_3; // @[Xbar.scala 270:24]
  wire  _T_2427_4; // @[Xbar.scala 270:24]
  wire  _T_2427_5; // @[Xbar.scala 270:24]
  wire  _T_2427_6; // @[Xbar.scala 270:24]
  wire  _T_2427_7; // @[Xbar.scala 270:24]
  wire  _T_2427_8; // @[Xbar.scala 270:24]
  wire  _T_2427_9; // @[Xbar.scala 270:24]
  wire  _T_2427_10; // @[Xbar.scala 270:24]
  wire  _T_2427_11; // @[Xbar.scala 270:24]
  wire  _T_2427_12; // @[Xbar.scala 270:24]
  wire  _T_2427_13; // @[Xbar.scala 270:24]
  wire  _T_2427_14; // @[Xbar.scala 270:24]
  wire  _T_2427_15; // @[Xbar.scala 270:24]
  wire  _T_2427_16; // @[Xbar.scala 270:24]
  wire  _T_2427_17; // @[Xbar.scala 270:24]
  wire  _T_2427_18; // @[Xbar.scala 270:24]
  wire  _T_2427_19; // @[Xbar.scala 270:24]
  wire  _T_2427_20; // @[Xbar.scala 270:24]
  wire  _T_2427_21; // @[Xbar.scala 270:24]
  wire [2:0] _T_2495; // @[Mux.scala 27:72]
  wire [2:0] _T_2496; // @[Mux.scala 27:72]
  wire [2:0] _T_2497; // @[Mux.scala 27:72]
  wire [2:0] _T_2498; // @[Mux.scala 27:72]
  wire [2:0] _T_2499; // @[Mux.scala 27:72]
  wire [2:0] _T_2500; // @[Mux.scala 27:72]
  wire [2:0] _T_2501; // @[Mux.scala 27:72]
  wire [2:0] _T_2502; // @[Mux.scala 27:72]
  wire [2:0] _T_2503; // @[Mux.scala 27:72]
  wire [2:0] _T_2504; // @[Mux.scala 27:72]
  wire [2:0] _T_2505; // @[Mux.scala 27:72]
  wire [2:0] _T_2506; // @[Mux.scala 27:72]
  wire [2:0] _T_2507; // @[Mux.scala 27:72]
  wire [2:0] _T_2508; // @[Mux.scala 27:72]
  wire [2:0] _T_2509; // @[Mux.scala 27:72]
  wire [2:0] _T_2510; // @[Mux.scala 27:72]
  wire [2:0] _T_2511; // @[Mux.scala 27:72]
  wire [2:0] _T_2512; // @[Mux.scala 27:72]
  wire [2:0] _T_2513; // @[Mux.scala 27:72]
  wire [2:0] _T_2514; // @[Mux.scala 27:72]
  wire [2:0] _T_2515; // @[Mux.scala 27:72]
  wire [2:0] _T_2516; // @[Mux.scala 27:72]
  wire [2:0] _T_2517; // @[Mux.scala 27:72]
  wire [2:0] _T_2518; // @[Mux.scala 27:72]
  wire [2:0] _T_2519; // @[Mux.scala 27:72]
  wire [2:0] _T_2520; // @[Mux.scala 27:72]
  wire [2:0] _T_2521; // @[Mux.scala 27:72]
  wire [2:0] _T_2522; // @[Mux.scala 27:72]
  wire [2:0] _T_2523; // @[Mux.scala 27:72]
  wire [2:0] _T_2524; // @[Mux.scala 27:72]
  wire [2:0] _T_2525; // @[Mux.scala 27:72]
  wire [2:0] _T_2526; // @[Mux.scala 27:72]
  wire [2:0] _T_2527; // @[Mux.scala 27:72]
  wire [2:0] _T_2528; // @[Mux.scala 27:72]
  wire [2:0] _T_2529; // @[Mux.scala 27:72]
  wire [2:0] _T_2530; // @[Mux.scala 27:72]
  wire [2:0] _T_2531; // @[Mux.scala 27:72]
  wire [2:0] _T_2532; // @[Mux.scala 27:72]
  wire [2:0] _T_2533; // @[Mux.scala 27:72]
  wire [2:0] _T_2534; // @[Mux.scala 27:72]
  wire [2:0] _T_2535; // @[Mux.scala 27:72]
  wire [2:0] _T_2536; // @[Mux.scala 27:72]
  wire [2:0] _T_2537; // @[Mux.scala 27:72]
  wire [2:0] _T_2538; // @[Mux.scala 27:72]
  wire [2:0] _T_2539; // @[Mux.scala 27:72]
  wire [2:0] _T_2540; // @[Mux.scala 27:72]
  wire [2:0] _T_2541; // @[Mux.scala 27:72]
  wire [2:0] _T_2542; // @[Mux.scala 27:72]
  wire [2:0] _T_2543; // @[Mux.scala 27:72]
  wire [2:0] _T_2544; // @[Mux.scala 27:72]
  wire [2:0] _T_2545; // @[Mux.scala 27:72]
  wire [2:0] _T_2546; // @[Mux.scala 27:72]
  wire [2:0] _T_2547; // @[Mux.scala 27:72]
  wire [2:0] _T_2548; // @[Mux.scala 27:72]
  wire [2:0] _T_2549; // @[Mux.scala 27:72]
  wire [2:0] _T_2550; // @[Mux.scala 27:72]
  wire [2:0] _T_2551; // @[Mux.scala 27:72]
  wire [2:0] _T_2552; // @[Mux.scala 27:72]
  wire [2:0] _T_2553; // @[Mux.scala 27:72]
  wire [2:0] _T_2554; // @[Mux.scala 27:72]
  wire [2:0] _T_2555; // @[Mux.scala 27:72]
  wire [2:0] _T_2556; // @[Mux.scala 27:72]
  wire [2:0] _T_2557; // @[Mux.scala 27:72]
  wire [2:0] _T_2558; // @[Mux.scala 27:72]
  wire [2:0] _T_2559; // @[Mux.scala 27:72]
  QueueCompatibility_8 awIn_0 ( // @[Xbar.scala 55:47]
    .clock(awIn_0_clock),
    .reset(awIn_0_reset),
    .io_enq_ready(awIn_0_io_enq_ready),
    .io_enq_valid(awIn_0_io_enq_valid),
    .io_enq_bits(awIn_0_io_enq_bits),
    .io_deq_ready(awIn_0_io_deq_ready),
    .io_deq_valid(awIn_0_io_deq_valid),
    .io_deq_bits(awIn_0_io_deq_bits)
  );
  assign _T_1 = {1'b0,$signed(auto_in_ar_bits_addr)}; // @[Parameters.scala 137:49]
  assign _T_3 = $signed(_T_1) & 31'shf130; // @[Parameters.scala 137:52]
  assign requestARIO_0_0 = $signed(_T_3) == 31'sh0; // @[Parameters.scala 137:67]
  assign _T_5 = auto_in_ar_bits_addr ^ 30'h1000; // @[Parameters.scala 137:31]
  assign _T_6 = {1'b0,$signed(_T_5)}; // @[Parameters.scala 137:49]
  assign _T_8 = $signed(_T_6) & 31'shf000; // @[Parameters.scala 137:52]
  assign _T_9 = $signed(_T_8) == 31'sh0; // @[Parameters.scala 137:67]
  assign _T_10 = auto_in_ar_bits_addr ^ 30'h2100; // @[Parameters.scala 137:31]
  assign _T_11 = {1'b0,$signed(_T_10)}; // @[Parameters.scala 137:49]
  assign _T_13 = $signed(_T_11) & 31'shf100; // @[Parameters.scala 137:52]
  assign _T_14 = $signed(_T_13) == 31'sh0; // @[Parameters.scala 137:67]
  assign requestARIO_0_1 = _T_9 | _T_14; // @[Xbar.scala 52:97]
  assign _T_16 = auto_in_ar_bits_addr ^ 30'h2000; // @[Parameters.scala 137:31]
  assign _T_17 = {1'b0,$signed(_T_16)}; // @[Parameters.scala 137:49]
  assign _T_19 = $signed(_T_17) & 31'shf130; // @[Parameters.scala 137:52]
  assign requestARIO_0_2 = $signed(_T_19) == 31'sh0; // @[Parameters.scala 137:67]
  assign _T_21 = auto_in_ar_bits_addr ^ 30'h2010; // @[Parameters.scala 137:31]
  assign _T_22 = {1'b0,$signed(_T_21)}; // @[Parameters.scala 137:49]
  assign _T_24 = $signed(_T_22) & 31'shf130; // @[Parameters.scala 137:52]
  assign requestARIO_0_3 = $signed(_T_24) == 31'sh0; // @[Parameters.scala 137:67]
  assign _T_26 = auto_in_ar_bits_addr ^ 30'h2020; // @[Parameters.scala 137:31]
  assign _T_27 = {1'b0,$signed(_T_26)}; // @[Parameters.scala 137:49]
  assign _T_29 = $signed(_T_27) & 31'shf130; // @[Parameters.scala 137:52]
  assign requestARIO_0_4 = $signed(_T_29) == 31'sh0; // @[Parameters.scala 137:67]
  assign _T_31 = auto_in_ar_bits_addr ^ 30'h3000; // @[Parameters.scala 137:31]
  assign _T_32 = {1'b0,$signed(_T_31)}; // @[Parameters.scala 137:49]
  assign _T_34 = $signed(_T_32) & 31'shf130; // @[Parameters.scala 137:52]
  assign requestARIO_0_5 = $signed(_T_34) == 31'sh0; // @[Parameters.scala 137:67]
  assign _T_36 = auto_in_ar_bits_addr ^ 30'h3100; // @[Parameters.scala 137:31]
  assign _T_37 = {1'b0,$signed(_T_36)}; // @[Parameters.scala 137:49]
  assign _T_39 = $signed(_T_37) & 31'shf130; // @[Parameters.scala 137:52]
  assign requestARIO_0_6 = $signed(_T_39) == 31'sh0; // @[Parameters.scala 137:67]
  assign _T_41 = auto_in_ar_bits_addr ^ 30'h3110; // @[Parameters.scala 137:31]
  assign _T_42 = {1'b0,$signed(_T_41)}; // @[Parameters.scala 137:49]
  assign _T_44 = $signed(_T_42) & 31'shf130; // @[Parameters.scala 137:52]
  assign requestARIO_0_7 = $signed(_T_44) == 31'sh0; // @[Parameters.scala 137:67]
  assign _T_46 = auto_in_ar_bits_addr ^ 30'h3120; // @[Parameters.scala 137:31]
  assign _T_47 = {1'b0,$signed(_T_46)}; // @[Parameters.scala 137:49]
  assign _T_49 = $signed(_T_47) & 31'shf130; // @[Parameters.scala 137:52]
  assign requestARIO_0_8 = $signed(_T_49) == 31'sh0; // @[Parameters.scala 137:67]
  assign _T_51 = auto_in_ar_bits_addr ^ 30'h4000; // @[Parameters.scala 137:31]
  assign _T_52 = {1'b0,$signed(_T_51)}; // @[Parameters.scala 137:49]
  assign _T_54 = $signed(_T_52) & 31'shf100; // @[Parameters.scala 137:52]
  assign requestARIO_0_9 = $signed(_T_54) == 31'sh0; // @[Parameters.scala 137:67]
  assign _T_56 = auto_in_ar_bits_addr ^ 30'h4100; // @[Parameters.scala 137:31]
  assign _T_57 = {1'b0,$signed(_T_56)}; // @[Parameters.scala 137:49]
  assign _T_59 = $signed(_T_57) & 31'shf130; // @[Parameters.scala 137:52]
  assign requestARIO_0_10 = $signed(_T_59) == 31'sh0; // @[Parameters.scala 137:67]
  assign _T_61 = auto_in_ar_bits_addr ^ 30'h4110; // @[Parameters.scala 137:31]
  assign _T_62 = {1'b0,$signed(_T_61)}; // @[Parameters.scala 137:49]
  assign _T_64 = $signed(_T_62) & 31'shf130; // @[Parameters.scala 137:52]
  assign requestARIO_0_11 = $signed(_T_64) == 31'sh0; // @[Parameters.scala 137:67]
  assign _T_66 = auto_in_ar_bits_addr ^ 30'h4120; // @[Parameters.scala 137:31]
  assign _T_67 = {1'b0,$signed(_T_66)}; // @[Parameters.scala 137:49]
  assign _T_69 = $signed(_T_67) & 31'shf130; // @[Parameters.scala 137:52]
  assign requestARIO_0_12 = $signed(_T_69) == 31'sh0; // @[Parameters.scala 137:67]
  assign _T_71 = auto_in_ar_bits_addr ^ 30'h5000; // @[Parameters.scala 137:31]
  assign _T_72 = {1'b0,$signed(_T_71)}; // @[Parameters.scala 137:49]
  assign _T_74 = $signed(_T_72) & 31'shf100; // @[Parameters.scala 137:52]
  assign requestARIO_0_13 = $signed(_T_74) == 31'sh0; // @[Parameters.scala 137:67]
  assign _T_76 = auto_in_ar_bits_addr ^ 30'h5100; // @[Parameters.scala 137:31]
  assign _T_77 = {1'b0,$signed(_T_76)}; // @[Parameters.scala 137:49]
  assign _T_79 = $signed(_T_77) & 31'shf130; // @[Parameters.scala 137:52]
  assign requestARIO_0_14 = $signed(_T_79) == 31'sh0; // @[Parameters.scala 137:67]
  assign _T_81 = auto_in_ar_bits_addr ^ 30'h5110; // @[Parameters.scala 137:31]
  assign _T_82 = {1'b0,$signed(_T_81)}; // @[Parameters.scala 137:49]
  assign _T_84 = $signed(_T_82) & 31'shf130; // @[Parameters.scala 137:52]
  assign requestARIO_0_15 = $signed(_T_84) == 31'sh0; // @[Parameters.scala 137:67]
  assign _T_86 = auto_in_ar_bits_addr ^ 30'h5120; // @[Parameters.scala 137:31]
  assign _T_87 = {1'b0,$signed(_T_86)}; // @[Parameters.scala 137:49]
  assign _T_89 = $signed(_T_87) & 31'shf130; // @[Parameters.scala 137:52]
  assign requestARIO_0_16 = $signed(_T_89) == 31'sh0; // @[Parameters.scala 137:67]
  assign _T_91 = auto_in_ar_bits_addr ^ 30'h8000; // @[Parameters.scala 137:31]
  assign _T_92 = {1'b0,$signed(_T_91)}; // @[Parameters.scala 137:49]
  assign _T_94 = $signed(_T_92) & 31'shf130; // @[Parameters.scala 137:52]
  assign requestARIO_0_17 = $signed(_T_94) == 31'sh0; // @[Parameters.scala 137:67]
  assign _T_96 = auto_in_ar_bits_addr ^ 30'h8010; // @[Parameters.scala 137:31]
  assign _T_97 = {1'b0,$signed(_T_96)}; // @[Parameters.scala 137:49]
  assign _T_99 = $signed(_T_97) & 31'shf130; // @[Parameters.scala 137:52]
  assign requestARIO_0_18 = $signed(_T_99) == 31'sh0; // @[Parameters.scala 137:67]
  assign _T_101 = auto_in_ar_bits_addr ^ 30'h9000; // @[Parameters.scala 137:31]
  assign _T_102 = {1'b0,$signed(_T_101)}; // @[Parameters.scala 137:49]
  assign _T_104 = $signed(_T_102) & 31'shf100; // @[Parameters.scala 137:52]
  assign requestARIO_0_19 = $signed(_T_104) == 31'sh0; // @[Parameters.scala 137:67]
  assign _T_106 = auto_in_ar_bits_addr ^ 30'h9100; // @[Parameters.scala 137:31]
  assign _T_107 = {1'b0,$signed(_T_106)}; // @[Parameters.scala 137:49]
  assign _T_109 = $signed(_T_107) & 31'shf130; // @[Parameters.scala 137:52]
  assign requestARIO_0_20 = $signed(_T_109) == 31'sh0; // @[Parameters.scala 137:67]
  assign _T_111 = auto_in_ar_bits_addr ^ 30'h6000; // @[Parameters.scala 137:31]
  assign _T_112 = {1'b0,$signed(_T_111)}; // @[Parameters.scala 137:49]
  assign _T_114 = $signed(_T_112) & 31'shf000; // @[Parameters.scala 137:52]
  assign _T_115 = $signed(_T_114) == 31'sh0; // @[Parameters.scala 137:67]
  assign _T_116 = auto_in_ar_bits_addr ^ 30'h7000; // @[Parameters.scala 137:31]
  assign _T_117 = {1'b0,$signed(_T_116)}; // @[Parameters.scala 137:49]
  assign _T_119 = $signed(_T_117) & 31'shf130; // @[Parameters.scala 137:52]
  assign _T_120 = $signed(_T_119) == 31'sh0; // @[Parameters.scala 137:67]
  assign requestARIO_0_21 = _T_115 | _T_120; // @[Xbar.scala 52:97]
  assign _T_123 = {1'b0,$signed(auto_in_aw_bits_addr)}; // @[Parameters.scala 137:49]
  assign _T_125 = $signed(_T_123) & 31'shf130; // @[Parameters.scala 137:52]
  assign requestAWIO_0_0 = $signed(_T_125) == 31'sh0; // @[Parameters.scala 137:67]
  assign _T_127 = auto_in_aw_bits_addr ^ 30'h1000; // @[Parameters.scala 137:31]
  assign _T_128 = {1'b0,$signed(_T_127)}; // @[Parameters.scala 137:49]
  assign _T_130 = $signed(_T_128) & 31'shf000; // @[Parameters.scala 137:52]
  assign _T_131 = $signed(_T_130) == 31'sh0; // @[Parameters.scala 137:67]
  assign _T_132 = auto_in_aw_bits_addr ^ 30'h2100; // @[Parameters.scala 137:31]
  assign _T_133 = {1'b0,$signed(_T_132)}; // @[Parameters.scala 137:49]
  assign _T_135 = $signed(_T_133) & 31'shf100; // @[Parameters.scala 137:52]
  assign _T_136 = $signed(_T_135) == 31'sh0; // @[Parameters.scala 137:67]
  assign requestAWIO_0_1 = _T_131 | _T_136; // @[Xbar.scala 52:97]
  assign _T_138 = auto_in_aw_bits_addr ^ 30'h2000; // @[Parameters.scala 137:31]
  assign _T_139 = {1'b0,$signed(_T_138)}; // @[Parameters.scala 137:49]
  assign _T_141 = $signed(_T_139) & 31'shf130; // @[Parameters.scala 137:52]
  assign requestAWIO_0_2 = $signed(_T_141) == 31'sh0; // @[Parameters.scala 137:67]
  assign _T_143 = auto_in_aw_bits_addr ^ 30'h2010; // @[Parameters.scala 137:31]
  assign _T_144 = {1'b0,$signed(_T_143)}; // @[Parameters.scala 137:49]
  assign _T_146 = $signed(_T_144) & 31'shf130; // @[Parameters.scala 137:52]
  assign requestAWIO_0_3 = $signed(_T_146) == 31'sh0; // @[Parameters.scala 137:67]
  assign _T_148 = auto_in_aw_bits_addr ^ 30'h2020; // @[Parameters.scala 137:31]
  assign _T_149 = {1'b0,$signed(_T_148)}; // @[Parameters.scala 137:49]
  assign _T_151 = $signed(_T_149) & 31'shf130; // @[Parameters.scala 137:52]
  assign requestAWIO_0_4 = $signed(_T_151) == 31'sh0; // @[Parameters.scala 137:67]
  assign _T_153 = auto_in_aw_bits_addr ^ 30'h3000; // @[Parameters.scala 137:31]
  assign _T_154 = {1'b0,$signed(_T_153)}; // @[Parameters.scala 137:49]
  assign _T_156 = $signed(_T_154) & 31'shf130; // @[Parameters.scala 137:52]
  assign requestAWIO_0_5 = $signed(_T_156) == 31'sh0; // @[Parameters.scala 137:67]
  assign _T_158 = auto_in_aw_bits_addr ^ 30'h3100; // @[Parameters.scala 137:31]
  assign _T_159 = {1'b0,$signed(_T_158)}; // @[Parameters.scala 137:49]
  assign _T_161 = $signed(_T_159) & 31'shf130; // @[Parameters.scala 137:52]
  assign requestAWIO_0_6 = $signed(_T_161) == 31'sh0; // @[Parameters.scala 137:67]
  assign _T_163 = auto_in_aw_bits_addr ^ 30'h3110; // @[Parameters.scala 137:31]
  assign _T_164 = {1'b0,$signed(_T_163)}; // @[Parameters.scala 137:49]
  assign _T_166 = $signed(_T_164) & 31'shf130; // @[Parameters.scala 137:52]
  assign requestAWIO_0_7 = $signed(_T_166) == 31'sh0; // @[Parameters.scala 137:67]
  assign _T_168 = auto_in_aw_bits_addr ^ 30'h3120; // @[Parameters.scala 137:31]
  assign _T_169 = {1'b0,$signed(_T_168)}; // @[Parameters.scala 137:49]
  assign _T_171 = $signed(_T_169) & 31'shf130; // @[Parameters.scala 137:52]
  assign requestAWIO_0_8 = $signed(_T_171) == 31'sh0; // @[Parameters.scala 137:67]
  assign _T_173 = auto_in_aw_bits_addr ^ 30'h4000; // @[Parameters.scala 137:31]
  assign _T_174 = {1'b0,$signed(_T_173)}; // @[Parameters.scala 137:49]
  assign _T_176 = $signed(_T_174) & 31'shf100; // @[Parameters.scala 137:52]
  assign requestAWIO_0_9 = $signed(_T_176) == 31'sh0; // @[Parameters.scala 137:67]
  assign _T_178 = auto_in_aw_bits_addr ^ 30'h4100; // @[Parameters.scala 137:31]
  assign _T_179 = {1'b0,$signed(_T_178)}; // @[Parameters.scala 137:49]
  assign _T_181 = $signed(_T_179) & 31'shf130; // @[Parameters.scala 137:52]
  assign requestAWIO_0_10 = $signed(_T_181) == 31'sh0; // @[Parameters.scala 137:67]
  assign _T_183 = auto_in_aw_bits_addr ^ 30'h4110; // @[Parameters.scala 137:31]
  assign _T_184 = {1'b0,$signed(_T_183)}; // @[Parameters.scala 137:49]
  assign _T_186 = $signed(_T_184) & 31'shf130; // @[Parameters.scala 137:52]
  assign requestAWIO_0_11 = $signed(_T_186) == 31'sh0; // @[Parameters.scala 137:67]
  assign _T_188 = auto_in_aw_bits_addr ^ 30'h4120; // @[Parameters.scala 137:31]
  assign _T_189 = {1'b0,$signed(_T_188)}; // @[Parameters.scala 137:49]
  assign _T_191 = $signed(_T_189) & 31'shf130; // @[Parameters.scala 137:52]
  assign requestAWIO_0_12 = $signed(_T_191) == 31'sh0; // @[Parameters.scala 137:67]
  assign _T_193 = auto_in_aw_bits_addr ^ 30'h5000; // @[Parameters.scala 137:31]
  assign _T_194 = {1'b0,$signed(_T_193)}; // @[Parameters.scala 137:49]
  assign _T_196 = $signed(_T_194) & 31'shf100; // @[Parameters.scala 137:52]
  assign requestAWIO_0_13 = $signed(_T_196) == 31'sh0; // @[Parameters.scala 137:67]
  assign _T_198 = auto_in_aw_bits_addr ^ 30'h5100; // @[Parameters.scala 137:31]
  assign _T_199 = {1'b0,$signed(_T_198)}; // @[Parameters.scala 137:49]
  assign _T_201 = $signed(_T_199) & 31'shf130; // @[Parameters.scala 137:52]
  assign requestAWIO_0_14 = $signed(_T_201) == 31'sh0; // @[Parameters.scala 137:67]
  assign _T_203 = auto_in_aw_bits_addr ^ 30'h5110; // @[Parameters.scala 137:31]
  assign _T_204 = {1'b0,$signed(_T_203)}; // @[Parameters.scala 137:49]
  assign _T_206 = $signed(_T_204) & 31'shf130; // @[Parameters.scala 137:52]
  assign requestAWIO_0_15 = $signed(_T_206) == 31'sh0; // @[Parameters.scala 137:67]
  assign _T_208 = auto_in_aw_bits_addr ^ 30'h5120; // @[Parameters.scala 137:31]
  assign _T_209 = {1'b0,$signed(_T_208)}; // @[Parameters.scala 137:49]
  assign _T_211 = $signed(_T_209) & 31'shf130; // @[Parameters.scala 137:52]
  assign requestAWIO_0_16 = $signed(_T_211) == 31'sh0; // @[Parameters.scala 137:67]
  assign _T_213 = auto_in_aw_bits_addr ^ 30'h8000; // @[Parameters.scala 137:31]
  assign _T_214 = {1'b0,$signed(_T_213)}; // @[Parameters.scala 137:49]
  assign _T_216 = $signed(_T_214) & 31'shf130; // @[Parameters.scala 137:52]
  assign requestAWIO_0_17 = $signed(_T_216) == 31'sh0; // @[Parameters.scala 137:67]
  assign _T_218 = auto_in_aw_bits_addr ^ 30'h8010; // @[Parameters.scala 137:31]
  assign _T_219 = {1'b0,$signed(_T_218)}; // @[Parameters.scala 137:49]
  assign _T_221 = $signed(_T_219) & 31'shf130; // @[Parameters.scala 137:52]
  assign requestAWIO_0_18 = $signed(_T_221) == 31'sh0; // @[Parameters.scala 137:67]
  assign _T_223 = auto_in_aw_bits_addr ^ 30'h9000; // @[Parameters.scala 137:31]
  assign _T_224 = {1'b0,$signed(_T_223)}; // @[Parameters.scala 137:49]
  assign _T_226 = $signed(_T_224) & 31'shf100; // @[Parameters.scala 137:52]
  assign requestAWIO_0_19 = $signed(_T_226) == 31'sh0; // @[Parameters.scala 137:67]
  assign _T_228 = auto_in_aw_bits_addr ^ 30'h9100; // @[Parameters.scala 137:31]
  assign _T_229 = {1'b0,$signed(_T_228)}; // @[Parameters.scala 137:49]
  assign _T_231 = $signed(_T_229) & 31'shf130; // @[Parameters.scala 137:52]
  assign requestAWIO_0_20 = $signed(_T_231) == 31'sh0; // @[Parameters.scala 137:67]
  assign _T_233 = auto_in_aw_bits_addr ^ 30'h6000; // @[Parameters.scala 137:31]
  assign _T_234 = {1'b0,$signed(_T_233)}; // @[Parameters.scala 137:49]
  assign _T_236 = $signed(_T_234) & 31'shf000; // @[Parameters.scala 137:52]
  assign _T_237 = $signed(_T_236) == 31'sh0; // @[Parameters.scala 137:67]
  assign _T_238 = auto_in_aw_bits_addr ^ 30'h7000; // @[Parameters.scala 137:31]
  assign _T_239 = {1'b0,$signed(_T_238)}; // @[Parameters.scala 137:49]
  assign _T_241 = $signed(_T_239) & 31'shf130; // @[Parameters.scala 137:52]
  assign _T_242 = $signed(_T_241) == 31'sh0; // @[Parameters.scala 137:67]
  assign requestAWIO_0_21 = _T_237 | _T_242; // @[Xbar.scala 52:97]
  assign requestROI_0_0 = ~auto_out_0_r_bits_id; // @[Parameters.scala 47:9]
  assign requestROI_1_0 = ~auto_out_1_r_bits_id; // @[Parameters.scala 47:9]
  assign requestROI_2_0 = ~auto_out_2_r_bits_id; // @[Parameters.scala 47:9]
  assign requestROI_3_0 = ~auto_out_3_r_bits_id; // @[Parameters.scala 47:9]
  assign requestROI_4_0 = ~auto_out_4_r_bits_id; // @[Parameters.scala 47:9]
  assign requestROI_5_0 = ~auto_out_5_r_bits_id; // @[Parameters.scala 47:9]
  assign requestROI_6_0 = ~auto_out_6_r_bits_id; // @[Parameters.scala 47:9]
  assign requestROI_7_0 = ~auto_out_7_r_bits_id; // @[Parameters.scala 47:9]
  assign requestROI_8_0 = ~auto_out_8_r_bits_id; // @[Parameters.scala 47:9]
  assign requestROI_9_0 = ~auto_out_9_r_bits_id; // @[Parameters.scala 47:9]
  assign requestROI_10_0 = ~auto_out_10_r_bits_id; // @[Parameters.scala 47:9]
  assign requestROI_11_0 = ~auto_out_11_r_bits_id; // @[Parameters.scala 47:9]
  assign requestROI_12_0 = ~auto_out_12_r_bits_id; // @[Parameters.scala 47:9]
  assign requestROI_13_0 = ~auto_out_13_r_bits_id; // @[Parameters.scala 47:9]
  assign requestROI_14_0 = ~auto_out_14_r_bits_id; // @[Parameters.scala 47:9]
  assign requestROI_15_0 = ~auto_out_15_r_bits_id; // @[Parameters.scala 47:9]
  assign requestROI_16_0 = ~auto_out_16_r_bits_id; // @[Parameters.scala 47:9]
  assign requestROI_17_0 = ~auto_out_17_r_bits_id; // @[Parameters.scala 47:9]
  assign requestROI_18_0 = ~auto_out_18_r_bits_id; // @[Parameters.scala 47:9]
  assign requestROI_19_0 = ~auto_out_19_r_bits_id; // @[Parameters.scala 47:9]
  assign requestROI_20_0 = ~auto_out_20_r_bits_id; // @[Parameters.scala 47:9]
  assign requestBOI_0_0 = ~auto_out_0_b_bits_id; // @[Parameters.scala 47:9]
  assign requestBOI_1_0 = ~auto_out_1_b_bits_id; // @[Parameters.scala 47:9]
  assign requestBOI_2_0 = ~auto_out_2_b_bits_id; // @[Parameters.scala 47:9]
  assign requestBOI_3_0 = ~auto_out_3_b_bits_id; // @[Parameters.scala 47:9]
  assign requestBOI_4_0 = ~auto_out_4_b_bits_id; // @[Parameters.scala 47:9]
  assign requestBOI_5_0 = ~auto_out_5_b_bits_id; // @[Parameters.scala 47:9]
  assign requestBOI_6_0 = ~auto_out_6_b_bits_id; // @[Parameters.scala 47:9]
  assign requestBOI_7_0 = ~auto_out_7_b_bits_id; // @[Parameters.scala 47:9]
  assign requestBOI_8_0 = ~auto_out_8_b_bits_id; // @[Parameters.scala 47:9]
  assign requestBOI_9_0 = ~auto_out_9_b_bits_id; // @[Parameters.scala 47:9]
  assign requestBOI_10_0 = ~auto_out_10_b_bits_id; // @[Parameters.scala 47:9]
  assign requestBOI_11_0 = ~auto_out_11_b_bits_id; // @[Parameters.scala 47:9]
  assign requestBOI_12_0 = ~auto_out_12_b_bits_id; // @[Parameters.scala 47:9]
  assign requestBOI_13_0 = ~auto_out_13_b_bits_id; // @[Parameters.scala 47:9]
  assign requestBOI_14_0 = ~auto_out_14_b_bits_id; // @[Parameters.scala 47:9]
  assign requestBOI_15_0 = ~auto_out_15_b_bits_id; // @[Parameters.scala 47:9]
  assign requestBOI_16_0 = ~auto_out_16_b_bits_id; // @[Parameters.scala 47:9]
  assign requestBOI_17_0 = ~auto_out_17_b_bits_id; // @[Parameters.scala 47:9]
  assign requestBOI_18_0 = ~auto_out_18_b_bits_id; // @[Parameters.scala 47:9]
  assign requestBOI_19_0 = ~auto_out_19_b_bits_id; // @[Parameters.scala 47:9]
  assign requestBOI_20_0 = ~auto_out_20_b_bits_id; // @[Parameters.scala 47:9]
  assign _T_247 = {requestAWIO_0_4,requestAWIO_0_3,requestAWIO_0_2,requestAWIO_0_1,requestAWIO_0_0}; // @[Xbar.scala 64:75]
  assign _T_253 = {requestAWIO_0_10,requestAWIO_0_9,requestAWIO_0_8,requestAWIO_0_7,requestAWIO_0_6,requestAWIO_0_5,_T_247}; // @[Xbar.scala 64:75]
  assign _T_257 = {requestAWIO_0_15,requestAWIO_0_14,requestAWIO_0_13,requestAWIO_0_12,requestAWIO_0_11}; // @[Xbar.scala 64:75]
  assign _T_263 = {requestAWIO_0_21,requestAWIO_0_20,requestAWIO_0_19,requestAWIO_0_18,requestAWIO_0_17,requestAWIO_0_16,_T_257}; // @[Xbar.scala 64:75]
  assign _T_264 = {requestAWIO_0_21,requestAWIO_0_20,requestAWIO_0_19,requestAWIO_0_18,requestAWIO_0_17,requestAWIO_0_16,_T_257,_T_253}; // @[Xbar.scala 64:75]
  assign requestWIO_0_0 = awIn_0_io_deq_bits[0]; // @[Xbar.scala 65:73]
  assign requestWIO_0_1 = awIn_0_io_deq_bits[1]; // @[Xbar.scala 65:73]
  assign requestWIO_0_2 = awIn_0_io_deq_bits[2]; // @[Xbar.scala 65:73]
  assign requestWIO_0_3 = awIn_0_io_deq_bits[3]; // @[Xbar.scala 65:73]
  assign requestWIO_0_4 = awIn_0_io_deq_bits[4]; // @[Xbar.scala 65:73]
  assign requestWIO_0_5 = awIn_0_io_deq_bits[5]; // @[Xbar.scala 65:73]
  assign requestWIO_0_6 = awIn_0_io_deq_bits[6]; // @[Xbar.scala 65:73]
  assign requestWIO_0_7 = awIn_0_io_deq_bits[7]; // @[Xbar.scala 65:73]
  assign requestWIO_0_8 = awIn_0_io_deq_bits[8]; // @[Xbar.scala 65:73]
  assign requestWIO_0_9 = awIn_0_io_deq_bits[9]; // @[Xbar.scala 65:73]
  assign requestWIO_0_10 = awIn_0_io_deq_bits[10]; // @[Xbar.scala 65:73]
  assign requestWIO_0_11 = awIn_0_io_deq_bits[11]; // @[Xbar.scala 65:73]
  assign requestWIO_0_12 = awIn_0_io_deq_bits[12]; // @[Xbar.scala 65:73]
  assign requestWIO_0_13 = awIn_0_io_deq_bits[13]; // @[Xbar.scala 65:73]
  assign requestWIO_0_14 = awIn_0_io_deq_bits[14]; // @[Xbar.scala 65:73]
  assign requestWIO_0_15 = awIn_0_io_deq_bits[15]; // @[Xbar.scala 65:73]
  assign requestWIO_0_16 = awIn_0_io_deq_bits[16]; // @[Xbar.scala 65:73]
  assign requestWIO_0_17 = awIn_0_io_deq_bits[17]; // @[Xbar.scala 65:73]
  assign requestWIO_0_18 = awIn_0_io_deq_bits[18]; // @[Xbar.scala 65:73]
  assign requestWIO_0_19 = awIn_0_io_deq_bits[19]; // @[Xbar.scala 65:73]
  assign requestWIO_0_20 = awIn_0_io_deq_bits[20]; // @[Xbar.scala 65:73]
  assign requestWIO_0_21 = awIn_0_io_deq_bits[21]; // @[Xbar.scala 65:73]
  assign _T_274 = {requestARIO_0_4,requestARIO_0_3,requestARIO_0_2,requestARIO_0_1,requestARIO_0_0}; // @[Xbar.scala 93:45]
  assign _T_280 = {requestARIO_0_10,requestARIO_0_9,requestARIO_0_8,requestARIO_0_7,requestARIO_0_6,requestARIO_0_5,_T_274}; // @[Xbar.scala 93:45]
  assign _T_284 = {requestARIO_0_15,requestARIO_0_14,requestARIO_0_13,requestARIO_0_12,requestARIO_0_11}; // @[Xbar.scala 93:45]
  assign _T_291 = {requestARIO_0_21,requestARIO_0_20,requestARIO_0_19,requestARIO_0_18,requestARIO_0_17,requestARIO_0_16,_T_284,_T_280}; // @[Xbar.scala 93:45]
  assign _T_294 = _T_291[21:16] != 6'h0; // @[OneHot.scala 32:14]
  assign _GEN_98 = {{10'd0}, _T_291[21:16]}; // @[OneHot.scala 32:28]
  assign _T_295 = _GEN_98 | _T_291[15:0]; // @[OneHot.scala 32:28]
  assign _T_298 = _T_295[15:8] != 8'h0; // @[OneHot.scala 32:14]
  assign _T_299 = _T_295[15:8] | _T_295[7:0]; // @[OneHot.scala 32:28]
  assign _T_302 = _T_299[7:4] != 4'h0; // @[OneHot.scala 32:14]
  assign _T_303 = _T_299[7:4] | _T_299[3:0]; // @[OneHot.scala 32:28]
  assign _T_306 = _T_303[3:2] != 2'h0; // @[OneHot.scala 32:14]
  assign _T_307 = _T_303[3:2] | _T_303[1:0]; // @[OneHot.scala 32:28]
  assign _T_312 = {_T_294,_T_298,_T_302,_T_306,_T_307[1]}; // @[Cat.scala 29:58]
  assign _T_336 = _T_264[21:16] != 6'h0; // @[OneHot.scala 32:14]
  assign _GEN_99 = {{10'd0}, _T_264[21:16]}; // @[OneHot.scala 32:28]
  assign _T_337 = _GEN_99 | _T_264[15:0]; // @[OneHot.scala 32:28]
  assign _T_340 = _T_337[15:8] != 8'h0; // @[OneHot.scala 32:14]
  assign _T_341 = _T_337[15:8] | _T_337[7:0]; // @[OneHot.scala 32:28]
  assign _T_344 = _T_341[7:4] != 4'h0; // @[OneHot.scala 32:14]
  assign _T_345 = _T_341[7:4] | _T_341[3:0]; // @[OneHot.scala 32:28]
  assign _T_348 = _T_345[3:2] != 2'h0; // @[OneHot.scala 32:14]
  assign _T_349 = _T_345[3:2] | _T_345[1:0]; // @[OneHot.scala 32:28]
  assign _T_354 = {_T_336,_T_340,_T_344,_T_348,_T_349[1]}; // @[Cat.scala 29:58]
  assign _T_452 = requestARIO_0_0 & auto_out_0_ar_ready; // @[Mux.scala 27:72]
  assign _T_453 = requestARIO_0_1 & auto_out_1_ar_ready; // @[Mux.scala 27:72]
  assign _T_474 = _T_452 | _T_453; // @[Mux.scala 27:72]
  assign _T_454 = requestARIO_0_2 & auto_out_2_ar_ready; // @[Mux.scala 27:72]
  assign _T_475 = _T_474 | _T_454; // @[Mux.scala 27:72]
  assign _T_455 = requestARIO_0_3 & auto_out_3_ar_ready; // @[Mux.scala 27:72]
  assign _T_476 = _T_475 | _T_455; // @[Mux.scala 27:72]
  assign _T_456 = requestARIO_0_4 & auto_out_4_ar_ready; // @[Mux.scala 27:72]
  assign _T_477 = _T_476 | _T_456; // @[Mux.scala 27:72]
  assign _T_457 = requestARIO_0_5 & auto_out_5_ar_ready; // @[Mux.scala 27:72]
  assign _T_478 = _T_477 | _T_457; // @[Mux.scala 27:72]
  assign _T_458 = requestARIO_0_6 & auto_out_6_ar_ready; // @[Mux.scala 27:72]
  assign _T_479 = _T_478 | _T_458; // @[Mux.scala 27:72]
  assign _T_459 = requestARIO_0_7 & auto_out_7_ar_ready; // @[Mux.scala 27:72]
  assign _T_480 = _T_479 | _T_459; // @[Mux.scala 27:72]
  assign _T_460 = requestARIO_0_8 & auto_out_8_ar_ready; // @[Mux.scala 27:72]
  assign _T_481 = _T_480 | _T_460; // @[Mux.scala 27:72]
  assign _T_461 = requestARIO_0_9 & auto_out_9_ar_ready; // @[Mux.scala 27:72]
  assign _T_482 = _T_481 | _T_461; // @[Mux.scala 27:72]
  assign _T_462 = requestARIO_0_10 & auto_out_10_ar_ready; // @[Mux.scala 27:72]
  assign _T_483 = _T_482 | _T_462; // @[Mux.scala 27:72]
  assign _T_463 = requestARIO_0_11 & auto_out_11_ar_ready; // @[Mux.scala 27:72]
  assign _T_484 = _T_483 | _T_463; // @[Mux.scala 27:72]
  assign _T_464 = requestARIO_0_12 & auto_out_12_ar_ready; // @[Mux.scala 27:72]
  assign _T_485 = _T_484 | _T_464; // @[Mux.scala 27:72]
  assign _T_465 = requestARIO_0_13 & auto_out_13_ar_ready; // @[Mux.scala 27:72]
  assign _T_486 = _T_485 | _T_465; // @[Mux.scala 27:72]
  assign _T_466 = requestARIO_0_14 & auto_out_14_ar_ready; // @[Mux.scala 27:72]
  assign _T_487 = _T_486 | _T_466; // @[Mux.scala 27:72]
  assign _T_467 = requestARIO_0_15 & auto_out_15_ar_ready; // @[Mux.scala 27:72]
  assign _T_488 = _T_487 | _T_467; // @[Mux.scala 27:72]
  assign _T_468 = requestARIO_0_16 & auto_out_16_ar_ready; // @[Mux.scala 27:72]
  assign _T_489 = _T_488 | _T_468; // @[Mux.scala 27:72]
  assign _T_469 = requestARIO_0_17 & auto_out_17_ar_ready; // @[Mux.scala 27:72]
  assign _T_490 = _T_489 | _T_469; // @[Mux.scala 27:72]
  assign _T_470 = requestARIO_0_18 & auto_out_18_ar_ready; // @[Mux.scala 27:72]
  assign _T_491 = _T_490 | _T_470; // @[Mux.scala 27:72]
  assign _T_471 = requestARIO_0_19 & auto_out_19_ar_ready; // @[Mux.scala 27:72]
  assign _T_492 = _T_491 | _T_471; // @[Mux.scala 27:72]
  assign _T_472 = requestARIO_0_20 & auto_out_20_ar_ready; // @[Mux.scala 27:72]
  assign _T_493 = _T_492 | _T_472; // @[Mux.scala 27:72]
  assign _T_473 = requestARIO_0_21 & auto_out_21_ar_ready; // @[Mux.scala 27:72]
  assign in_0_ar_ready = _T_493 | _T_473; // @[Mux.scala 27:72]
  assign _T_379 = _T_360 == 3'h0; // @[Xbar.scala 112:22]
  assign _T_378 = _T_361 == _T_312; // @[Xbar.scala 111:75]
  assign _T_380 = _T_379 | _T_378; // @[Xbar.scala 112:34]
  assign _T_381 = _T_360 != 3'h7; // @[Xbar.scala 112:80]
  assign _T_383 = _T_380 & _T_381; // @[Xbar.scala 112:48]
  assign io_in_0_ar_ready = in_0_ar_ready & _T_383; // @[Xbar.scala 130:45]
  assign _T_355 = io_in_0_ar_ready & auto_in_ar_valid; // @[Decoupled.scala 40:37]
  assign _T_631 = auto_out_0_r_valid & requestROI_0_0; // @[Xbar.scala 222:40]
  assign _T_633 = auto_out_1_r_valid & requestROI_1_0; // @[Xbar.scala 222:40]
  assign _T_1687 = _T_631 | _T_633; // @[Xbar.scala 246:36]
  assign _T_635 = auto_out_2_r_valid & requestROI_2_0; // @[Xbar.scala 222:40]
  assign _T_1688 = _T_1687 | _T_635; // @[Xbar.scala 246:36]
  assign _T_637 = auto_out_3_r_valid & requestROI_3_0; // @[Xbar.scala 222:40]
  assign _T_1689 = _T_1688 | _T_637; // @[Xbar.scala 246:36]
  assign _T_639 = auto_out_4_r_valid & requestROI_4_0; // @[Xbar.scala 222:40]
  assign _T_1690 = _T_1689 | _T_639; // @[Xbar.scala 246:36]
  assign _T_641 = auto_out_5_r_valid & requestROI_5_0; // @[Xbar.scala 222:40]
  assign _T_1691 = _T_1690 | _T_641; // @[Xbar.scala 246:36]
  assign _T_643 = auto_out_6_r_valid & requestROI_6_0; // @[Xbar.scala 222:40]
  assign _T_1692 = _T_1691 | _T_643; // @[Xbar.scala 246:36]
  assign _T_645 = auto_out_7_r_valid & requestROI_7_0; // @[Xbar.scala 222:40]
  assign _T_1693 = _T_1692 | _T_645; // @[Xbar.scala 246:36]
  assign _T_647 = auto_out_8_r_valid & requestROI_8_0; // @[Xbar.scala 222:40]
  assign _T_1694 = _T_1693 | _T_647; // @[Xbar.scala 246:36]
  assign _T_649 = auto_out_9_r_valid & requestROI_9_0; // @[Xbar.scala 222:40]
  assign _T_1695 = _T_1694 | _T_649; // @[Xbar.scala 246:36]
  assign _T_651 = auto_out_10_r_valid & requestROI_10_0; // @[Xbar.scala 222:40]
  assign _T_1696 = _T_1695 | _T_651; // @[Xbar.scala 246:36]
  assign _T_653 = auto_out_11_r_valid & requestROI_11_0; // @[Xbar.scala 222:40]
  assign _T_1697 = _T_1696 | _T_653; // @[Xbar.scala 246:36]
  assign _T_655 = auto_out_12_r_valid & requestROI_12_0; // @[Xbar.scala 222:40]
  assign _T_1698 = _T_1697 | _T_655; // @[Xbar.scala 246:36]
  assign _T_657 = auto_out_13_r_valid & requestROI_13_0; // @[Xbar.scala 222:40]
  assign _T_1699 = _T_1698 | _T_657; // @[Xbar.scala 246:36]
  assign _T_659 = auto_out_14_r_valid & requestROI_14_0; // @[Xbar.scala 222:40]
  assign _T_1700 = _T_1699 | _T_659; // @[Xbar.scala 246:36]
  assign _T_661 = auto_out_15_r_valid & requestROI_15_0; // @[Xbar.scala 222:40]
  assign _T_1701 = _T_1700 | _T_661; // @[Xbar.scala 246:36]
  assign _T_663 = auto_out_16_r_valid & requestROI_16_0; // @[Xbar.scala 222:40]
  assign _T_1702 = _T_1701 | _T_663; // @[Xbar.scala 246:36]
  assign _T_665 = auto_out_17_r_valid & requestROI_17_0; // @[Xbar.scala 222:40]
  assign _T_1703 = _T_1702 | _T_665; // @[Xbar.scala 246:36]
  assign _T_667 = auto_out_18_r_valid & requestROI_18_0; // @[Xbar.scala 222:40]
  assign _T_1704 = _T_1703 | _T_667; // @[Xbar.scala 246:36]
  assign _T_669 = auto_out_19_r_valid & requestROI_19_0; // @[Xbar.scala 222:40]
  assign _T_1705 = _T_1704 | _T_669; // @[Xbar.scala 246:36]
  assign _T_671 = auto_out_20_r_valid & requestROI_20_0; // @[Xbar.scala 222:40]
  assign _T_1706 = _T_1705 | _T_671; // @[Xbar.scala 246:36]
  assign _T_1707 = _T_1706 | auto_out_21_r_valid; // @[Xbar.scala 246:36]
  assign _T_1988 = _T_1962_0 & _T_631; // @[Mux.scala 27:72]
  assign _T_1989 = _T_1962_1 & _T_633; // @[Mux.scala 27:72]
  assign _T_2010 = _T_1988 | _T_1989; // @[Mux.scala 27:72]
  assign _T_1990 = _T_1962_2 & _T_635; // @[Mux.scala 27:72]
  assign _T_2011 = _T_2010 | _T_1990; // @[Mux.scala 27:72]
  assign _T_1991 = _T_1962_3 & _T_637; // @[Mux.scala 27:72]
  assign _T_2012 = _T_2011 | _T_1991; // @[Mux.scala 27:72]
  assign _T_1992 = _T_1962_4 & _T_639; // @[Mux.scala 27:72]
  assign _T_2013 = _T_2012 | _T_1992; // @[Mux.scala 27:72]
  assign _T_1993 = _T_1962_5 & _T_641; // @[Mux.scala 27:72]
  assign _T_2014 = _T_2013 | _T_1993; // @[Mux.scala 27:72]
  assign _T_1994 = _T_1962_6 & _T_643; // @[Mux.scala 27:72]
  assign _T_2015 = _T_2014 | _T_1994; // @[Mux.scala 27:72]
  assign _T_1995 = _T_1962_7 & _T_645; // @[Mux.scala 27:72]
  assign _T_2016 = _T_2015 | _T_1995; // @[Mux.scala 27:72]
  assign _T_1996 = _T_1962_8 & _T_647; // @[Mux.scala 27:72]
  assign _T_2017 = _T_2016 | _T_1996; // @[Mux.scala 27:72]
  assign _T_1997 = _T_1962_9 & _T_649; // @[Mux.scala 27:72]
  assign _T_2018 = _T_2017 | _T_1997; // @[Mux.scala 27:72]
  assign _T_1998 = _T_1962_10 & _T_651; // @[Mux.scala 27:72]
  assign _T_2019 = _T_2018 | _T_1998; // @[Mux.scala 27:72]
  assign _T_1999 = _T_1962_11 & _T_653; // @[Mux.scala 27:72]
  assign _T_2020 = _T_2019 | _T_1999; // @[Mux.scala 27:72]
  assign _T_2000 = _T_1962_12 & _T_655; // @[Mux.scala 27:72]
  assign _T_2021 = _T_2020 | _T_2000; // @[Mux.scala 27:72]
  assign _T_2001 = _T_1962_13 & _T_657; // @[Mux.scala 27:72]
  assign _T_2022 = _T_2021 | _T_2001; // @[Mux.scala 27:72]
  assign _T_2002 = _T_1962_14 & _T_659; // @[Mux.scala 27:72]
  assign _T_2023 = _T_2022 | _T_2002; // @[Mux.scala 27:72]
  assign _T_2003 = _T_1962_15 & _T_661; // @[Mux.scala 27:72]
  assign _T_2024 = _T_2023 | _T_2003; // @[Mux.scala 27:72]
  assign _T_2004 = _T_1962_16 & _T_663; // @[Mux.scala 27:72]
  assign _T_2025 = _T_2024 | _T_2004; // @[Mux.scala 27:72]
  assign _T_2005 = _T_1962_17 & _T_665; // @[Mux.scala 27:72]
  assign _T_2026 = _T_2025 | _T_2005; // @[Mux.scala 27:72]
  assign _T_2006 = _T_1962_18 & _T_667; // @[Mux.scala 27:72]
  assign _T_2027 = _T_2026 | _T_2006; // @[Mux.scala 27:72]
  assign _T_2007 = _T_1962_19 & _T_669; // @[Mux.scala 27:72]
  assign _T_2028 = _T_2027 | _T_2007; // @[Mux.scala 27:72]
  assign _T_2008 = _T_1962_20 & _T_671; // @[Mux.scala 27:72]
  assign _T_2029 = _T_2028 | _T_2008; // @[Mux.scala 27:72]
  assign _T_2009 = _T_1962_21 & auto_out_21_r_valid; // @[Mux.scala 27:72]
  assign _T_2030 = _T_2029 | _T_2009; // @[Mux.scala 27:72]
  assign in_0_r_valid = _T_1686 ? _T_1707 : _T_2030; // @[Xbar.scala 278:22]
  assign _T_357 = auto_in_r_ready & in_0_r_valid; // @[Decoupled.scala 40:37]
  assign _T_1721 = {_T_661,_T_659,_T_657,_T_655,_T_653}; // @[Cat.scala 29:58]
  assign _T_1711 = {_T_639,_T_637,_T_635,_T_633,_T_631}; // @[Cat.scala 29:58]
  assign _T_1717 = {_T_651,_T_649,_T_647,_T_645,_T_643,_T_641,_T_1711}; // @[Cat.scala 29:58]
  assign _T_1728 = {auto_out_21_r_valid,_T_671,_T_669,_T_667,_T_665,_T_663,_T_1721,_T_1717}; // @[Cat.scala 29:58]
  assign _T_1736 = ~_T_1735; // @[Arbiter.scala 21:30]
  assign _T_1737 = _T_1728 & _T_1736; // @[Arbiter.scala 21:28]
  assign _T_1738 = {_T_1737,auto_out_21_r_valid,_T_671,_T_669,_T_667,_T_665,_T_663,_T_1721,_T_1717}; // @[Cat.scala 29:58]
  assign _GEN_100 = {{1'd0}, _T_1738[43:1]}; // @[package.scala 208:43]
  assign _T_1740 = _T_1738 | _GEN_100; // @[package.scala 208:43]
  assign _GEN_101 = {{2'd0}, _T_1740[43:2]}; // @[package.scala 208:43]
  assign _T_1742 = _T_1740 | _GEN_101; // @[package.scala 208:43]
  assign _GEN_102 = {{4'd0}, _T_1742[43:4]}; // @[package.scala 208:43]
  assign _T_1744 = _T_1742 | _GEN_102; // @[package.scala 208:43]
  assign _GEN_103 = {{8'd0}, _T_1744[43:8]}; // @[package.scala 208:43]
  assign _T_1746 = _T_1744 | _GEN_103; // @[package.scala 208:43]
  assign _GEN_104 = {{16'd0}, _T_1746[43:16]}; // @[package.scala 208:43]
  assign _T_1748 = _T_1746 | _GEN_104; // @[package.scala 208:43]
  assign _T_1751 = {_T_1735, 22'h0}; // @[Arbiter.scala 22:66]
  assign _GEN_105 = {{1'd0}, _T_1748[43:1]}; // @[Arbiter.scala 22:58]
  assign _T_1752 = _GEN_105 | _T_1751; // @[Arbiter.scala 22:58]
  assign _T_1755 = _T_1752[43:22] & _T_1752[21:0]; // @[Arbiter.scala 23:39]
  assign _T_1756 = ~_T_1755; // @[Arbiter.scala 23:18]
  assign _T_1800 = _T_1756[0] & _T_631; // @[Xbar.scala 250:63]
  assign _T_1963_0 = _T_1686 ? _T_1800 : _T_1962_0; // @[Xbar.scala 262:23]
  assign _T_2035 = {auto_out_0_r_bits_id,auto_out_0_r_bits_data,auto_out_0_r_bits_resp,auto_out_0_r_bits_last}; // @[Mux.scala 27:72]
  assign _T_2036 = _T_1963_0 ? _T_2035 : 36'h0; // @[Mux.scala 27:72]
  assign _T_1801 = _T_1756[1] & _T_633; // @[Xbar.scala 250:63]
  assign _T_1963_1 = _T_1686 ? _T_1801 : _T_1962_1; // @[Xbar.scala 262:23]
  assign _T_2039 = {auto_out_1_r_bits_id,auto_out_1_r_bits_data,auto_out_1_r_bits_resp,auto_out_1_r_bits_last}; // @[Mux.scala 27:72]
  assign _T_2040 = _T_1963_1 ? _T_2039 : 36'h0; // @[Mux.scala 27:72]
  assign _T_2121 = _T_2036 | _T_2040; // @[Mux.scala 27:72]
  assign _T_1802 = _T_1756[2] & _T_635; // @[Xbar.scala 250:63]
  assign _T_1963_2 = _T_1686 ? _T_1802 : _T_1962_2; // @[Xbar.scala 262:23]
  assign _T_2043 = {auto_out_2_r_bits_id,auto_out_2_r_bits_data,auto_out_2_r_bits_resp,auto_out_2_r_bits_last}; // @[Mux.scala 27:72]
  assign _T_2044 = _T_1963_2 ? _T_2043 : 36'h0; // @[Mux.scala 27:72]
  assign _T_2122 = _T_2121 | _T_2044; // @[Mux.scala 27:72]
  assign _T_1803 = _T_1756[3] & _T_637; // @[Xbar.scala 250:63]
  assign _T_1963_3 = _T_1686 ? _T_1803 : _T_1962_3; // @[Xbar.scala 262:23]
  assign _T_2047 = {auto_out_3_r_bits_id,auto_out_3_r_bits_data,auto_out_3_r_bits_resp,auto_out_3_r_bits_last}; // @[Mux.scala 27:72]
  assign _T_2048 = _T_1963_3 ? _T_2047 : 36'h0; // @[Mux.scala 27:72]
  assign _T_2123 = _T_2122 | _T_2048; // @[Mux.scala 27:72]
  assign _T_1804 = _T_1756[4] & _T_639; // @[Xbar.scala 250:63]
  assign _T_1963_4 = _T_1686 ? _T_1804 : _T_1962_4; // @[Xbar.scala 262:23]
  assign _T_2051 = {auto_out_4_r_bits_id,auto_out_4_r_bits_data,auto_out_4_r_bits_resp,auto_out_4_r_bits_last}; // @[Mux.scala 27:72]
  assign _T_2052 = _T_1963_4 ? _T_2051 : 36'h0; // @[Mux.scala 27:72]
  assign _T_2124 = _T_2123 | _T_2052; // @[Mux.scala 27:72]
  assign _T_1805 = _T_1756[5] & _T_641; // @[Xbar.scala 250:63]
  assign _T_1963_5 = _T_1686 ? _T_1805 : _T_1962_5; // @[Xbar.scala 262:23]
  assign _T_2055 = {auto_out_5_r_bits_id,auto_out_5_r_bits_data,auto_out_5_r_bits_resp,auto_out_5_r_bits_last}; // @[Mux.scala 27:72]
  assign _T_2056 = _T_1963_5 ? _T_2055 : 36'h0; // @[Mux.scala 27:72]
  assign _T_2125 = _T_2124 | _T_2056; // @[Mux.scala 27:72]
  assign _T_1806 = _T_1756[6] & _T_643; // @[Xbar.scala 250:63]
  assign _T_1963_6 = _T_1686 ? _T_1806 : _T_1962_6; // @[Xbar.scala 262:23]
  assign _T_2059 = {auto_out_6_r_bits_id,auto_out_6_r_bits_data,auto_out_6_r_bits_resp,auto_out_6_r_bits_last}; // @[Mux.scala 27:72]
  assign _T_2060 = _T_1963_6 ? _T_2059 : 36'h0; // @[Mux.scala 27:72]
  assign _T_2126 = _T_2125 | _T_2060; // @[Mux.scala 27:72]
  assign _T_1807 = _T_1756[7] & _T_645; // @[Xbar.scala 250:63]
  assign _T_1963_7 = _T_1686 ? _T_1807 : _T_1962_7; // @[Xbar.scala 262:23]
  assign _T_2063 = {auto_out_7_r_bits_id,auto_out_7_r_bits_data,auto_out_7_r_bits_resp,auto_out_7_r_bits_last}; // @[Mux.scala 27:72]
  assign _T_2064 = _T_1963_7 ? _T_2063 : 36'h0; // @[Mux.scala 27:72]
  assign _T_2127 = _T_2126 | _T_2064; // @[Mux.scala 27:72]
  assign _T_1808 = _T_1756[8] & _T_647; // @[Xbar.scala 250:63]
  assign _T_1963_8 = _T_1686 ? _T_1808 : _T_1962_8; // @[Xbar.scala 262:23]
  assign _T_2067 = {auto_out_8_r_bits_id,auto_out_8_r_bits_data,auto_out_8_r_bits_resp,auto_out_8_r_bits_last}; // @[Mux.scala 27:72]
  assign _T_2068 = _T_1963_8 ? _T_2067 : 36'h0; // @[Mux.scala 27:72]
  assign _T_2128 = _T_2127 | _T_2068; // @[Mux.scala 27:72]
  assign _T_1809 = _T_1756[9] & _T_649; // @[Xbar.scala 250:63]
  assign _T_1963_9 = _T_1686 ? _T_1809 : _T_1962_9; // @[Xbar.scala 262:23]
  assign _T_2071 = {auto_out_9_r_bits_id,auto_out_9_r_bits_data,auto_out_9_r_bits_resp,auto_out_9_r_bits_last}; // @[Mux.scala 27:72]
  assign _T_2072 = _T_1963_9 ? _T_2071 : 36'h0; // @[Mux.scala 27:72]
  assign _T_2129 = _T_2128 | _T_2072; // @[Mux.scala 27:72]
  assign _T_1810 = _T_1756[10] & _T_651; // @[Xbar.scala 250:63]
  assign _T_1963_10 = _T_1686 ? _T_1810 : _T_1962_10; // @[Xbar.scala 262:23]
  assign _T_2075 = {auto_out_10_r_bits_id,auto_out_10_r_bits_data,auto_out_10_r_bits_resp,auto_out_10_r_bits_last}; // @[Mux.scala 27:72]
  assign _T_2076 = _T_1963_10 ? _T_2075 : 36'h0; // @[Mux.scala 27:72]
  assign _T_2130 = _T_2129 | _T_2076; // @[Mux.scala 27:72]
  assign _T_1811 = _T_1756[11] & _T_653; // @[Xbar.scala 250:63]
  assign _T_1963_11 = _T_1686 ? _T_1811 : _T_1962_11; // @[Xbar.scala 262:23]
  assign _T_2079 = {auto_out_11_r_bits_id,auto_out_11_r_bits_data,auto_out_11_r_bits_resp,auto_out_11_r_bits_last}; // @[Mux.scala 27:72]
  assign _T_2080 = _T_1963_11 ? _T_2079 : 36'h0; // @[Mux.scala 27:72]
  assign _T_2131 = _T_2130 | _T_2080; // @[Mux.scala 27:72]
  assign _T_1812 = _T_1756[12] & _T_655; // @[Xbar.scala 250:63]
  assign _T_1963_12 = _T_1686 ? _T_1812 : _T_1962_12; // @[Xbar.scala 262:23]
  assign _T_2083 = {auto_out_12_r_bits_id,auto_out_12_r_bits_data,auto_out_12_r_bits_resp,auto_out_12_r_bits_last}; // @[Mux.scala 27:72]
  assign _T_2084 = _T_1963_12 ? _T_2083 : 36'h0; // @[Mux.scala 27:72]
  assign _T_2132 = _T_2131 | _T_2084; // @[Mux.scala 27:72]
  assign _T_1813 = _T_1756[13] & _T_657; // @[Xbar.scala 250:63]
  assign _T_1963_13 = _T_1686 ? _T_1813 : _T_1962_13; // @[Xbar.scala 262:23]
  assign _T_2087 = {auto_out_13_r_bits_id,auto_out_13_r_bits_data,auto_out_13_r_bits_resp,auto_out_13_r_bits_last}; // @[Mux.scala 27:72]
  assign _T_2088 = _T_1963_13 ? _T_2087 : 36'h0; // @[Mux.scala 27:72]
  assign _T_2133 = _T_2132 | _T_2088; // @[Mux.scala 27:72]
  assign _T_1814 = _T_1756[14] & _T_659; // @[Xbar.scala 250:63]
  assign _T_1963_14 = _T_1686 ? _T_1814 : _T_1962_14; // @[Xbar.scala 262:23]
  assign _T_2091 = {auto_out_14_r_bits_id,auto_out_14_r_bits_data,auto_out_14_r_bits_resp,auto_out_14_r_bits_last}; // @[Mux.scala 27:72]
  assign _T_2092 = _T_1963_14 ? _T_2091 : 36'h0; // @[Mux.scala 27:72]
  assign _T_2134 = _T_2133 | _T_2092; // @[Mux.scala 27:72]
  assign _T_1815 = _T_1756[15] & _T_661; // @[Xbar.scala 250:63]
  assign _T_1963_15 = _T_1686 ? _T_1815 : _T_1962_15; // @[Xbar.scala 262:23]
  assign _T_2095 = {auto_out_15_r_bits_id,auto_out_15_r_bits_data,auto_out_15_r_bits_resp,auto_out_15_r_bits_last}; // @[Mux.scala 27:72]
  assign _T_2096 = _T_1963_15 ? _T_2095 : 36'h0; // @[Mux.scala 27:72]
  assign _T_2135 = _T_2134 | _T_2096; // @[Mux.scala 27:72]
  assign _T_1816 = _T_1756[16] & _T_663; // @[Xbar.scala 250:63]
  assign _T_1963_16 = _T_1686 ? _T_1816 : _T_1962_16; // @[Xbar.scala 262:23]
  assign _T_2099 = {auto_out_16_r_bits_id,auto_out_16_r_bits_data,auto_out_16_r_bits_resp,auto_out_16_r_bits_last}; // @[Mux.scala 27:72]
  assign _T_2100 = _T_1963_16 ? _T_2099 : 36'h0; // @[Mux.scala 27:72]
  assign _T_2136 = _T_2135 | _T_2100; // @[Mux.scala 27:72]
  assign _T_1817 = _T_1756[17] & _T_665; // @[Xbar.scala 250:63]
  assign _T_1963_17 = _T_1686 ? _T_1817 : _T_1962_17; // @[Xbar.scala 262:23]
  assign _T_2103 = {auto_out_17_r_bits_id,auto_out_17_r_bits_data,auto_out_17_r_bits_resp,auto_out_17_r_bits_last}; // @[Mux.scala 27:72]
  assign _T_2104 = _T_1963_17 ? _T_2103 : 36'h0; // @[Mux.scala 27:72]
  assign _T_2137 = _T_2136 | _T_2104; // @[Mux.scala 27:72]
  assign _T_1818 = _T_1756[18] & _T_667; // @[Xbar.scala 250:63]
  assign _T_1963_18 = _T_1686 ? _T_1818 : _T_1962_18; // @[Xbar.scala 262:23]
  assign _T_2107 = {auto_out_18_r_bits_id,auto_out_18_r_bits_data,auto_out_18_r_bits_resp,auto_out_18_r_bits_last}; // @[Mux.scala 27:72]
  assign _T_2108 = _T_1963_18 ? _T_2107 : 36'h0; // @[Mux.scala 27:72]
  assign _T_2138 = _T_2137 | _T_2108; // @[Mux.scala 27:72]
  assign _T_1819 = _T_1756[19] & _T_669; // @[Xbar.scala 250:63]
  assign _T_1963_19 = _T_1686 ? _T_1819 : _T_1962_19; // @[Xbar.scala 262:23]
  assign _T_2111 = {auto_out_19_r_bits_id,auto_out_19_r_bits_data,auto_out_19_r_bits_resp,auto_out_19_r_bits_last}; // @[Mux.scala 27:72]
  assign _T_2112 = _T_1963_19 ? _T_2111 : 36'h0; // @[Mux.scala 27:72]
  assign _T_2139 = _T_2138 | _T_2112; // @[Mux.scala 27:72]
  assign _T_1820 = _T_1756[20] & _T_671; // @[Xbar.scala 250:63]
  assign _T_1963_20 = _T_1686 ? _T_1820 : _T_1962_20; // @[Xbar.scala 262:23]
  assign _T_2115 = {auto_out_20_r_bits_id,auto_out_20_r_bits_data,auto_out_20_r_bits_resp,auto_out_20_r_bits_last}; // @[Mux.scala 27:72]
  assign _T_2116 = _T_1963_20 ? _T_2115 : 36'h0; // @[Mux.scala 27:72]
  assign _T_2140 = _T_2139 | _T_2116; // @[Mux.scala 27:72]
  assign _T_1821 = _T_1756[21] & auto_out_21_r_valid; // @[Xbar.scala 250:63]
  assign _T_1963_21 = _T_1686 ? _T_1821 : _T_1962_21; // @[Xbar.scala 262:23]
  assign _T_2119 = {1'h0,auto_out_21_r_bits_data,auto_out_21_r_bits_resp,auto_out_21_r_bits_last}; // @[Mux.scala 27:72]
  assign _T_2120 = _T_1963_21 ? _T_2119 : 36'h0; // @[Mux.scala 27:72]
  assign _T_2141 = _T_2140 | _T_2120; // @[Mux.scala 27:72]
  assign in_0_r_bits_last = _T_2141[0]; // @[Mux.scala 27:72]
  assign _T_359 = _T_357 & in_0_r_bits_last; // @[Xbar.scala 120:45]
  assign _GEN_106 = {{2'd0}, _T_355}; // @[Xbar.scala 106:30]
  assign _T_363 = _T_360 + _GEN_106; // @[Xbar.scala 106:30]
  assign _GEN_107 = {{2'd0}, _T_359}; // @[Xbar.scala 106:48]
  assign _T_365 = _T_363 - _GEN_107; // @[Xbar.scala 106:48]
  assign _T_366 = ~_T_359; // @[Xbar.scala 107:23]
  assign _T_367 = _T_360 != 3'h0; // @[Xbar.scala 107:43]
  assign _T_368 = _T_366 | _T_367; // @[Xbar.scala 107:34]
  assign _T_370 = _T_368 | reset; // @[Xbar.scala 107:22]
  assign _T_371 = ~_T_370; // @[Xbar.scala 107:22]
  assign _T_372 = ~_T_355; // @[Xbar.scala 108:23]
  assign _T_374 = _T_372 | _T_381; // @[Xbar.scala 108:34]
  assign _T_376 = _T_374 | reset; // @[Xbar.scala 108:22]
  assign _T_377 = ~_T_376; // @[Xbar.scala 108:22]
  assign _T_519 = requestAWIO_0_0 & auto_out_0_aw_ready; // @[Mux.scala 27:72]
  assign _T_520 = requestAWIO_0_1 & auto_out_1_aw_ready; // @[Mux.scala 27:72]
  assign _T_541 = _T_519 | _T_520; // @[Mux.scala 27:72]
  assign _T_521 = requestAWIO_0_2 & auto_out_2_aw_ready; // @[Mux.scala 27:72]
  assign _T_542 = _T_541 | _T_521; // @[Mux.scala 27:72]
  assign _T_522 = requestAWIO_0_3 & auto_out_3_aw_ready; // @[Mux.scala 27:72]
  assign _T_543 = _T_542 | _T_522; // @[Mux.scala 27:72]
  assign _T_523 = requestAWIO_0_4 & auto_out_4_aw_ready; // @[Mux.scala 27:72]
  assign _T_544 = _T_543 | _T_523; // @[Mux.scala 27:72]
  assign _T_524 = requestAWIO_0_5 & auto_out_5_aw_ready; // @[Mux.scala 27:72]
  assign _T_545 = _T_544 | _T_524; // @[Mux.scala 27:72]
  assign _T_525 = requestAWIO_0_6 & auto_out_6_aw_ready; // @[Mux.scala 27:72]
  assign _T_546 = _T_545 | _T_525; // @[Mux.scala 27:72]
  assign _T_526 = requestAWIO_0_7 & auto_out_7_aw_ready; // @[Mux.scala 27:72]
  assign _T_547 = _T_546 | _T_526; // @[Mux.scala 27:72]
  assign _T_527 = requestAWIO_0_8 & auto_out_8_aw_ready; // @[Mux.scala 27:72]
  assign _T_548 = _T_547 | _T_527; // @[Mux.scala 27:72]
  assign _T_528 = requestAWIO_0_9 & auto_out_9_aw_ready; // @[Mux.scala 27:72]
  assign _T_549 = _T_548 | _T_528; // @[Mux.scala 27:72]
  assign _T_529 = requestAWIO_0_10 & auto_out_10_aw_ready; // @[Mux.scala 27:72]
  assign _T_550 = _T_549 | _T_529; // @[Mux.scala 27:72]
  assign _T_530 = requestAWIO_0_11 & auto_out_11_aw_ready; // @[Mux.scala 27:72]
  assign _T_551 = _T_550 | _T_530; // @[Mux.scala 27:72]
  assign _T_531 = requestAWIO_0_12 & auto_out_12_aw_ready; // @[Mux.scala 27:72]
  assign _T_552 = _T_551 | _T_531; // @[Mux.scala 27:72]
  assign _T_532 = requestAWIO_0_13 & auto_out_13_aw_ready; // @[Mux.scala 27:72]
  assign _T_553 = _T_552 | _T_532; // @[Mux.scala 27:72]
  assign _T_533 = requestAWIO_0_14 & auto_out_14_aw_ready; // @[Mux.scala 27:72]
  assign _T_554 = _T_553 | _T_533; // @[Mux.scala 27:72]
  assign _T_534 = requestAWIO_0_15 & auto_out_15_aw_ready; // @[Mux.scala 27:72]
  assign _T_555 = _T_554 | _T_534; // @[Mux.scala 27:72]
  assign _T_535 = requestAWIO_0_16 & auto_out_16_aw_ready; // @[Mux.scala 27:72]
  assign _T_556 = _T_555 | _T_535; // @[Mux.scala 27:72]
  assign _T_536 = requestAWIO_0_17 & auto_out_17_aw_ready; // @[Mux.scala 27:72]
  assign _T_557 = _T_556 | _T_536; // @[Mux.scala 27:72]
  assign _T_537 = requestAWIO_0_18 & auto_out_18_aw_ready; // @[Mux.scala 27:72]
  assign _T_558 = _T_557 | _T_537; // @[Mux.scala 27:72]
  assign _T_538 = requestAWIO_0_19 & auto_out_19_aw_ready; // @[Mux.scala 27:72]
  assign _T_559 = _T_558 | _T_538; // @[Mux.scala 27:72]
  assign _T_539 = requestAWIO_0_20 & auto_out_20_aw_ready; // @[Mux.scala 27:72]
  assign _T_560 = _T_559 | _T_539; // @[Mux.scala 27:72]
  assign _T_540 = requestAWIO_0_21 & auto_out_21_aw_ready; // @[Mux.scala 27:72]
  assign in_0_aw_ready = _T_560 | _T_540; // @[Mux.scala 27:72]
  assign _T_418 = _T_414 | awIn_0_io_enq_ready; // @[Xbar.scala 139:57]
  assign _T_419 = in_0_aw_ready & _T_418; // @[Xbar.scala 139:45]
  assign _T_407 = _T_388 == 3'h0; // @[Xbar.scala 112:22]
  assign _T_406 = _T_389 == _T_354; // @[Xbar.scala 111:75]
  assign _T_408 = _T_407 | _T_406; // @[Xbar.scala 112:34]
  assign _T_409 = _T_388 != 3'h7; // @[Xbar.scala 112:80]
  assign _T_411 = _T_408 & _T_409; // @[Xbar.scala 112:48]
  assign io_in_0_aw_ready = _T_419 & _T_411; // @[Xbar.scala 139:82]
  assign _T_384 = io_in_0_aw_ready & auto_in_aw_valid; // @[Decoupled.scala 40:37]
  assign _T_675 = auto_out_0_b_valid & requestBOI_0_0; // @[Xbar.scala 222:40]
  assign _T_677 = auto_out_1_b_valid & requestBOI_1_0; // @[Xbar.scala 222:40]
  assign _T_2149 = _T_675 | _T_677; // @[Xbar.scala 246:36]
  assign _T_679 = auto_out_2_b_valid & requestBOI_2_0; // @[Xbar.scala 222:40]
  assign _T_2150 = _T_2149 | _T_679; // @[Xbar.scala 246:36]
  assign _T_681 = auto_out_3_b_valid & requestBOI_3_0; // @[Xbar.scala 222:40]
  assign _T_2151 = _T_2150 | _T_681; // @[Xbar.scala 246:36]
  assign _T_683 = auto_out_4_b_valid & requestBOI_4_0; // @[Xbar.scala 222:40]
  assign _T_2152 = _T_2151 | _T_683; // @[Xbar.scala 246:36]
  assign _T_685 = auto_out_5_b_valid & requestBOI_5_0; // @[Xbar.scala 222:40]
  assign _T_2153 = _T_2152 | _T_685; // @[Xbar.scala 246:36]
  assign _T_687 = auto_out_6_b_valid & requestBOI_6_0; // @[Xbar.scala 222:40]
  assign _T_2154 = _T_2153 | _T_687; // @[Xbar.scala 246:36]
  assign _T_689 = auto_out_7_b_valid & requestBOI_7_0; // @[Xbar.scala 222:40]
  assign _T_2155 = _T_2154 | _T_689; // @[Xbar.scala 246:36]
  assign _T_691 = auto_out_8_b_valid & requestBOI_8_0; // @[Xbar.scala 222:40]
  assign _T_2156 = _T_2155 | _T_691; // @[Xbar.scala 246:36]
  assign _T_693 = auto_out_9_b_valid & requestBOI_9_0; // @[Xbar.scala 222:40]
  assign _T_2157 = _T_2156 | _T_693; // @[Xbar.scala 246:36]
  assign _T_695 = auto_out_10_b_valid & requestBOI_10_0; // @[Xbar.scala 222:40]
  assign _T_2158 = _T_2157 | _T_695; // @[Xbar.scala 246:36]
  assign _T_697 = auto_out_11_b_valid & requestBOI_11_0; // @[Xbar.scala 222:40]
  assign _T_2159 = _T_2158 | _T_697; // @[Xbar.scala 246:36]
  assign _T_699 = auto_out_12_b_valid & requestBOI_12_0; // @[Xbar.scala 222:40]
  assign _T_2160 = _T_2159 | _T_699; // @[Xbar.scala 246:36]
  assign _T_701 = auto_out_13_b_valid & requestBOI_13_0; // @[Xbar.scala 222:40]
  assign _T_2161 = _T_2160 | _T_701; // @[Xbar.scala 246:36]
  assign _T_703 = auto_out_14_b_valid & requestBOI_14_0; // @[Xbar.scala 222:40]
  assign _T_2162 = _T_2161 | _T_703; // @[Xbar.scala 246:36]
  assign _T_705 = auto_out_15_b_valid & requestBOI_15_0; // @[Xbar.scala 222:40]
  assign _T_2163 = _T_2162 | _T_705; // @[Xbar.scala 246:36]
  assign _T_707 = auto_out_16_b_valid & requestBOI_16_0; // @[Xbar.scala 222:40]
  assign _T_2164 = _T_2163 | _T_707; // @[Xbar.scala 246:36]
  assign _T_709 = auto_out_17_b_valid & requestBOI_17_0; // @[Xbar.scala 222:40]
  assign _T_2165 = _T_2164 | _T_709; // @[Xbar.scala 246:36]
  assign _T_711 = auto_out_18_b_valid & requestBOI_18_0; // @[Xbar.scala 222:40]
  assign _T_2166 = _T_2165 | _T_711; // @[Xbar.scala 246:36]
  assign _T_713 = auto_out_19_b_valid & requestBOI_19_0; // @[Xbar.scala 222:40]
  assign _T_2167 = _T_2166 | _T_713; // @[Xbar.scala 246:36]
  assign _T_715 = auto_out_20_b_valid & requestBOI_20_0; // @[Xbar.scala 222:40]
  assign _T_2168 = _T_2167 | _T_715; // @[Xbar.scala 246:36]
  assign _T_2169 = _T_2168 | auto_out_21_b_valid; // @[Xbar.scala 246:36]
  assign _T_2450 = _T_2424_0 & _T_675; // @[Mux.scala 27:72]
  assign _T_2451 = _T_2424_1 & _T_677; // @[Mux.scala 27:72]
  assign _T_2472 = _T_2450 | _T_2451; // @[Mux.scala 27:72]
  assign _T_2452 = _T_2424_2 & _T_679; // @[Mux.scala 27:72]
  assign _T_2473 = _T_2472 | _T_2452; // @[Mux.scala 27:72]
  assign _T_2453 = _T_2424_3 & _T_681; // @[Mux.scala 27:72]
  assign _T_2474 = _T_2473 | _T_2453; // @[Mux.scala 27:72]
  assign _T_2454 = _T_2424_4 & _T_683; // @[Mux.scala 27:72]
  assign _T_2475 = _T_2474 | _T_2454; // @[Mux.scala 27:72]
  assign _T_2455 = _T_2424_5 & _T_685; // @[Mux.scala 27:72]
  assign _T_2476 = _T_2475 | _T_2455; // @[Mux.scala 27:72]
  assign _T_2456 = _T_2424_6 & _T_687; // @[Mux.scala 27:72]
  assign _T_2477 = _T_2476 | _T_2456; // @[Mux.scala 27:72]
  assign _T_2457 = _T_2424_7 & _T_689; // @[Mux.scala 27:72]
  assign _T_2478 = _T_2477 | _T_2457; // @[Mux.scala 27:72]
  assign _T_2458 = _T_2424_8 & _T_691; // @[Mux.scala 27:72]
  assign _T_2479 = _T_2478 | _T_2458; // @[Mux.scala 27:72]
  assign _T_2459 = _T_2424_9 & _T_693; // @[Mux.scala 27:72]
  assign _T_2480 = _T_2479 | _T_2459; // @[Mux.scala 27:72]
  assign _T_2460 = _T_2424_10 & _T_695; // @[Mux.scala 27:72]
  assign _T_2481 = _T_2480 | _T_2460; // @[Mux.scala 27:72]
  assign _T_2461 = _T_2424_11 & _T_697; // @[Mux.scala 27:72]
  assign _T_2482 = _T_2481 | _T_2461; // @[Mux.scala 27:72]
  assign _T_2462 = _T_2424_12 & _T_699; // @[Mux.scala 27:72]
  assign _T_2483 = _T_2482 | _T_2462; // @[Mux.scala 27:72]
  assign _T_2463 = _T_2424_13 & _T_701; // @[Mux.scala 27:72]
  assign _T_2484 = _T_2483 | _T_2463; // @[Mux.scala 27:72]
  assign _T_2464 = _T_2424_14 & _T_703; // @[Mux.scala 27:72]
  assign _T_2485 = _T_2484 | _T_2464; // @[Mux.scala 27:72]
  assign _T_2465 = _T_2424_15 & _T_705; // @[Mux.scala 27:72]
  assign _T_2486 = _T_2485 | _T_2465; // @[Mux.scala 27:72]
  assign _T_2466 = _T_2424_16 & _T_707; // @[Mux.scala 27:72]
  assign _T_2487 = _T_2486 | _T_2466; // @[Mux.scala 27:72]
  assign _T_2467 = _T_2424_17 & _T_709; // @[Mux.scala 27:72]
  assign _T_2488 = _T_2487 | _T_2467; // @[Mux.scala 27:72]
  assign _T_2468 = _T_2424_18 & _T_711; // @[Mux.scala 27:72]
  assign _T_2489 = _T_2488 | _T_2468; // @[Mux.scala 27:72]
  assign _T_2469 = _T_2424_19 & _T_713; // @[Mux.scala 27:72]
  assign _T_2490 = _T_2489 | _T_2469; // @[Mux.scala 27:72]
  assign _T_2470 = _T_2424_20 & _T_715; // @[Mux.scala 27:72]
  assign _T_2491 = _T_2490 | _T_2470; // @[Mux.scala 27:72]
  assign _T_2471 = _T_2424_21 & auto_out_21_b_valid; // @[Mux.scala 27:72]
  assign _T_2492 = _T_2491 | _T_2471; // @[Mux.scala 27:72]
  assign in_0_b_valid = _T_2148 ? _T_2169 : _T_2492; // @[Xbar.scala 278:22]
  assign _T_386 = auto_in_b_ready & in_0_b_valid; // @[Decoupled.scala 40:37]
  assign _GEN_108 = {{2'd0}, _T_384}; // @[Xbar.scala 106:30]
  assign _T_391 = _T_388 + _GEN_108; // @[Xbar.scala 106:30]
  assign _GEN_109 = {{2'd0}, _T_386}; // @[Xbar.scala 106:48]
  assign _T_393 = _T_391 - _GEN_109; // @[Xbar.scala 106:48]
  assign _T_394 = ~_T_386; // @[Xbar.scala 107:23]
  assign _T_395 = _T_388 != 3'h0; // @[Xbar.scala 107:43]
  assign _T_396 = _T_394 | _T_395; // @[Xbar.scala 107:34]
  assign _T_398 = _T_396 | reset; // @[Xbar.scala 107:22]
  assign _T_399 = ~_T_398; // @[Xbar.scala 107:22]
  assign _T_400 = ~_T_384; // @[Xbar.scala 108:23]
  assign _T_402 = _T_400 | _T_409; // @[Xbar.scala 108:34]
  assign _T_404 = _T_402 | reset; // @[Xbar.scala 108:22]
  assign _T_405 = ~_T_404; // @[Xbar.scala 108:22]
  assign in_0_ar_valid = auto_in_ar_valid & _T_383; // @[Xbar.scala 129:45]
  assign _T_416 = auto_in_aw_valid & _T_418; // @[Xbar.scala 138:45]
  assign in_0_aw_valid = _T_416 & _T_411; // @[Xbar.scala 138:82]
  assign _T_421 = ~_T_414; // @[Xbar.scala 140:54]
  assign _T_423 = awIn_0_io_enq_ready & awIn_0_io_enq_valid; // @[Decoupled.scala 40:37]
  assign _GEN_2 = _T_423 | _T_414; // @[Xbar.scala 141:38]
  assign _T_424 = in_0_aw_ready & in_0_aw_valid; // @[Decoupled.scala 40:37]
  assign in_0_w_valid = auto_in_w_valid & awIn_0_io_deq_valid; // @[Xbar.scala 145:43]
  assign _T_586 = requestWIO_0_0 & auto_out_0_w_ready; // @[Mux.scala 27:72]
  assign _T_587 = requestWIO_0_1 & auto_out_1_w_ready; // @[Mux.scala 27:72]
  assign _T_608 = _T_586 | _T_587; // @[Mux.scala 27:72]
  assign _T_588 = requestWIO_0_2 & auto_out_2_w_ready; // @[Mux.scala 27:72]
  assign _T_609 = _T_608 | _T_588; // @[Mux.scala 27:72]
  assign _T_589 = requestWIO_0_3 & auto_out_3_w_ready; // @[Mux.scala 27:72]
  assign _T_610 = _T_609 | _T_589; // @[Mux.scala 27:72]
  assign _T_590 = requestWIO_0_4 & auto_out_4_w_ready; // @[Mux.scala 27:72]
  assign _T_611 = _T_610 | _T_590; // @[Mux.scala 27:72]
  assign _T_591 = requestWIO_0_5 & auto_out_5_w_ready; // @[Mux.scala 27:72]
  assign _T_612 = _T_611 | _T_591; // @[Mux.scala 27:72]
  assign _T_592 = requestWIO_0_6 & auto_out_6_w_ready; // @[Mux.scala 27:72]
  assign _T_613 = _T_612 | _T_592; // @[Mux.scala 27:72]
  assign _T_593 = requestWIO_0_7 & auto_out_7_w_ready; // @[Mux.scala 27:72]
  assign _T_614 = _T_613 | _T_593; // @[Mux.scala 27:72]
  assign _T_594 = requestWIO_0_8 & auto_out_8_w_ready; // @[Mux.scala 27:72]
  assign _T_615 = _T_614 | _T_594; // @[Mux.scala 27:72]
  assign _T_595 = requestWIO_0_9 & auto_out_9_w_ready; // @[Mux.scala 27:72]
  assign _T_616 = _T_615 | _T_595; // @[Mux.scala 27:72]
  assign _T_596 = requestWIO_0_10 & auto_out_10_w_ready; // @[Mux.scala 27:72]
  assign _T_617 = _T_616 | _T_596; // @[Mux.scala 27:72]
  assign _T_597 = requestWIO_0_11 & auto_out_11_w_ready; // @[Mux.scala 27:72]
  assign _T_618 = _T_617 | _T_597; // @[Mux.scala 27:72]
  assign _T_598 = requestWIO_0_12 & auto_out_12_w_ready; // @[Mux.scala 27:72]
  assign _T_619 = _T_618 | _T_598; // @[Mux.scala 27:72]
  assign _T_599 = requestWIO_0_13 & auto_out_13_w_ready; // @[Mux.scala 27:72]
  assign _T_620 = _T_619 | _T_599; // @[Mux.scala 27:72]
  assign _T_600 = requestWIO_0_14 & auto_out_14_w_ready; // @[Mux.scala 27:72]
  assign _T_621 = _T_620 | _T_600; // @[Mux.scala 27:72]
  assign _T_601 = requestWIO_0_15 & auto_out_15_w_ready; // @[Mux.scala 27:72]
  assign _T_622 = _T_621 | _T_601; // @[Mux.scala 27:72]
  assign _T_602 = requestWIO_0_16 & auto_out_16_w_ready; // @[Mux.scala 27:72]
  assign _T_623 = _T_622 | _T_602; // @[Mux.scala 27:72]
  assign _T_603 = requestWIO_0_17 & auto_out_17_w_ready; // @[Mux.scala 27:72]
  assign _T_624 = _T_623 | _T_603; // @[Mux.scala 27:72]
  assign _T_604 = requestWIO_0_18 & auto_out_18_w_ready; // @[Mux.scala 27:72]
  assign _T_625 = _T_624 | _T_604; // @[Mux.scala 27:72]
  assign _T_605 = requestWIO_0_19 & auto_out_19_w_ready; // @[Mux.scala 27:72]
  assign _T_626 = _T_625 | _T_605; // @[Mux.scala 27:72]
  assign _T_606 = requestWIO_0_20 & auto_out_20_w_ready; // @[Mux.scala 27:72]
  assign _T_627 = _T_626 | _T_606; // @[Mux.scala 27:72]
  assign _T_607 = requestWIO_0_21 & auto_out_21_w_ready; // @[Mux.scala 27:72]
  assign in_0_w_ready = _T_627 | _T_607; // @[Mux.scala 27:72]
  assign _T_427 = auto_in_w_valid & auto_in_w_bits_last; // @[Xbar.scala 147:50]
  assign out_0_ar_valid = in_0_ar_valid & requestARIO_0_0; // @[Xbar.scala 222:40]
  assign out_1_ar_valid = in_0_ar_valid & requestARIO_0_1; // @[Xbar.scala 222:40]
  assign out_2_ar_valid = in_0_ar_valid & requestARIO_0_2; // @[Xbar.scala 222:40]
  assign out_3_ar_valid = in_0_ar_valid & requestARIO_0_3; // @[Xbar.scala 222:40]
  assign out_4_ar_valid = in_0_ar_valid & requestARIO_0_4; // @[Xbar.scala 222:40]
  assign out_5_ar_valid = in_0_ar_valid & requestARIO_0_5; // @[Xbar.scala 222:40]
  assign out_6_ar_valid = in_0_ar_valid & requestARIO_0_6; // @[Xbar.scala 222:40]
  assign out_7_ar_valid = in_0_ar_valid & requestARIO_0_7; // @[Xbar.scala 222:40]
  assign out_8_ar_valid = in_0_ar_valid & requestARIO_0_8; // @[Xbar.scala 222:40]
  assign out_9_ar_valid = in_0_ar_valid & requestARIO_0_9; // @[Xbar.scala 222:40]
  assign out_10_ar_valid = in_0_ar_valid & requestARIO_0_10; // @[Xbar.scala 222:40]
  assign out_11_ar_valid = in_0_ar_valid & requestARIO_0_11; // @[Xbar.scala 222:40]
  assign out_12_ar_valid = in_0_ar_valid & requestARIO_0_12; // @[Xbar.scala 222:40]
  assign out_13_ar_valid = in_0_ar_valid & requestARIO_0_13; // @[Xbar.scala 222:40]
  assign out_14_ar_valid = in_0_ar_valid & requestARIO_0_14; // @[Xbar.scala 222:40]
  assign out_15_ar_valid = in_0_ar_valid & requestARIO_0_15; // @[Xbar.scala 222:40]
  assign out_16_ar_valid = in_0_ar_valid & requestARIO_0_16; // @[Xbar.scala 222:40]
  assign out_17_ar_valid = in_0_ar_valid & requestARIO_0_17; // @[Xbar.scala 222:40]
  assign out_18_ar_valid = in_0_ar_valid & requestARIO_0_18; // @[Xbar.scala 222:40]
  assign out_19_ar_valid = in_0_ar_valid & requestARIO_0_19; // @[Xbar.scala 222:40]
  assign out_20_ar_valid = in_0_ar_valid & requestARIO_0_20; // @[Xbar.scala 222:40]
  assign out_21_ar_valid = in_0_ar_valid & requestARIO_0_21; // @[Xbar.scala 222:40]
  assign out_0_aw_valid = in_0_aw_valid & requestAWIO_0_0; // @[Xbar.scala 222:40]
  assign out_1_aw_valid = in_0_aw_valid & requestAWIO_0_1; // @[Xbar.scala 222:40]
  assign out_2_aw_valid = in_0_aw_valid & requestAWIO_0_2; // @[Xbar.scala 222:40]
  assign out_3_aw_valid = in_0_aw_valid & requestAWIO_0_3; // @[Xbar.scala 222:40]
  assign out_4_aw_valid = in_0_aw_valid & requestAWIO_0_4; // @[Xbar.scala 222:40]
  assign out_5_aw_valid = in_0_aw_valid & requestAWIO_0_5; // @[Xbar.scala 222:40]
  assign out_6_aw_valid = in_0_aw_valid & requestAWIO_0_6; // @[Xbar.scala 222:40]
  assign out_7_aw_valid = in_0_aw_valid & requestAWIO_0_7; // @[Xbar.scala 222:40]
  assign out_8_aw_valid = in_0_aw_valid & requestAWIO_0_8; // @[Xbar.scala 222:40]
  assign out_9_aw_valid = in_0_aw_valid & requestAWIO_0_9; // @[Xbar.scala 222:40]
  assign out_10_aw_valid = in_0_aw_valid & requestAWIO_0_10; // @[Xbar.scala 222:40]
  assign out_11_aw_valid = in_0_aw_valid & requestAWIO_0_11; // @[Xbar.scala 222:40]
  assign out_12_aw_valid = in_0_aw_valid & requestAWIO_0_12; // @[Xbar.scala 222:40]
  assign out_13_aw_valid = in_0_aw_valid & requestAWIO_0_13; // @[Xbar.scala 222:40]
  assign out_14_aw_valid = in_0_aw_valid & requestAWIO_0_14; // @[Xbar.scala 222:40]
  assign out_15_aw_valid = in_0_aw_valid & requestAWIO_0_15; // @[Xbar.scala 222:40]
  assign out_16_aw_valid = in_0_aw_valid & requestAWIO_0_16; // @[Xbar.scala 222:40]
  assign out_17_aw_valid = in_0_aw_valid & requestAWIO_0_17; // @[Xbar.scala 222:40]
  assign out_18_aw_valid = in_0_aw_valid & requestAWIO_0_18; // @[Xbar.scala 222:40]
  assign out_19_aw_valid = in_0_aw_valid & requestAWIO_0_19; // @[Xbar.scala 222:40]
  assign out_20_aw_valid = in_0_aw_valid & requestAWIO_0_20; // @[Xbar.scala 222:40]
  assign out_21_aw_valid = in_0_aw_valid & requestAWIO_0_21; // @[Xbar.scala 222:40]
  assign _T_724 = ~out_0_aw_valid; // @[Xbar.scala 256:60]
  assign _T_730 = _T_724 | out_0_aw_valid; // @[Xbar.scala 258:23]
  assign _T_732 = _T_730 | reset; // @[Xbar.scala 258:12]
  assign _T_733 = ~_T_732; // @[Xbar.scala 258:12]
  assign _T_745 = ~out_0_ar_valid; // @[Xbar.scala 256:60]
  assign _T_751 = _T_745 | out_0_ar_valid; // @[Xbar.scala 258:23]
  assign _T_753 = _T_751 | reset; // @[Xbar.scala 258:12]
  assign _T_754 = ~_T_753; // @[Xbar.scala 258:12]
  assign _T_768 = ~out_1_aw_valid; // @[Xbar.scala 256:60]
  assign _T_774 = _T_768 | out_1_aw_valid; // @[Xbar.scala 258:23]
  assign _T_776 = _T_774 | reset; // @[Xbar.scala 258:12]
  assign _T_777 = ~_T_776; // @[Xbar.scala 258:12]
  assign _T_789 = ~out_1_ar_valid; // @[Xbar.scala 256:60]
  assign _T_795 = _T_789 | out_1_ar_valid; // @[Xbar.scala 258:23]
  assign _T_797 = _T_795 | reset; // @[Xbar.scala 258:12]
  assign _T_798 = ~_T_797; // @[Xbar.scala 258:12]
  assign _T_812 = ~out_2_aw_valid; // @[Xbar.scala 256:60]
  assign _T_818 = _T_812 | out_2_aw_valid; // @[Xbar.scala 258:23]
  assign _T_820 = _T_818 | reset; // @[Xbar.scala 258:12]
  assign _T_821 = ~_T_820; // @[Xbar.scala 258:12]
  assign _T_833 = ~out_2_ar_valid; // @[Xbar.scala 256:60]
  assign _T_839 = _T_833 | out_2_ar_valid; // @[Xbar.scala 258:23]
  assign _T_841 = _T_839 | reset; // @[Xbar.scala 258:12]
  assign _T_842 = ~_T_841; // @[Xbar.scala 258:12]
  assign _T_856 = ~out_3_aw_valid; // @[Xbar.scala 256:60]
  assign _T_862 = _T_856 | out_3_aw_valid; // @[Xbar.scala 258:23]
  assign _T_864 = _T_862 | reset; // @[Xbar.scala 258:12]
  assign _T_865 = ~_T_864; // @[Xbar.scala 258:12]
  assign _T_877 = ~out_3_ar_valid; // @[Xbar.scala 256:60]
  assign _T_883 = _T_877 | out_3_ar_valid; // @[Xbar.scala 258:23]
  assign _T_885 = _T_883 | reset; // @[Xbar.scala 258:12]
  assign _T_886 = ~_T_885; // @[Xbar.scala 258:12]
  assign _T_900 = ~out_4_aw_valid; // @[Xbar.scala 256:60]
  assign _T_906 = _T_900 | out_4_aw_valid; // @[Xbar.scala 258:23]
  assign _T_908 = _T_906 | reset; // @[Xbar.scala 258:12]
  assign _T_909 = ~_T_908; // @[Xbar.scala 258:12]
  assign _T_921 = ~out_4_ar_valid; // @[Xbar.scala 256:60]
  assign _T_927 = _T_921 | out_4_ar_valid; // @[Xbar.scala 258:23]
  assign _T_929 = _T_927 | reset; // @[Xbar.scala 258:12]
  assign _T_930 = ~_T_929; // @[Xbar.scala 258:12]
  assign _T_944 = ~out_5_aw_valid; // @[Xbar.scala 256:60]
  assign _T_950 = _T_944 | out_5_aw_valid; // @[Xbar.scala 258:23]
  assign _T_952 = _T_950 | reset; // @[Xbar.scala 258:12]
  assign _T_953 = ~_T_952; // @[Xbar.scala 258:12]
  assign _T_965 = ~out_5_ar_valid; // @[Xbar.scala 256:60]
  assign _T_971 = _T_965 | out_5_ar_valid; // @[Xbar.scala 258:23]
  assign _T_973 = _T_971 | reset; // @[Xbar.scala 258:12]
  assign _T_974 = ~_T_973; // @[Xbar.scala 258:12]
  assign _T_988 = ~out_6_aw_valid; // @[Xbar.scala 256:60]
  assign _T_994 = _T_988 | out_6_aw_valid; // @[Xbar.scala 258:23]
  assign _T_996 = _T_994 | reset; // @[Xbar.scala 258:12]
  assign _T_997 = ~_T_996; // @[Xbar.scala 258:12]
  assign _T_1009 = ~out_6_ar_valid; // @[Xbar.scala 256:60]
  assign _T_1015 = _T_1009 | out_6_ar_valid; // @[Xbar.scala 258:23]
  assign _T_1017 = _T_1015 | reset; // @[Xbar.scala 258:12]
  assign _T_1018 = ~_T_1017; // @[Xbar.scala 258:12]
  assign _T_1032 = ~out_7_aw_valid; // @[Xbar.scala 256:60]
  assign _T_1038 = _T_1032 | out_7_aw_valid; // @[Xbar.scala 258:23]
  assign _T_1040 = _T_1038 | reset; // @[Xbar.scala 258:12]
  assign _T_1041 = ~_T_1040; // @[Xbar.scala 258:12]
  assign _T_1053 = ~out_7_ar_valid; // @[Xbar.scala 256:60]
  assign _T_1059 = _T_1053 | out_7_ar_valid; // @[Xbar.scala 258:23]
  assign _T_1061 = _T_1059 | reset; // @[Xbar.scala 258:12]
  assign _T_1062 = ~_T_1061; // @[Xbar.scala 258:12]
  assign _T_1076 = ~out_8_aw_valid; // @[Xbar.scala 256:60]
  assign _T_1082 = _T_1076 | out_8_aw_valid; // @[Xbar.scala 258:23]
  assign _T_1084 = _T_1082 | reset; // @[Xbar.scala 258:12]
  assign _T_1085 = ~_T_1084; // @[Xbar.scala 258:12]
  assign _T_1097 = ~out_8_ar_valid; // @[Xbar.scala 256:60]
  assign _T_1103 = _T_1097 | out_8_ar_valid; // @[Xbar.scala 258:23]
  assign _T_1105 = _T_1103 | reset; // @[Xbar.scala 258:12]
  assign _T_1106 = ~_T_1105; // @[Xbar.scala 258:12]
  assign _T_1120 = ~out_9_aw_valid; // @[Xbar.scala 256:60]
  assign _T_1126 = _T_1120 | out_9_aw_valid; // @[Xbar.scala 258:23]
  assign _T_1128 = _T_1126 | reset; // @[Xbar.scala 258:12]
  assign _T_1129 = ~_T_1128; // @[Xbar.scala 258:12]
  assign _T_1141 = ~out_9_ar_valid; // @[Xbar.scala 256:60]
  assign _T_1147 = _T_1141 | out_9_ar_valid; // @[Xbar.scala 258:23]
  assign _T_1149 = _T_1147 | reset; // @[Xbar.scala 258:12]
  assign _T_1150 = ~_T_1149; // @[Xbar.scala 258:12]
  assign _T_1164 = ~out_10_aw_valid; // @[Xbar.scala 256:60]
  assign _T_1170 = _T_1164 | out_10_aw_valid; // @[Xbar.scala 258:23]
  assign _T_1172 = _T_1170 | reset; // @[Xbar.scala 258:12]
  assign _T_1173 = ~_T_1172; // @[Xbar.scala 258:12]
  assign _T_1185 = ~out_10_ar_valid; // @[Xbar.scala 256:60]
  assign _T_1191 = _T_1185 | out_10_ar_valid; // @[Xbar.scala 258:23]
  assign _T_1193 = _T_1191 | reset; // @[Xbar.scala 258:12]
  assign _T_1194 = ~_T_1193; // @[Xbar.scala 258:12]
  assign _T_1208 = ~out_11_aw_valid; // @[Xbar.scala 256:60]
  assign _T_1214 = _T_1208 | out_11_aw_valid; // @[Xbar.scala 258:23]
  assign _T_1216 = _T_1214 | reset; // @[Xbar.scala 258:12]
  assign _T_1217 = ~_T_1216; // @[Xbar.scala 258:12]
  assign _T_1229 = ~out_11_ar_valid; // @[Xbar.scala 256:60]
  assign _T_1235 = _T_1229 | out_11_ar_valid; // @[Xbar.scala 258:23]
  assign _T_1237 = _T_1235 | reset; // @[Xbar.scala 258:12]
  assign _T_1238 = ~_T_1237; // @[Xbar.scala 258:12]
  assign _T_1252 = ~out_12_aw_valid; // @[Xbar.scala 256:60]
  assign _T_1258 = _T_1252 | out_12_aw_valid; // @[Xbar.scala 258:23]
  assign _T_1260 = _T_1258 | reset; // @[Xbar.scala 258:12]
  assign _T_1261 = ~_T_1260; // @[Xbar.scala 258:12]
  assign _T_1273 = ~out_12_ar_valid; // @[Xbar.scala 256:60]
  assign _T_1279 = _T_1273 | out_12_ar_valid; // @[Xbar.scala 258:23]
  assign _T_1281 = _T_1279 | reset; // @[Xbar.scala 258:12]
  assign _T_1282 = ~_T_1281; // @[Xbar.scala 258:12]
  assign _T_1296 = ~out_13_aw_valid; // @[Xbar.scala 256:60]
  assign _T_1302 = _T_1296 | out_13_aw_valid; // @[Xbar.scala 258:23]
  assign _T_1304 = _T_1302 | reset; // @[Xbar.scala 258:12]
  assign _T_1305 = ~_T_1304; // @[Xbar.scala 258:12]
  assign _T_1317 = ~out_13_ar_valid; // @[Xbar.scala 256:60]
  assign _T_1323 = _T_1317 | out_13_ar_valid; // @[Xbar.scala 258:23]
  assign _T_1325 = _T_1323 | reset; // @[Xbar.scala 258:12]
  assign _T_1326 = ~_T_1325; // @[Xbar.scala 258:12]
  assign _T_1340 = ~out_14_aw_valid; // @[Xbar.scala 256:60]
  assign _T_1346 = _T_1340 | out_14_aw_valid; // @[Xbar.scala 258:23]
  assign _T_1348 = _T_1346 | reset; // @[Xbar.scala 258:12]
  assign _T_1349 = ~_T_1348; // @[Xbar.scala 258:12]
  assign _T_1361 = ~out_14_ar_valid; // @[Xbar.scala 256:60]
  assign _T_1367 = _T_1361 | out_14_ar_valid; // @[Xbar.scala 258:23]
  assign _T_1369 = _T_1367 | reset; // @[Xbar.scala 258:12]
  assign _T_1370 = ~_T_1369; // @[Xbar.scala 258:12]
  assign _T_1384 = ~out_15_aw_valid; // @[Xbar.scala 256:60]
  assign _T_1390 = _T_1384 | out_15_aw_valid; // @[Xbar.scala 258:23]
  assign _T_1392 = _T_1390 | reset; // @[Xbar.scala 258:12]
  assign _T_1393 = ~_T_1392; // @[Xbar.scala 258:12]
  assign _T_1405 = ~out_15_ar_valid; // @[Xbar.scala 256:60]
  assign _T_1411 = _T_1405 | out_15_ar_valid; // @[Xbar.scala 258:23]
  assign _T_1413 = _T_1411 | reset; // @[Xbar.scala 258:12]
  assign _T_1414 = ~_T_1413; // @[Xbar.scala 258:12]
  assign _T_1428 = ~out_16_aw_valid; // @[Xbar.scala 256:60]
  assign _T_1434 = _T_1428 | out_16_aw_valid; // @[Xbar.scala 258:23]
  assign _T_1436 = _T_1434 | reset; // @[Xbar.scala 258:12]
  assign _T_1437 = ~_T_1436; // @[Xbar.scala 258:12]
  assign _T_1449 = ~out_16_ar_valid; // @[Xbar.scala 256:60]
  assign _T_1455 = _T_1449 | out_16_ar_valid; // @[Xbar.scala 258:23]
  assign _T_1457 = _T_1455 | reset; // @[Xbar.scala 258:12]
  assign _T_1458 = ~_T_1457; // @[Xbar.scala 258:12]
  assign _T_1472 = ~out_17_aw_valid; // @[Xbar.scala 256:60]
  assign _T_1478 = _T_1472 | out_17_aw_valid; // @[Xbar.scala 258:23]
  assign _T_1480 = _T_1478 | reset; // @[Xbar.scala 258:12]
  assign _T_1481 = ~_T_1480; // @[Xbar.scala 258:12]
  assign _T_1493 = ~out_17_ar_valid; // @[Xbar.scala 256:60]
  assign _T_1499 = _T_1493 | out_17_ar_valid; // @[Xbar.scala 258:23]
  assign _T_1501 = _T_1499 | reset; // @[Xbar.scala 258:12]
  assign _T_1502 = ~_T_1501; // @[Xbar.scala 258:12]
  assign _T_1516 = ~out_18_aw_valid; // @[Xbar.scala 256:60]
  assign _T_1522 = _T_1516 | out_18_aw_valid; // @[Xbar.scala 258:23]
  assign _T_1524 = _T_1522 | reset; // @[Xbar.scala 258:12]
  assign _T_1525 = ~_T_1524; // @[Xbar.scala 258:12]
  assign _T_1537 = ~out_18_ar_valid; // @[Xbar.scala 256:60]
  assign _T_1543 = _T_1537 | out_18_ar_valid; // @[Xbar.scala 258:23]
  assign _T_1545 = _T_1543 | reset; // @[Xbar.scala 258:12]
  assign _T_1546 = ~_T_1545; // @[Xbar.scala 258:12]
  assign _T_1560 = ~out_19_aw_valid; // @[Xbar.scala 256:60]
  assign _T_1566 = _T_1560 | out_19_aw_valid; // @[Xbar.scala 258:23]
  assign _T_1568 = _T_1566 | reset; // @[Xbar.scala 258:12]
  assign _T_1569 = ~_T_1568; // @[Xbar.scala 258:12]
  assign _T_1581 = ~out_19_ar_valid; // @[Xbar.scala 256:60]
  assign _T_1587 = _T_1581 | out_19_ar_valid; // @[Xbar.scala 258:23]
  assign _T_1589 = _T_1587 | reset; // @[Xbar.scala 258:12]
  assign _T_1590 = ~_T_1589; // @[Xbar.scala 258:12]
  assign _T_1604 = ~out_20_aw_valid; // @[Xbar.scala 256:60]
  assign _T_1610 = _T_1604 | out_20_aw_valid; // @[Xbar.scala 258:23]
  assign _T_1612 = _T_1610 | reset; // @[Xbar.scala 258:12]
  assign _T_1613 = ~_T_1612; // @[Xbar.scala 258:12]
  assign _T_1625 = ~out_20_ar_valid; // @[Xbar.scala 256:60]
  assign _T_1631 = _T_1625 | out_20_ar_valid; // @[Xbar.scala 258:23]
  assign _T_1633 = _T_1631 | reset; // @[Xbar.scala 258:12]
  assign _T_1634 = ~_T_1633; // @[Xbar.scala 258:12]
  assign _T_1648 = ~out_21_aw_valid; // @[Xbar.scala 256:60]
  assign _T_1654 = _T_1648 | out_21_aw_valid; // @[Xbar.scala 258:23]
  assign _T_1656 = _T_1654 | reset; // @[Xbar.scala 258:12]
  assign _T_1657 = ~_T_1656; // @[Xbar.scala 258:12]
  assign _T_1669 = ~out_21_ar_valid; // @[Xbar.scala 256:60]
  assign _T_1675 = _T_1669 | out_21_ar_valid; // @[Xbar.scala 258:23]
  assign _T_1677 = _T_1675 | reset; // @[Xbar.scala 258:12]
  assign _T_1678 = ~_T_1677; // @[Xbar.scala 258:12]
  assign _T_1757 = _T_1728 != 22'h0; // @[Arbiter.scala 24:27]
  assign _T_1758 = _T_1686 & _T_1757; // @[Arbiter.scala 24:18]
  assign _T_1759 = _T_1756 & _T_1728; // @[Arbiter.scala 25:29]
  assign _T_1760 = {_T_1759, 1'h0}; // @[package.scala 199:48]
  assign _T_1762 = _T_1759 | _T_1760[21:0]; // @[package.scala 199:43]
  assign _T_1763 = {_T_1762, 2'h0}; // @[package.scala 199:48]
  assign _T_1765 = _T_1762 | _T_1763[21:0]; // @[package.scala 199:43]
  assign _T_1766 = {_T_1765, 4'h0}; // @[package.scala 199:48]
  assign _T_1768 = _T_1765 | _T_1766[21:0]; // @[package.scala 199:43]
  assign _T_1769 = {_T_1768, 8'h0}; // @[package.scala 199:48]
  assign _T_1771 = _T_1768 | _T_1769[21:0]; // @[package.scala 199:43]
  assign _T_1772 = {_T_1771, 16'h0}; // @[package.scala 199:48]
  assign _T_1774 = _T_1771 | _T_1772[21:0]; // @[package.scala 199:43]
  assign _T_1824 = _T_1800 | _T_1801; // @[Xbar.scala 255:50]
  assign _T_1825 = _T_1824 | _T_1802; // @[Xbar.scala 255:50]
  assign _T_1826 = _T_1825 | _T_1803; // @[Xbar.scala 255:50]
  assign _T_1827 = _T_1826 | _T_1804; // @[Xbar.scala 255:50]
  assign _T_1828 = _T_1827 | _T_1805; // @[Xbar.scala 255:50]
  assign _T_1829 = _T_1828 | _T_1806; // @[Xbar.scala 255:50]
  assign _T_1830 = _T_1829 | _T_1807; // @[Xbar.scala 255:50]
  assign _T_1831 = _T_1830 | _T_1808; // @[Xbar.scala 255:50]
  assign _T_1832 = _T_1831 | _T_1809; // @[Xbar.scala 255:50]
  assign _T_1833 = _T_1832 | _T_1810; // @[Xbar.scala 255:50]
  assign _T_1834 = _T_1833 | _T_1811; // @[Xbar.scala 255:50]
  assign _T_1835 = _T_1834 | _T_1812; // @[Xbar.scala 255:50]
  assign _T_1836 = _T_1835 | _T_1813; // @[Xbar.scala 255:50]
  assign _T_1837 = _T_1836 | _T_1814; // @[Xbar.scala 255:50]
  assign _T_1838 = _T_1837 | _T_1815; // @[Xbar.scala 255:50]
  assign _T_1839 = _T_1838 | _T_1816; // @[Xbar.scala 255:50]
  assign _T_1840 = _T_1839 | _T_1817; // @[Xbar.scala 255:50]
  assign _T_1841 = _T_1840 | _T_1818; // @[Xbar.scala 255:50]
  assign _T_1842 = _T_1841 | _T_1819; // @[Xbar.scala 255:50]
  assign _T_1843 = _T_1842 | _T_1820; // @[Xbar.scala 255:50]
  assign _T_1844 = _T_1843 | _T_1821; // @[Xbar.scala 255:50]
  assign _T_1846 = ~_T_1800; // @[Xbar.scala 256:60]
  assign _T_1849 = ~_T_1801; // @[Xbar.scala 256:60]
  assign _T_1850 = _T_1846 | _T_1849; // @[Xbar.scala 256:57]
  assign _T_1851 = ~_T_1824; // @[Xbar.scala 256:54]
  assign _T_1852 = ~_T_1802; // @[Xbar.scala 256:60]
  assign _T_1853 = _T_1851 | _T_1852; // @[Xbar.scala 256:57]
  assign _T_1854 = ~_T_1825; // @[Xbar.scala 256:54]
  assign _T_1855 = ~_T_1803; // @[Xbar.scala 256:60]
  assign _T_1856 = _T_1854 | _T_1855; // @[Xbar.scala 256:57]
  assign _T_1857 = ~_T_1826; // @[Xbar.scala 256:54]
  assign _T_1858 = ~_T_1804; // @[Xbar.scala 256:60]
  assign _T_1859 = _T_1857 | _T_1858; // @[Xbar.scala 256:57]
  assign _T_1860 = ~_T_1827; // @[Xbar.scala 256:54]
  assign _T_1861 = ~_T_1805; // @[Xbar.scala 256:60]
  assign _T_1862 = _T_1860 | _T_1861; // @[Xbar.scala 256:57]
  assign _T_1863 = ~_T_1828; // @[Xbar.scala 256:54]
  assign _T_1864 = ~_T_1806; // @[Xbar.scala 256:60]
  assign _T_1865 = _T_1863 | _T_1864; // @[Xbar.scala 256:57]
  assign _T_1866 = ~_T_1829; // @[Xbar.scala 256:54]
  assign _T_1867 = ~_T_1807; // @[Xbar.scala 256:60]
  assign _T_1868 = _T_1866 | _T_1867; // @[Xbar.scala 256:57]
  assign _T_1869 = ~_T_1830; // @[Xbar.scala 256:54]
  assign _T_1870 = ~_T_1808; // @[Xbar.scala 256:60]
  assign _T_1871 = _T_1869 | _T_1870; // @[Xbar.scala 256:57]
  assign _T_1872 = ~_T_1831; // @[Xbar.scala 256:54]
  assign _T_1873 = ~_T_1809; // @[Xbar.scala 256:60]
  assign _T_1874 = _T_1872 | _T_1873; // @[Xbar.scala 256:57]
  assign _T_1875 = ~_T_1832; // @[Xbar.scala 256:54]
  assign _T_1876 = ~_T_1810; // @[Xbar.scala 256:60]
  assign _T_1877 = _T_1875 | _T_1876; // @[Xbar.scala 256:57]
  assign _T_1878 = ~_T_1833; // @[Xbar.scala 256:54]
  assign _T_1879 = ~_T_1811; // @[Xbar.scala 256:60]
  assign _T_1880 = _T_1878 | _T_1879; // @[Xbar.scala 256:57]
  assign _T_1881 = ~_T_1834; // @[Xbar.scala 256:54]
  assign _T_1882 = ~_T_1812; // @[Xbar.scala 256:60]
  assign _T_1883 = _T_1881 | _T_1882; // @[Xbar.scala 256:57]
  assign _T_1884 = ~_T_1835; // @[Xbar.scala 256:54]
  assign _T_1885 = ~_T_1813; // @[Xbar.scala 256:60]
  assign _T_1886 = _T_1884 | _T_1885; // @[Xbar.scala 256:57]
  assign _T_1887 = ~_T_1836; // @[Xbar.scala 256:54]
  assign _T_1888 = ~_T_1814; // @[Xbar.scala 256:60]
  assign _T_1889 = _T_1887 | _T_1888; // @[Xbar.scala 256:57]
  assign _T_1890 = ~_T_1837; // @[Xbar.scala 256:54]
  assign _T_1891 = ~_T_1815; // @[Xbar.scala 256:60]
  assign _T_1892 = _T_1890 | _T_1891; // @[Xbar.scala 256:57]
  assign _T_1893 = ~_T_1838; // @[Xbar.scala 256:54]
  assign _T_1894 = ~_T_1816; // @[Xbar.scala 256:60]
  assign _T_1895 = _T_1893 | _T_1894; // @[Xbar.scala 256:57]
  assign _T_1896 = ~_T_1839; // @[Xbar.scala 256:54]
  assign _T_1897 = ~_T_1817; // @[Xbar.scala 256:60]
  assign _T_1898 = _T_1896 | _T_1897; // @[Xbar.scala 256:57]
  assign _T_1899 = ~_T_1840; // @[Xbar.scala 256:54]
  assign _T_1900 = ~_T_1818; // @[Xbar.scala 256:60]
  assign _T_1901 = _T_1899 | _T_1900; // @[Xbar.scala 256:57]
  assign _T_1902 = ~_T_1841; // @[Xbar.scala 256:54]
  assign _T_1903 = ~_T_1819; // @[Xbar.scala 256:60]
  assign _T_1904 = _T_1902 | _T_1903; // @[Xbar.scala 256:57]
  assign _T_1905 = ~_T_1842; // @[Xbar.scala 256:54]
  assign _T_1906 = ~_T_1820; // @[Xbar.scala 256:60]
  assign _T_1907 = _T_1905 | _T_1906; // @[Xbar.scala 256:57]
  assign _T_1908 = ~_T_1843; // @[Xbar.scala 256:54]
  assign _T_1909 = ~_T_1821; // @[Xbar.scala 256:60]
  assign _T_1910 = _T_1908 | _T_1909; // @[Xbar.scala 256:57]
  assign _T_1912 = _T_1850 & _T_1853; // @[Xbar.scala 256:75]
  assign _T_1913 = _T_1912 & _T_1856; // @[Xbar.scala 256:75]
  assign _T_1914 = _T_1913 & _T_1859; // @[Xbar.scala 256:75]
  assign _T_1915 = _T_1914 & _T_1862; // @[Xbar.scala 256:75]
  assign _T_1916 = _T_1915 & _T_1865; // @[Xbar.scala 256:75]
  assign _T_1917 = _T_1916 & _T_1868; // @[Xbar.scala 256:75]
  assign _T_1918 = _T_1917 & _T_1871; // @[Xbar.scala 256:75]
  assign _T_1919 = _T_1918 & _T_1874; // @[Xbar.scala 256:75]
  assign _T_1920 = _T_1919 & _T_1877; // @[Xbar.scala 256:75]
  assign _T_1921 = _T_1920 & _T_1880; // @[Xbar.scala 256:75]
  assign _T_1922 = _T_1921 & _T_1883; // @[Xbar.scala 256:75]
  assign _T_1923 = _T_1922 & _T_1886; // @[Xbar.scala 256:75]
  assign _T_1924 = _T_1923 & _T_1889; // @[Xbar.scala 256:75]
  assign _T_1925 = _T_1924 & _T_1892; // @[Xbar.scala 256:75]
  assign _T_1926 = _T_1925 & _T_1895; // @[Xbar.scala 256:75]
  assign _T_1927 = _T_1926 & _T_1898; // @[Xbar.scala 256:75]
  assign _T_1928 = _T_1927 & _T_1901; // @[Xbar.scala 256:75]
  assign _T_1929 = _T_1928 & _T_1904; // @[Xbar.scala 256:75]
  assign _T_1930 = _T_1929 & _T_1907; // @[Xbar.scala 256:75]
  assign _T_1931 = _T_1930 & _T_1910; // @[Xbar.scala 256:75]
  assign _T_1933 = _T_1931 | reset; // @[Xbar.scala 256:11]
  assign _T_1934 = ~_T_1933; // @[Xbar.scala 256:11]
  assign _T_1935 = ~_T_1707; // @[Xbar.scala 258:13]
  assign _T_1957 = _T_1935 | _T_1844; // @[Xbar.scala 258:23]
  assign _T_1959 = _T_1957 | reset; // @[Xbar.scala 258:12]
  assign _T_1960 = ~_T_1959; // @[Xbar.scala 258:12]
  assign _GEN_93 = _T_1707 ? 1'h0 : _T_1686; // @[Xbar.scala 266:21]
  assign _GEN_94 = _T_357 | _GEN_93; // @[Xbar.scala 267:24]
  assign _T_1965_0 = _T_1686 ? _T_1756[0] : _T_1962_0; // @[Xbar.scala 270:24]
  assign _T_1965_1 = _T_1686 ? _T_1756[1] : _T_1962_1; // @[Xbar.scala 270:24]
  assign _T_1965_2 = _T_1686 ? _T_1756[2] : _T_1962_2; // @[Xbar.scala 270:24]
  assign _T_1965_3 = _T_1686 ? _T_1756[3] : _T_1962_3; // @[Xbar.scala 270:24]
  assign _T_1965_4 = _T_1686 ? _T_1756[4] : _T_1962_4; // @[Xbar.scala 270:24]
  assign _T_1965_5 = _T_1686 ? _T_1756[5] : _T_1962_5; // @[Xbar.scala 270:24]
  assign _T_1965_6 = _T_1686 ? _T_1756[6] : _T_1962_6; // @[Xbar.scala 270:24]
  assign _T_1965_7 = _T_1686 ? _T_1756[7] : _T_1962_7; // @[Xbar.scala 270:24]
  assign _T_1965_8 = _T_1686 ? _T_1756[8] : _T_1962_8; // @[Xbar.scala 270:24]
  assign _T_1965_9 = _T_1686 ? _T_1756[9] : _T_1962_9; // @[Xbar.scala 270:24]
  assign _T_1965_10 = _T_1686 ? _T_1756[10] : _T_1962_10; // @[Xbar.scala 270:24]
  assign _T_1965_11 = _T_1686 ? _T_1756[11] : _T_1962_11; // @[Xbar.scala 270:24]
  assign _T_1965_12 = _T_1686 ? _T_1756[12] : _T_1962_12; // @[Xbar.scala 270:24]
  assign _T_1965_13 = _T_1686 ? _T_1756[13] : _T_1962_13; // @[Xbar.scala 270:24]
  assign _T_1965_14 = _T_1686 ? _T_1756[14] : _T_1962_14; // @[Xbar.scala 270:24]
  assign _T_1965_15 = _T_1686 ? _T_1756[15] : _T_1962_15; // @[Xbar.scala 270:24]
  assign _T_1965_16 = _T_1686 ? _T_1756[16] : _T_1962_16; // @[Xbar.scala 270:24]
  assign _T_1965_17 = _T_1686 ? _T_1756[17] : _T_1962_17; // @[Xbar.scala 270:24]
  assign _T_1965_18 = _T_1686 ? _T_1756[18] : _T_1962_18; // @[Xbar.scala 270:24]
  assign _T_1965_19 = _T_1686 ? _T_1756[19] : _T_1962_19; // @[Xbar.scala 270:24]
  assign _T_1965_20 = _T_1686 ? _T_1756[20] : _T_1962_20; // @[Xbar.scala 270:24]
  assign _T_1965_21 = _T_1686 ? _T_1756[21] : _T_1962_21; // @[Xbar.scala 270:24]
  assign _T_2173 = {_T_683,_T_681,_T_679,_T_677,_T_675}; // @[Cat.scala 29:58]
  assign _T_2179 = {_T_695,_T_693,_T_691,_T_689,_T_687,_T_685,_T_2173}; // @[Cat.scala 29:58]
  assign _T_2183 = {_T_705,_T_703,_T_701,_T_699,_T_697}; // @[Cat.scala 29:58]
  assign _T_2190 = {auto_out_21_b_valid,_T_715,_T_713,_T_711,_T_709,_T_707,_T_2183,_T_2179}; // @[Cat.scala 29:58]
  assign _T_2198 = ~_T_2197; // @[Arbiter.scala 21:30]
  assign _T_2199 = _T_2190 & _T_2198; // @[Arbiter.scala 21:28]
  assign _T_2200 = {_T_2199,auto_out_21_b_valid,_T_715,_T_713,_T_711,_T_709,_T_707,_T_2183,_T_2179}; // @[Cat.scala 29:58]
  assign _GEN_110 = {{1'd0}, _T_2200[43:1]}; // @[package.scala 208:43]
  assign _T_2202 = _T_2200 | _GEN_110; // @[package.scala 208:43]
  assign _GEN_111 = {{2'd0}, _T_2202[43:2]}; // @[package.scala 208:43]
  assign _T_2204 = _T_2202 | _GEN_111; // @[package.scala 208:43]
  assign _GEN_112 = {{4'd0}, _T_2204[43:4]}; // @[package.scala 208:43]
  assign _T_2206 = _T_2204 | _GEN_112; // @[package.scala 208:43]
  assign _GEN_113 = {{8'd0}, _T_2206[43:8]}; // @[package.scala 208:43]
  assign _T_2208 = _T_2206 | _GEN_113; // @[package.scala 208:43]
  assign _GEN_114 = {{16'd0}, _T_2208[43:16]}; // @[package.scala 208:43]
  assign _T_2210 = _T_2208 | _GEN_114; // @[package.scala 208:43]
  assign _T_2213 = {_T_2197, 22'h0}; // @[Arbiter.scala 22:66]
  assign _GEN_115 = {{1'd0}, _T_2210[43:1]}; // @[Arbiter.scala 22:58]
  assign _T_2214 = _GEN_115 | _T_2213; // @[Arbiter.scala 22:58]
  assign _T_2217 = _T_2214[43:22] & _T_2214[21:0]; // @[Arbiter.scala 23:39]
  assign _T_2218 = ~_T_2217; // @[Arbiter.scala 23:18]
  assign _T_2219 = _T_2190 != 22'h0; // @[Arbiter.scala 24:27]
  assign _T_2220 = _T_2148 & _T_2219; // @[Arbiter.scala 24:18]
  assign _T_2221 = _T_2218 & _T_2190; // @[Arbiter.scala 25:29]
  assign _T_2222 = {_T_2221, 1'h0}; // @[package.scala 199:48]
  assign _T_2224 = _T_2221 | _T_2222[21:0]; // @[package.scala 199:43]
  assign _T_2225 = {_T_2224, 2'h0}; // @[package.scala 199:48]
  assign _T_2227 = _T_2224 | _T_2225[21:0]; // @[package.scala 199:43]
  assign _T_2228 = {_T_2227, 4'h0}; // @[package.scala 199:48]
  assign _T_2230 = _T_2227 | _T_2228[21:0]; // @[package.scala 199:43]
  assign _T_2231 = {_T_2230, 8'h0}; // @[package.scala 199:48]
  assign _T_2233 = _T_2230 | _T_2231[21:0]; // @[package.scala 199:43]
  assign _T_2234 = {_T_2233, 16'h0}; // @[package.scala 199:48]
  assign _T_2236 = _T_2233 | _T_2234[21:0]; // @[package.scala 199:43]
  assign _T_2262 = _T_2218[0] & _T_675; // @[Xbar.scala 250:63]
  assign _T_2263 = _T_2218[1] & _T_677; // @[Xbar.scala 250:63]
  assign _T_2264 = _T_2218[2] & _T_679; // @[Xbar.scala 250:63]
  assign _T_2265 = _T_2218[3] & _T_681; // @[Xbar.scala 250:63]
  assign _T_2266 = _T_2218[4] & _T_683; // @[Xbar.scala 250:63]
  assign _T_2267 = _T_2218[5] & _T_685; // @[Xbar.scala 250:63]
  assign _T_2268 = _T_2218[6] & _T_687; // @[Xbar.scala 250:63]
  assign _T_2269 = _T_2218[7] & _T_689; // @[Xbar.scala 250:63]
  assign _T_2270 = _T_2218[8] & _T_691; // @[Xbar.scala 250:63]
  assign _T_2271 = _T_2218[9] & _T_693; // @[Xbar.scala 250:63]
  assign _T_2272 = _T_2218[10] & _T_695; // @[Xbar.scala 250:63]
  assign _T_2273 = _T_2218[11] & _T_697; // @[Xbar.scala 250:63]
  assign _T_2274 = _T_2218[12] & _T_699; // @[Xbar.scala 250:63]
  assign _T_2275 = _T_2218[13] & _T_701; // @[Xbar.scala 250:63]
  assign _T_2276 = _T_2218[14] & _T_703; // @[Xbar.scala 250:63]
  assign _T_2277 = _T_2218[15] & _T_705; // @[Xbar.scala 250:63]
  assign _T_2278 = _T_2218[16] & _T_707; // @[Xbar.scala 250:63]
  assign _T_2279 = _T_2218[17] & _T_709; // @[Xbar.scala 250:63]
  assign _T_2280 = _T_2218[18] & _T_711; // @[Xbar.scala 250:63]
  assign _T_2281 = _T_2218[19] & _T_713; // @[Xbar.scala 250:63]
  assign _T_2282 = _T_2218[20] & _T_715; // @[Xbar.scala 250:63]
  assign _T_2283 = _T_2218[21] & auto_out_21_b_valid; // @[Xbar.scala 250:63]
  assign _T_2286 = _T_2262 | _T_2263; // @[Xbar.scala 255:50]
  assign _T_2287 = _T_2286 | _T_2264; // @[Xbar.scala 255:50]
  assign _T_2288 = _T_2287 | _T_2265; // @[Xbar.scala 255:50]
  assign _T_2289 = _T_2288 | _T_2266; // @[Xbar.scala 255:50]
  assign _T_2290 = _T_2289 | _T_2267; // @[Xbar.scala 255:50]
  assign _T_2291 = _T_2290 | _T_2268; // @[Xbar.scala 255:50]
  assign _T_2292 = _T_2291 | _T_2269; // @[Xbar.scala 255:50]
  assign _T_2293 = _T_2292 | _T_2270; // @[Xbar.scala 255:50]
  assign _T_2294 = _T_2293 | _T_2271; // @[Xbar.scala 255:50]
  assign _T_2295 = _T_2294 | _T_2272; // @[Xbar.scala 255:50]
  assign _T_2296 = _T_2295 | _T_2273; // @[Xbar.scala 255:50]
  assign _T_2297 = _T_2296 | _T_2274; // @[Xbar.scala 255:50]
  assign _T_2298 = _T_2297 | _T_2275; // @[Xbar.scala 255:50]
  assign _T_2299 = _T_2298 | _T_2276; // @[Xbar.scala 255:50]
  assign _T_2300 = _T_2299 | _T_2277; // @[Xbar.scala 255:50]
  assign _T_2301 = _T_2300 | _T_2278; // @[Xbar.scala 255:50]
  assign _T_2302 = _T_2301 | _T_2279; // @[Xbar.scala 255:50]
  assign _T_2303 = _T_2302 | _T_2280; // @[Xbar.scala 255:50]
  assign _T_2304 = _T_2303 | _T_2281; // @[Xbar.scala 255:50]
  assign _T_2305 = _T_2304 | _T_2282; // @[Xbar.scala 255:50]
  assign _T_2306 = _T_2305 | _T_2283; // @[Xbar.scala 255:50]
  assign _T_2308 = ~_T_2262; // @[Xbar.scala 256:60]
  assign _T_2311 = ~_T_2263; // @[Xbar.scala 256:60]
  assign _T_2312 = _T_2308 | _T_2311; // @[Xbar.scala 256:57]
  assign _T_2313 = ~_T_2286; // @[Xbar.scala 256:54]
  assign _T_2314 = ~_T_2264; // @[Xbar.scala 256:60]
  assign _T_2315 = _T_2313 | _T_2314; // @[Xbar.scala 256:57]
  assign _T_2316 = ~_T_2287; // @[Xbar.scala 256:54]
  assign _T_2317 = ~_T_2265; // @[Xbar.scala 256:60]
  assign _T_2318 = _T_2316 | _T_2317; // @[Xbar.scala 256:57]
  assign _T_2319 = ~_T_2288; // @[Xbar.scala 256:54]
  assign _T_2320 = ~_T_2266; // @[Xbar.scala 256:60]
  assign _T_2321 = _T_2319 | _T_2320; // @[Xbar.scala 256:57]
  assign _T_2322 = ~_T_2289; // @[Xbar.scala 256:54]
  assign _T_2323 = ~_T_2267; // @[Xbar.scala 256:60]
  assign _T_2324 = _T_2322 | _T_2323; // @[Xbar.scala 256:57]
  assign _T_2325 = ~_T_2290; // @[Xbar.scala 256:54]
  assign _T_2326 = ~_T_2268; // @[Xbar.scala 256:60]
  assign _T_2327 = _T_2325 | _T_2326; // @[Xbar.scala 256:57]
  assign _T_2328 = ~_T_2291; // @[Xbar.scala 256:54]
  assign _T_2329 = ~_T_2269; // @[Xbar.scala 256:60]
  assign _T_2330 = _T_2328 | _T_2329; // @[Xbar.scala 256:57]
  assign _T_2331 = ~_T_2292; // @[Xbar.scala 256:54]
  assign _T_2332 = ~_T_2270; // @[Xbar.scala 256:60]
  assign _T_2333 = _T_2331 | _T_2332; // @[Xbar.scala 256:57]
  assign _T_2334 = ~_T_2293; // @[Xbar.scala 256:54]
  assign _T_2335 = ~_T_2271; // @[Xbar.scala 256:60]
  assign _T_2336 = _T_2334 | _T_2335; // @[Xbar.scala 256:57]
  assign _T_2337 = ~_T_2294; // @[Xbar.scala 256:54]
  assign _T_2338 = ~_T_2272; // @[Xbar.scala 256:60]
  assign _T_2339 = _T_2337 | _T_2338; // @[Xbar.scala 256:57]
  assign _T_2340 = ~_T_2295; // @[Xbar.scala 256:54]
  assign _T_2341 = ~_T_2273; // @[Xbar.scala 256:60]
  assign _T_2342 = _T_2340 | _T_2341; // @[Xbar.scala 256:57]
  assign _T_2343 = ~_T_2296; // @[Xbar.scala 256:54]
  assign _T_2344 = ~_T_2274; // @[Xbar.scala 256:60]
  assign _T_2345 = _T_2343 | _T_2344; // @[Xbar.scala 256:57]
  assign _T_2346 = ~_T_2297; // @[Xbar.scala 256:54]
  assign _T_2347 = ~_T_2275; // @[Xbar.scala 256:60]
  assign _T_2348 = _T_2346 | _T_2347; // @[Xbar.scala 256:57]
  assign _T_2349 = ~_T_2298; // @[Xbar.scala 256:54]
  assign _T_2350 = ~_T_2276; // @[Xbar.scala 256:60]
  assign _T_2351 = _T_2349 | _T_2350; // @[Xbar.scala 256:57]
  assign _T_2352 = ~_T_2299; // @[Xbar.scala 256:54]
  assign _T_2353 = ~_T_2277; // @[Xbar.scala 256:60]
  assign _T_2354 = _T_2352 | _T_2353; // @[Xbar.scala 256:57]
  assign _T_2355 = ~_T_2300; // @[Xbar.scala 256:54]
  assign _T_2356 = ~_T_2278; // @[Xbar.scala 256:60]
  assign _T_2357 = _T_2355 | _T_2356; // @[Xbar.scala 256:57]
  assign _T_2358 = ~_T_2301; // @[Xbar.scala 256:54]
  assign _T_2359 = ~_T_2279; // @[Xbar.scala 256:60]
  assign _T_2360 = _T_2358 | _T_2359; // @[Xbar.scala 256:57]
  assign _T_2361 = ~_T_2302; // @[Xbar.scala 256:54]
  assign _T_2362 = ~_T_2280; // @[Xbar.scala 256:60]
  assign _T_2363 = _T_2361 | _T_2362; // @[Xbar.scala 256:57]
  assign _T_2364 = ~_T_2303; // @[Xbar.scala 256:54]
  assign _T_2365 = ~_T_2281; // @[Xbar.scala 256:60]
  assign _T_2366 = _T_2364 | _T_2365; // @[Xbar.scala 256:57]
  assign _T_2367 = ~_T_2304; // @[Xbar.scala 256:54]
  assign _T_2368 = ~_T_2282; // @[Xbar.scala 256:60]
  assign _T_2369 = _T_2367 | _T_2368; // @[Xbar.scala 256:57]
  assign _T_2370 = ~_T_2305; // @[Xbar.scala 256:54]
  assign _T_2371 = ~_T_2283; // @[Xbar.scala 256:60]
  assign _T_2372 = _T_2370 | _T_2371; // @[Xbar.scala 256:57]
  assign _T_2374 = _T_2312 & _T_2315; // @[Xbar.scala 256:75]
  assign _T_2375 = _T_2374 & _T_2318; // @[Xbar.scala 256:75]
  assign _T_2376 = _T_2375 & _T_2321; // @[Xbar.scala 256:75]
  assign _T_2377 = _T_2376 & _T_2324; // @[Xbar.scala 256:75]
  assign _T_2378 = _T_2377 & _T_2327; // @[Xbar.scala 256:75]
  assign _T_2379 = _T_2378 & _T_2330; // @[Xbar.scala 256:75]
  assign _T_2380 = _T_2379 & _T_2333; // @[Xbar.scala 256:75]
  assign _T_2381 = _T_2380 & _T_2336; // @[Xbar.scala 256:75]
  assign _T_2382 = _T_2381 & _T_2339; // @[Xbar.scala 256:75]
  assign _T_2383 = _T_2382 & _T_2342; // @[Xbar.scala 256:75]
  assign _T_2384 = _T_2383 & _T_2345; // @[Xbar.scala 256:75]
  assign _T_2385 = _T_2384 & _T_2348; // @[Xbar.scala 256:75]
  assign _T_2386 = _T_2385 & _T_2351; // @[Xbar.scala 256:75]
  assign _T_2387 = _T_2386 & _T_2354; // @[Xbar.scala 256:75]
  assign _T_2388 = _T_2387 & _T_2357; // @[Xbar.scala 256:75]
  assign _T_2389 = _T_2388 & _T_2360; // @[Xbar.scala 256:75]
  assign _T_2390 = _T_2389 & _T_2363; // @[Xbar.scala 256:75]
  assign _T_2391 = _T_2390 & _T_2366; // @[Xbar.scala 256:75]
  assign _T_2392 = _T_2391 & _T_2369; // @[Xbar.scala 256:75]
  assign _T_2393 = _T_2392 & _T_2372; // @[Xbar.scala 256:75]
  assign _T_2395 = _T_2393 | reset; // @[Xbar.scala 256:11]
  assign _T_2396 = ~_T_2395; // @[Xbar.scala 256:11]
  assign _T_2397 = ~_T_2169; // @[Xbar.scala 258:13]
  assign _T_2419 = _T_2397 | _T_2306; // @[Xbar.scala 258:23]
  assign _T_2421 = _T_2419 | reset; // @[Xbar.scala 258:12]
  assign _T_2422 = ~_T_2421; // @[Xbar.scala 258:12]
  assign _T_2425_0 = _T_2148 ? _T_2262 : _T_2424_0; // @[Xbar.scala 262:23]
  assign _T_2425_1 = _T_2148 ? _T_2263 : _T_2424_1; // @[Xbar.scala 262:23]
  assign _T_2425_2 = _T_2148 ? _T_2264 : _T_2424_2; // @[Xbar.scala 262:23]
  assign _T_2425_3 = _T_2148 ? _T_2265 : _T_2424_3; // @[Xbar.scala 262:23]
  assign _T_2425_4 = _T_2148 ? _T_2266 : _T_2424_4; // @[Xbar.scala 262:23]
  assign _T_2425_5 = _T_2148 ? _T_2267 : _T_2424_5; // @[Xbar.scala 262:23]
  assign _T_2425_6 = _T_2148 ? _T_2268 : _T_2424_6; // @[Xbar.scala 262:23]
  assign _T_2425_7 = _T_2148 ? _T_2269 : _T_2424_7; // @[Xbar.scala 262:23]
  assign _T_2425_8 = _T_2148 ? _T_2270 : _T_2424_8; // @[Xbar.scala 262:23]
  assign _T_2425_9 = _T_2148 ? _T_2271 : _T_2424_9; // @[Xbar.scala 262:23]
  assign _T_2425_10 = _T_2148 ? _T_2272 : _T_2424_10; // @[Xbar.scala 262:23]
  assign _T_2425_11 = _T_2148 ? _T_2273 : _T_2424_11; // @[Xbar.scala 262:23]
  assign _T_2425_12 = _T_2148 ? _T_2274 : _T_2424_12; // @[Xbar.scala 262:23]
  assign _T_2425_13 = _T_2148 ? _T_2275 : _T_2424_13; // @[Xbar.scala 262:23]
  assign _T_2425_14 = _T_2148 ? _T_2276 : _T_2424_14; // @[Xbar.scala 262:23]
  assign _T_2425_15 = _T_2148 ? _T_2277 : _T_2424_15; // @[Xbar.scala 262:23]
  assign _T_2425_16 = _T_2148 ? _T_2278 : _T_2424_16; // @[Xbar.scala 262:23]
  assign _T_2425_17 = _T_2148 ? _T_2279 : _T_2424_17; // @[Xbar.scala 262:23]
  assign _T_2425_18 = _T_2148 ? _T_2280 : _T_2424_18; // @[Xbar.scala 262:23]
  assign _T_2425_19 = _T_2148 ? _T_2281 : _T_2424_19; // @[Xbar.scala 262:23]
  assign _T_2425_20 = _T_2148 ? _T_2282 : _T_2424_20; // @[Xbar.scala 262:23]
  assign _T_2425_21 = _T_2148 ? _T_2283 : _T_2424_21; // @[Xbar.scala 262:23]
  assign _GEN_96 = _T_2169 ? 1'h0 : _T_2148; // @[Xbar.scala 266:21]
  assign _GEN_97 = _T_386 | _GEN_96; // @[Xbar.scala 267:24]
  assign _T_2427_0 = _T_2148 ? _T_2218[0] : _T_2424_0; // @[Xbar.scala 270:24]
  assign _T_2427_1 = _T_2148 ? _T_2218[1] : _T_2424_1; // @[Xbar.scala 270:24]
  assign _T_2427_2 = _T_2148 ? _T_2218[2] : _T_2424_2; // @[Xbar.scala 270:24]
  assign _T_2427_3 = _T_2148 ? _T_2218[3] : _T_2424_3; // @[Xbar.scala 270:24]
  assign _T_2427_4 = _T_2148 ? _T_2218[4] : _T_2424_4; // @[Xbar.scala 270:24]
  assign _T_2427_5 = _T_2148 ? _T_2218[5] : _T_2424_5; // @[Xbar.scala 270:24]
  assign _T_2427_6 = _T_2148 ? _T_2218[6] : _T_2424_6; // @[Xbar.scala 270:24]
  assign _T_2427_7 = _T_2148 ? _T_2218[7] : _T_2424_7; // @[Xbar.scala 270:24]
  assign _T_2427_8 = _T_2148 ? _T_2218[8] : _T_2424_8; // @[Xbar.scala 270:24]
  assign _T_2427_9 = _T_2148 ? _T_2218[9] : _T_2424_9; // @[Xbar.scala 270:24]
  assign _T_2427_10 = _T_2148 ? _T_2218[10] : _T_2424_10; // @[Xbar.scala 270:24]
  assign _T_2427_11 = _T_2148 ? _T_2218[11] : _T_2424_11; // @[Xbar.scala 270:24]
  assign _T_2427_12 = _T_2148 ? _T_2218[12] : _T_2424_12; // @[Xbar.scala 270:24]
  assign _T_2427_13 = _T_2148 ? _T_2218[13] : _T_2424_13; // @[Xbar.scala 270:24]
  assign _T_2427_14 = _T_2148 ? _T_2218[14] : _T_2424_14; // @[Xbar.scala 270:24]
  assign _T_2427_15 = _T_2148 ? _T_2218[15] : _T_2424_15; // @[Xbar.scala 270:24]
  assign _T_2427_16 = _T_2148 ? _T_2218[16] : _T_2424_16; // @[Xbar.scala 270:24]
  assign _T_2427_17 = _T_2148 ? _T_2218[17] : _T_2424_17; // @[Xbar.scala 270:24]
  assign _T_2427_18 = _T_2148 ? _T_2218[18] : _T_2424_18; // @[Xbar.scala 270:24]
  assign _T_2427_19 = _T_2148 ? _T_2218[19] : _T_2424_19; // @[Xbar.scala 270:24]
  assign _T_2427_20 = _T_2148 ? _T_2218[20] : _T_2424_20; // @[Xbar.scala 270:24]
  assign _T_2427_21 = _T_2148 ? _T_2218[21] : _T_2424_21; // @[Xbar.scala 270:24]
  assign _T_2495 = {auto_out_0_b_bits_id,auto_out_0_b_bits_resp}; // @[Mux.scala 27:72]
  assign _T_2496 = _T_2425_0 ? _T_2495 : 3'h0; // @[Mux.scala 27:72]
  assign _T_2497 = {auto_out_1_b_bits_id,auto_out_1_b_bits_resp}; // @[Mux.scala 27:72]
  assign _T_2498 = _T_2425_1 ? _T_2497 : 3'h0; // @[Mux.scala 27:72]
  assign _T_2499 = {auto_out_2_b_bits_id,auto_out_2_b_bits_resp}; // @[Mux.scala 27:72]
  assign _T_2500 = _T_2425_2 ? _T_2499 : 3'h0; // @[Mux.scala 27:72]
  assign _T_2501 = {auto_out_3_b_bits_id,auto_out_3_b_bits_resp}; // @[Mux.scala 27:72]
  assign _T_2502 = _T_2425_3 ? _T_2501 : 3'h0; // @[Mux.scala 27:72]
  assign _T_2503 = {auto_out_4_b_bits_id,auto_out_4_b_bits_resp}; // @[Mux.scala 27:72]
  assign _T_2504 = _T_2425_4 ? _T_2503 : 3'h0; // @[Mux.scala 27:72]
  assign _T_2505 = {auto_out_5_b_bits_id,auto_out_5_b_bits_resp}; // @[Mux.scala 27:72]
  assign _T_2506 = _T_2425_5 ? _T_2505 : 3'h0; // @[Mux.scala 27:72]
  assign _T_2507 = {auto_out_6_b_bits_id,auto_out_6_b_bits_resp}; // @[Mux.scala 27:72]
  assign _T_2508 = _T_2425_6 ? _T_2507 : 3'h0; // @[Mux.scala 27:72]
  assign _T_2509 = {auto_out_7_b_bits_id,auto_out_7_b_bits_resp}; // @[Mux.scala 27:72]
  assign _T_2510 = _T_2425_7 ? _T_2509 : 3'h0; // @[Mux.scala 27:72]
  assign _T_2511 = {auto_out_8_b_bits_id,auto_out_8_b_bits_resp}; // @[Mux.scala 27:72]
  assign _T_2512 = _T_2425_8 ? _T_2511 : 3'h0; // @[Mux.scala 27:72]
  assign _T_2513 = {auto_out_9_b_bits_id,auto_out_9_b_bits_resp}; // @[Mux.scala 27:72]
  assign _T_2514 = _T_2425_9 ? _T_2513 : 3'h0; // @[Mux.scala 27:72]
  assign _T_2515 = {auto_out_10_b_bits_id,auto_out_10_b_bits_resp}; // @[Mux.scala 27:72]
  assign _T_2516 = _T_2425_10 ? _T_2515 : 3'h0; // @[Mux.scala 27:72]
  assign _T_2517 = {auto_out_11_b_bits_id,auto_out_11_b_bits_resp}; // @[Mux.scala 27:72]
  assign _T_2518 = _T_2425_11 ? _T_2517 : 3'h0; // @[Mux.scala 27:72]
  assign _T_2519 = {auto_out_12_b_bits_id,auto_out_12_b_bits_resp}; // @[Mux.scala 27:72]
  assign _T_2520 = _T_2425_12 ? _T_2519 : 3'h0; // @[Mux.scala 27:72]
  assign _T_2521 = {auto_out_13_b_bits_id,auto_out_13_b_bits_resp}; // @[Mux.scala 27:72]
  assign _T_2522 = _T_2425_13 ? _T_2521 : 3'h0; // @[Mux.scala 27:72]
  assign _T_2523 = {auto_out_14_b_bits_id,auto_out_14_b_bits_resp}; // @[Mux.scala 27:72]
  assign _T_2524 = _T_2425_14 ? _T_2523 : 3'h0; // @[Mux.scala 27:72]
  assign _T_2525 = {auto_out_15_b_bits_id,auto_out_15_b_bits_resp}; // @[Mux.scala 27:72]
  assign _T_2526 = _T_2425_15 ? _T_2525 : 3'h0; // @[Mux.scala 27:72]
  assign _T_2527 = {auto_out_16_b_bits_id,auto_out_16_b_bits_resp}; // @[Mux.scala 27:72]
  assign _T_2528 = _T_2425_16 ? _T_2527 : 3'h0; // @[Mux.scala 27:72]
  assign _T_2529 = {auto_out_17_b_bits_id,auto_out_17_b_bits_resp}; // @[Mux.scala 27:72]
  assign _T_2530 = _T_2425_17 ? _T_2529 : 3'h0; // @[Mux.scala 27:72]
  assign _T_2531 = {auto_out_18_b_bits_id,auto_out_18_b_bits_resp}; // @[Mux.scala 27:72]
  assign _T_2532 = _T_2425_18 ? _T_2531 : 3'h0; // @[Mux.scala 27:72]
  assign _T_2533 = {auto_out_19_b_bits_id,auto_out_19_b_bits_resp}; // @[Mux.scala 27:72]
  assign _T_2534 = _T_2425_19 ? _T_2533 : 3'h0; // @[Mux.scala 27:72]
  assign _T_2535 = {auto_out_20_b_bits_id,auto_out_20_b_bits_resp}; // @[Mux.scala 27:72]
  assign _T_2536 = _T_2425_20 ? _T_2535 : 3'h0; // @[Mux.scala 27:72]
  assign _T_2537 = {1'h0,auto_out_21_b_bits_resp}; // @[Mux.scala 27:72]
  assign _T_2538 = _T_2425_21 ? _T_2537 : 3'h0; // @[Mux.scala 27:72]
  assign _T_2539 = _T_2496 | _T_2498; // @[Mux.scala 27:72]
  assign _T_2540 = _T_2539 | _T_2500; // @[Mux.scala 27:72]
  assign _T_2541 = _T_2540 | _T_2502; // @[Mux.scala 27:72]
  assign _T_2542 = _T_2541 | _T_2504; // @[Mux.scala 27:72]
  assign _T_2543 = _T_2542 | _T_2506; // @[Mux.scala 27:72]
  assign _T_2544 = _T_2543 | _T_2508; // @[Mux.scala 27:72]
  assign _T_2545 = _T_2544 | _T_2510; // @[Mux.scala 27:72]
  assign _T_2546 = _T_2545 | _T_2512; // @[Mux.scala 27:72]
  assign _T_2547 = _T_2546 | _T_2514; // @[Mux.scala 27:72]
  assign _T_2548 = _T_2547 | _T_2516; // @[Mux.scala 27:72]
  assign _T_2549 = _T_2548 | _T_2518; // @[Mux.scala 27:72]
  assign _T_2550 = _T_2549 | _T_2520; // @[Mux.scala 27:72]
  assign _T_2551 = _T_2550 | _T_2522; // @[Mux.scala 27:72]
  assign _T_2552 = _T_2551 | _T_2524; // @[Mux.scala 27:72]
  assign _T_2553 = _T_2552 | _T_2526; // @[Mux.scala 27:72]
  assign _T_2554 = _T_2553 | _T_2528; // @[Mux.scala 27:72]
  assign _T_2555 = _T_2554 | _T_2530; // @[Mux.scala 27:72]
  assign _T_2556 = _T_2555 | _T_2532; // @[Mux.scala 27:72]
  assign _T_2557 = _T_2556 | _T_2534; // @[Mux.scala 27:72]
  assign _T_2558 = _T_2557 | _T_2536; // @[Mux.scala 27:72]
  assign _T_2559 = _T_2558 | _T_2538; // @[Mux.scala 27:72]
  assign auto_in_aw_ready = _T_419 & _T_411; // @[LazyModule.scala 173:31]
  assign auto_in_w_ready = in_0_w_ready & awIn_0_io_deq_valid; // @[LazyModule.scala 173:31]
  assign auto_in_b_valid = _T_2148 ? _T_2169 : _T_2492; // @[LazyModule.scala 173:31]
  assign auto_in_b_bits_resp = _T_2559[1:0]; // @[LazyModule.scala 173:31]
  assign auto_in_ar_ready = in_0_ar_ready & _T_383; // @[LazyModule.scala 173:31]
  assign auto_in_r_valid = _T_1686 ? _T_1707 : _T_2030; // @[LazyModule.scala 173:31]
  assign auto_in_r_bits_data = _T_2141[34:3]; // @[LazyModule.scala 173:31]
  assign auto_in_r_bits_resp = _T_2141[2:1]; // @[LazyModule.scala 173:31]
  assign auto_in_r_bits_last = _T_2141[0]; // @[LazyModule.scala 173:31]
  assign auto_out_21_aw_valid = in_0_aw_valid & requestAWIO_0_21; // @[LazyModule.scala 173:49]
  assign auto_out_21_aw_bits_id = auto_in_aw_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_21_aw_bits_addr = auto_in_aw_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_21_aw_bits_size = auto_in_aw_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_21_w_valid = in_0_w_valid & requestWIO_0_21; // @[LazyModule.scala 173:49]
  assign auto_out_21_w_bits_data = auto_in_w_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_21_w_bits_strb = auto_in_w_bits_strb; // @[LazyModule.scala 173:49]
  assign auto_out_21_w_bits_last = auto_in_w_bits_last; // @[LazyModule.scala 173:49]
  assign auto_out_21_b_ready = auto_in_b_ready & _T_2427_21; // @[LazyModule.scala 173:49]
  assign auto_out_21_ar_valid = in_0_ar_valid & requestARIO_0_21; // @[LazyModule.scala 173:49]
  assign auto_out_21_ar_bits_id = auto_in_ar_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_21_ar_bits_addr = auto_in_ar_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_21_ar_bits_size = auto_in_ar_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_21_r_ready = auto_in_r_ready & _T_1965_21; // @[LazyModule.scala 173:49]
  assign auto_out_20_aw_valid = in_0_aw_valid & requestAWIO_0_20; // @[LazyModule.scala 173:49]
  assign auto_out_20_aw_bits_id = auto_in_aw_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_20_aw_bits_addr = auto_in_aw_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_20_aw_bits_size = auto_in_aw_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_20_w_valid = in_0_w_valid & requestWIO_0_20; // @[LazyModule.scala 173:49]
  assign auto_out_20_w_bits_data = auto_in_w_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_20_w_bits_strb = auto_in_w_bits_strb; // @[LazyModule.scala 173:49]
  assign auto_out_20_w_bits_last = auto_in_w_bits_last; // @[LazyModule.scala 173:49]
  assign auto_out_20_b_ready = auto_in_b_ready & _T_2427_20; // @[LazyModule.scala 173:49]
  assign auto_out_20_ar_valid = in_0_ar_valid & requestARIO_0_20; // @[LazyModule.scala 173:49]
  assign auto_out_20_ar_bits_id = auto_in_ar_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_20_ar_bits_addr = auto_in_ar_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_20_ar_bits_size = auto_in_ar_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_20_r_ready = auto_in_r_ready & _T_1965_20; // @[LazyModule.scala 173:49]
  assign auto_out_19_aw_valid = in_0_aw_valid & requestAWIO_0_19; // @[LazyModule.scala 173:49]
  assign auto_out_19_aw_bits_id = auto_in_aw_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_19_aw_bits_addr = auto_in_aw_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_19_aw_bits_size = auto_in_aw_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_19_w_valid = in_0_w_valid & requestWIO_0_19; // @[LazyModule.scala 173:49]
  assign auto_out_19_w_bits_data = auto_in_w_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_19_w_bits_strb = auto_in_w_bits_strb; // @[LazyModule.scala 173:49]
  assign auto_out_19_w_bits_last = auto_in_w_bits_last; // @[LazyModule.scala 173:49]
  assign auto_out_19_b_ready = auto_in_b_ready & _T_2427_19; // @[LazyModule.scala 173:49]
  assign auto_out_19_ar_valid = in_0_ar_valid & requestARIO_0_19; // @[LazyModule.scala 173:49]
  assign auto_out_19_ar_bits_id = auto_in_ar_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_19_ar_bits_addr = auto_in_ar_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_19_ar_bits_size = auto_in_ar_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_19_r_ready = auto_in_r_ready & _T_1965_19; // @[LazyModule.scala 173:49]
  assign auto_out_18_aw_valid = in_0_aw_valid & requestAWIO_0_18; // @[LazyModule.scala 173:49]
  assign auto_out_18_aw_bits_id = auto_in_aw_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_18_aw_bits_addr = auto_in_aw_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_18_aw_bits_size = auto_in_aw_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_18_w_valid = in_0_w_valid & requestWIO_0_18; // @[LazyModule.scala 173:49]
  assign auto_out_18_w_bits_data = auto_in_w_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_18_w_bits_strb = auto_in_w_bits_strb; // @[LazyModule.scala 173:49]
  assign auto_out_18_w_bits_last = auto_in_w_bits_last; // @[LazyModule.scala 173:49]
  assign auto_out_18_b_ready = auto_in_b_ready & _T_2427_18; // @[LazyModule.scala 173:49]
  assign auto_out_18_ar_valid = in_0_ar_valid & requestARIO_0_18; // @[LazyModule.scala 173:49]
  assign auto_out_18_ar_bits_id = auto_in_ar_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_18_ar_bits_addr = auto_in_ar_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_18_ar_bits_size = auto_in_ar_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_18_r_ready = auto_in_r_ready & _T_1965_18; // @[LazyModule.scala 173:49]
  assign auto_out_17_aw_valid = in_0_aw_valid & requestAWIO_0_17; // @[LazyModule.scala 173:49]
  assign auto_out_17_aw_bits_id = auto_in_aw_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_17_aw_bits_addr = auto_in_aw_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_17_aw_bits_size = auto_in_aw_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_17_w_valid = in_0_w_valid & requestWIO_0_17; // @[LazyModule.scala 173:49]
  assign auto_out_17_w_bits_data = auto_in_w_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_17_w_bits_strb = auto_in_w_bits_strb; // @[LazyModule.scala 173:49]
  assign auto_out_17_w_bits_last = auto_in_w_bits_last; // @[LazyModule.scala 173:49]
  assign auto_out_17_b_ready = auto_in_b_ready & _T_2427_17; // @[LazyModule.scala 173:49]
  assign auto_out_17_ar_valid = in_0_ar_valid & requestARIO_0_17; // @[LazyModule.scala 173:49]
  assign auto_out_17_ar_bits_id = auto_in_ar_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_17_ar_bits_addr = auto_in_ar_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_17_ar_bits_size = auto_in_ar_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_17_r_ready = auto_in_r_ready & _T_1965_17; // @[LazyModule.scala 173:49]
  assign auto_out_16_aw_valid = in_0_aw_valid & requestAWIO_0_16; // @[LazyModule.scala 173:49]
  assign auto_out_16_aw_bits_id = auto_in_aw_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_16_aw_bits_addr = auto_in_aw_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_16_aw_bits_size = auto_in_aw_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_16_w_valid = in_0_w_valid & requestWIO_0_16; // @[LazyModule.scala 173:49]
  assign auto_out_16_w_bits_data = auto_in_w_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_16_w_bits_strb = auto_in_w_bits_strb; // @[LazyModule.scala 173:49]
  assign auto_out_16_w_bits_last = auto_in_w_bits_last; // @[LazyModule.scala 173:49]
  assign auto_out_16_b_ready = auto_in_b_ready & _T_2427_16; // @[LazyModule.scala 173:49]
  assign auto_out_16_ar_valid = in_0_ar_valid & requestARIO_0_16; // @[LazyModule.scala 173:49]
  assign auto_out_16_ar_bits_id = auto_in_ar_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_16_ar_bits_addr = auto_in_ar_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_16_ar_bits_size = auto_in_ar_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_16_r_ready = auto_in_r_ready & _T_1965_16; // @[LazyModule.scala 173:49]
  assign auto_out_15_aw_valid = in_0_aw_valid & requestAWIO_0_15; // @[LazyModule.scala 173:49]
  assign auto_out_15_aw_bits_id = auto_in_aw_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_15_aw_bits_addr = auto_in_aw_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_15_aw_bits_size = auto_in_aw_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_15_w_valid = in_0_w_valid & requestWIO_0_15; // @[LazyModule.scala 173:49]
  assign auto_out_15_w_bits_data = auto_in_w_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_15_w_bits_strb = auto_in_w_bits_strb; // @[LazyModule.scala 173:49]
  assign auto_out_15_w_bits_last = auto_in_w_bits_last; // @[LazyModule.scala 173:49]
  assign auto_out_15_b_ready = auto_in_b_ready & _T_2427_15; // @[LazyModule.scala 173:49]
  assign auto_out_15_ar_valid = in_0_ar_valid & requestARIO_0_15; // @[LazyModule.scala 173:49]
  assign auto_out_15_ar_bits_id = auto_in_ar_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_15_ar_bits_addr = auto_in_ar_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_15_ar_bits_size = auto_in_ar_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_15_r_ready = auto_in_r_ready & _T_1965_15; // @[LazyModule.scala 173:49]
  assign auto_out_14_aw_valid = in_0_aw_valid & requestAWIO_0_14; // @[LazyModule.scala 173:49]
  assign auto_out_14_aw_bits_id = auto_in_aw_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_14_aw_bits_addr = auto_in_aw_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_14_aw_bits_size = auto_in_aw_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_14_w_valid = in_0_w_valid & requestWIO_0_14; // @[LazyModule.scala 173:49]
  assign auto_out_14_w_bits_data = auto_in_w_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_14_w_bits_strb = auto_in_w_bits_strb; // @[LazyModule.scala 173:49]
  assign auto_out_14_w_bits_last = auto_in_w_bits_last; // @[LazyModule.scala 173:49]
  assign auto_out_14_b_ready = auto_in_b_ready & _T_2427_14; // @[LazyModule.scala 173:49]
  assign auto_out_14_ar_valid = in_0_ar_valid & requestARIO_0_14; // @[LazyModule.scala 173:49]
  assign auto_out_14_ar_bits_id = auto_in_ar_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_14_ar_bits_addr = auto_in_ar_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_14_ar_bits_size = auto_in_ar_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_14_r_ready = auto_in_r_ready & _T_1965_14; // @[LazyModule.scala 173:49]
  assign auto_out_13_aw_valid = in_0_aw_valid & requestAWIO_0_13; // @[LazyModule.scala 173:49]
  assign auto_out_13_aw_bits_id = auto_in_aw_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_13_aw_bits_addr = auto_in_aw_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_13_aw_bits_size = auto_in_aw_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_13_w_valid = in_0_w_valid & requestWIO_0_13; // @[LazyModule.scala 173:49]
  assign auto_out_13_w_bits_data = auto_in_w_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_13_w_bits_strb = auto_in_w_bits_strb; // @[LazyModule.scala 173:49]
  assign auto_out_13_w_bits_last = auto_in_w_bits_last; // @[LazyModule.scala 173:49]
  assign auto_out_13_b_ready = auto_in_b_ready & _T_2427_13; // @[LazyModule.scala 173:49]
  assign auto_out_13_ar_valid = in_0_ar_valid & requestARIO_0_13; // @[LazyModule.scala 173:49]
  assign auto_out_13_ar_bits_id = auto_in_ar_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_13_ar_bits_addr = auto_in_ar_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_13_ar_bits_size = auto_in_ar_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_13_r_ready = auto_in_r_ready & _T_1965_13; // @[LazyModule.scala 173:49]
  assign auto_out_12_aw_valid = in_0_aw_valid & requestAWIO_0_12; // @[LazyModule.scala 173:49]
  assign auto_out_12_aw_bits_id = auto_in_aw_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_12_aw_bits_addr = auto_in_aw_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_12_aw_bits_size = auto_in_aw_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_12_w_valid = in_0_w_valid & requestWIO_0_12; // @[LazyModule.scala 173:49]
  assign auto_out_12_w_bits_data = auto_in_w_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_12_w_bits_strb = auto_in_w_bits_strb; // @[LazyModule.scala 173:49]
  assign auto_out_12_w_bits_last = auto_in_w_bits_last; // @[LazyModule.scala 173:49]
  assign auto_out_12_b_ready = auto_in_b_ready & _T_2427_12; // @[LazyModule.scala 173:49]
  assign auto_out_12_ar_valid = in_0_ar_valid & requestARIO_0_12; // @[LazyModule.scala 173:49]
  assign auto_out_12_ar_bits_id = auto_in_ar_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_12_ar_bits_addr = auto_in_ar_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_12_ar_bits_size = auto_in_ar_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_12_r_ready = auto_in_r_ready & _T_1965_12; // @[LazyModule.scala 173:49]
  assign auto_out_11_aw_valid = in_0_aw_valid & requestAWIO_0_11; // @[LazyModule.scala 173:49]
  assign auto_out_11_aw_bits_id = auto_in_aw_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_11_aw_bits_addr = auto_in_aw_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_11_aw_bits_size = auto_in_aw_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_11_w_valid = in_0_w_valid & requestWIO_0_11; // @[LazyModule.scala 173:49]
  assign auto_out_11_w_bits_data = auto_in_w_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_11_w_bits_strb = auto_in_w_bits_strb; // @[LazyModule.scala 173:49]
  assign auto_out_11_w_bits_last = auto_in_w_bits_last; // @[LazyModule.scala 173:49]
  assign auto_out_11_b_ready = auto_in_b_ready & _T_2427_11; // @[LazyModule.scala 173:49]
  assign auto_out_11_ar_valid = in_0_ar_valid & requestARIO_0_11; // @[LazyModule.scala 173:49]
  assign auto_out_11_ar_bits_id = auto_in_ar_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_11_ar_bits_addr = auto_in_ar_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_11_ar_bits_size = auto_in_ar_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_11_r_ready = auto_in_r_ready & _T_1965_11; // @[LazyModule.scala 173:49]
  assign auto_out_10_aw_valid = in_0_aw_valid & requestAWIO_0_10; // @[LazyModule.scala 173:49]
  assign auto_out_10_aw_bits_id = auto_in_aw_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_10_aw_bits_addr = auto_in_aw_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_10_aw_bits_size = auto_in_aw_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_10_w_valid = in_0_w_valid & requestWIO_0_10; // @[LazyModule.scala 173:49]
  assign auto_out_10_w_bits_data = auto_in_w_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_10_w_bits_strb = auto_in_w_bits_strb; // @[LazyModule.scala 173:49]
  assign auto_out_10_w_bits_last = auto_in_w_bits_last; // @[LazyModule.scala 173:49]
  assign auto_out_10_b_ready = auto_in_b_ready & _T_2427_10; // @[LazyModule.scala 173:49]
  assign auto_out_10_ar_valid = in_0_ar_valid & requestARIO_0_10; // @[LazyModule.scala 173:49]
  assign auto_out_10_ar_bits_id = auto_in_ar_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_10_ar_bits_addr = auto_in_ar_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_10_ar_bits_size = auto_in_ar_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_10_r_ready = auto_in_r_ready & _T_1965_10; // @[LazyModule.scala 173:49]
  assign auto_out_9_aw_valid = in_0_aw_valid & requestAWIO_0_9; // @[LazyModule.scala 173:49]
  assign auto_out_9_aw_bits_id = auto_in_aw_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_9_aw_bits_addr = auto_in_aw_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_9_aw_bits_size = auto_in_aw_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_9_w_valid = in_0_w_valid & requestWIO_0_9; // @[LazyModule.scala 173:49]
  assign auto_out_9_w_bits_data = auto_in_w_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_9_w_bits_strb = auto_in_w_bits_strb; // @[LazyModule.scala 173:49]
  assign auto_out_9_w_bits_last = auto_in_w_bits_last; // @[LazyModule.scala 173:49]
  assign auto_out_9_b_ready = auto_in_b_ready & _T_2427_9; // @[LazyModule.scala 173:49]
  assign auto_out_9_ar_valid = in_0_ar_valid & requestARIO_0_9; // @[LazyModule.scala 173:49]
  assign auto_out_9_ar_bits_id = auto_in_ar_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_9_ar_bits_addr = auto_in_ar_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_9_ar_bits_size = auto_in_ar_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_9_r_ready = auto_in_r_ready & _T_1965_9; // @[LazyModule.scala 173:49]
  assign auto_out_8_aw_valid = in_0_aw_valid & requestAWIO_0_8; // @[LazyModule.scala 173:49]
  assign auto_out_8_aw_bits_id = auto_in_aw_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_8_aw_bits_addr = auto_in_aw_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_8_aw_bits_size = auto_in_aw_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_8_w_valid = in_0_w_valid & requestWIO_0_8; // @[LazyModule.scala 173:49]
  assign auto_out_8_w_bits_data = auto_in_w_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_8_w_bits_strb = auto_in_w_bits_strb; // @[LazyModule.scala 173:49]
  assign auto_out_8_w_bits_last = auto_in_w_bits_last; // @[LazyModule.scala 173:49]
  assign auto_out_8_b_ready = auto_in_b_ready & _T_2427_8; // @[LazyModule.scala 173:49]
  assign auto_out_8_ar_valid = in_0_ar_valid & requestARIO_0_8; // @[LazyModule.scala 173:49]
  assign auto_out_8_ar_bits_id = auto_in_ar_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_8_ar_bits_addr = auto_in_ar_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_8_ar_bits_size = auto_in_ar_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_8_r_ready = auto_in_r_ready & _T_1965_8; // @[LazyModule.scala 173:49]
  assign auto_out_7_aw_valid = in_0_aw_valid & requestAWIO_0_7; // @[LazyModule.scala 173:49]
  assign auto_out_7_aw_bits_id = auto_in_aw_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_7_aw_bits_addr = auto_in_aw_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_7_aw_bits_size = auto_in_aw_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_7_w_valid = in_0_w_valid & requestWIO_0_7; // @[LazyModule.scala 173:49]
  assign auto_out_7_w_bits_data = auto_in_w_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_7_w_bits_strb = auto_in_w_bits_strb; // @[LazyModule.scala 173:49]
  assign auto_out_7_w_bits_last = auto_in_w_bits_last; // @[LazyModule.scala 173:49]
  assign auto_out_7_b_ready = auto_in_b_ready & _T_2427_7; // @[LazyModule.scala 173:49]
  assign auto_out_7_ar_valid = in_0_ar_valid & requestARIO_0_7; // @[LazyModule.scala 173:49]
  assign auto_out_7_ar_bits_id = auto_in_ar_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_7_ar_bits_addr = auto_in_ar_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_7_ar_bits_size = auto_in_ar_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_7_r_ready = auto_in_r_ready & _T_1965_7; // @[LazyModule.scala 173:49]
  assign auto_out_6_aw_valid = in_0_aw_valid & requestAWIO_0_6; // @[LazyModule.scala 173:49]
  assign auto_out_6_aw_bits_id = auto_in_aw_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_6_aw_bits_addr = auto_in_aw_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_6_aw_bits_size = auto_in_aw_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_6_w_valid = in_0_w_valid & requestWIO_0_6; // @[LazyModule.scala 173:49]
  assign auto_out_6_w_bits_data = auto_in_w_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_6_w_bits_strb = auto_in_w_bits_strb; // @[LazyModule.scala 173:49]
  assign auto_out_6_w_bits_last = auto_in_w_bits_last; // @[LazyModule.scala 173:49]
  assign auto_out_6_b_ready = auto_in_b_ready & _T_2427_6; // @[LazyModule.scala 173:49]
  assign auto_out_6_ar_valid = in_0_ar_valid & requestARIO_0_6; // @[LazyModule.scala 173:49]
  assign auto_out_6_ar_bits_id = auto_in_ar_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_6_ar_bits_addr = auto_in_ar_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_6_ar_bits_size = auto_in_ar_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_6_r_ready = auto_in_r_ready & _T_1965_6; // @[LazyModule.scala 173:49]
  assign auto_out_5_aw_valid = in_0_aw_valid & requestAWIO_0_5; // @[LazyModule.scala 173:49]
  assign auto_out_5_aw_bits_id = auto_in_aw_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_5_aw_bits_addr = auto_in_aw_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_5_aw_bits_size = auto_in_aw_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_5_w_valid = in_0_w_valid & requestWIO_0_5; // @[LazyModule.scala 173:49]
  assign auto_out_5_w_bits_data = auto_in_w_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_5_w_bits_strb = auto_in_w_bits_strb; // @[LazyModule.scala 173:49]
  assign auto_out_5_w_bits_last = auto_in_w_bits_last; // @[LazyModule.scala 173:49]
  assign auto_out_5_b_ready = auto_in_b_ready & _T_2427_5; // @[LazyModule.scala 173:49]
  assign auto_out_5_ar_valid = in_0_ar_valid & requestARIO_0_5; // @[LazyModule.scala 173:49]
  assign auto_out_5_ar_bits_id = auto_in_ar_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_5_ar_bits_addr = auto_in_ar_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_5_ar_bits_size = auto_in_ar_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_5_r_ready = auto_in_r_ready & _T_1965_5; // @[LazyModule.scala 173:49]
  assign auto_out_4_aw_valid = in_0_aw_valid & requestAWIO_0_4; // @[LazyModule.scala 173:49]
  assign auto_out_4_aw_bits_id = auto_in_aw_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_4_aw_bits_addr = auto_in_aw_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_4_aw_bits_size = auto_in_aw_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_4_w_valid = in_0_w_valid & requestWIO_0_4; // @[LazyModule.scala 173:49]
  assign auto_out_4_w_bits_data = auto_in_w_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_4_w_bits_strb = auto_in_w_bits_strb; // @[LazyModule.scala 173:49]
  assign auto_out_4_w_bits_last = auto_in_w_bits_last; // @[LazyModule.scala 173:49]
  assign auto_out_4_b_ready = auto_in_b_ready & _T_2427_4; // @[LazyModule.scala 173:49]
  assign auto_out_4_ar_valid = in_0_ar_valid & requestARIO_0_4; // @[LazyModule.scala 173:49]
  assign auto_out_4_ar_bits_id = auto_in_ar_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_4_ar_bits_addr = auto_in_ar_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_4_ar_bits_size = auto_in_ar_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_4_r_ready = auto_in_r_ready & _T_1965_4; // @[LazyModule.scala 173:49]
  assign auto_out_3_aw_valid = in_0_aw_valid & requestAWIO_0_3; // @[LazyModule.scala 173:49]
  assign auto_out_3_aw_bits_id = auto_in_aw_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_3_aw_bits_addr = auto_in_aw_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_3_aw_bits_size = auto_in_aw_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_3_w_valid = in_0_w_valid & requestWIO_0_3; // @[LazyModule.scala 173:49]
  assign auto_out_3_w_bits_data = auto_in_w_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_3_w_bits_strb = auto_in_w_bits_strb; // @[LazyModule.scala 173:49]
  assign auto_out_3_w_bits_last = auto_in_w_bits_last; // @[LazyModule.scala 173:49]
  assign auto_out_3_b_ready = auto_in_b_ready & _T_2427_3; // @[LazyModule.scala 173:49]
  assign auto_out_3_ar_valid = in_0_ar_valid & requestARIO_0_3; // @[LazyModule.scala 173:49]
  assign auto_out_3_ar_bits_id = auto_in_ar_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_3_ar_bits_addr = auto_in_ar_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_3_ar_bits_size = auto_in_ar_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_3_r_ready = auto_in_r_ready & _T_1965_3; // @[LazyModule.scala 173:49]
  assign auto_out_2_aw_valid = in_0_aw_valid & requestAWIO_0_2; // @[LazyModule.scala 173:49]
  assign auto_out_2_aw_bits_id = auto_in_aw_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_2_aw_bits_addr = auto_in_aw_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_2_aw_bits_size = auto_in_aw_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_2_w_valid = in_0_w_valid & requestWIO_0_2; // @[LazyModule.scala 173:49]
  assign auto_out_2_w_bits_data = auto_in_w_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_2_w_bits_strb = auto_in_w_bits_strb; // @[LazyModule.scala 173:49]
  assign auto_out_2_w_bits_last = auto_in_w_bits_last; // @[LazyModule.scala 173:49]
  assign auto_out_2_b_ready = auto_in_b_ready & _T_2427_2; // @[LazyModule.scala 173:49]
  assign auto_out_2_ar_valid = in_0_ar_valid & requestARIO_0_2; // @[LazyModule.scala 173:49]
  assign auto_out_2_ar_bits_id = auto_in_ar_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_2_ar_bits_addr = auto_in_ar_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_2_ar_bits_size = auto_in_ar_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_2_r_ready = auto_in_r_ready & _T_1965_2; // @[LazyModule.scala 173:49]
  assign auto_out_1_aw_valid = in_0_aw_valid & requestAWIO_0_1; // @[LazyModule.scala 173:49]
  assign auto_out_1_aw_bits_id = auto_in_aw_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_1_aw_bits_addr = auto_in_aw_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_1_aw_bits_size = auto_in_aw_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_1_w_valid = in_0_w_valid & requestWIO_0_1; // @[LazyModule.scala 173:49]
  assign auto_out_1_w_bits_data = auto_in_w_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_1_w_bits_strb = auto_in_w_bits_strb; // @[LazyModule.scala 173:49]
  assign auto_out_1_w_bits_last = auto_in_w_bits_last; // @[LazyModule.scala 173:49]
  assign auto_out_1_b_ready = auto_in_b_ready & _T_2427_1; // @[LazyModule.scala 173:49]
  assign auto_out_1_ar_valid = in_0_ar_valid & requestARIO_0_1; // @[LazyModule.scala 173:49]
  assign auto_out_1_ar_bits_id = auto_in_ar_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_1_ar_bits_addr = auto_in_ar_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_1_ar_bits_size = auto_in_ar_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_1_r_ready = auto_in_r_ready & _T_1965_1; // @[LazyModule.scala 173:49]
  assign auto_out_0_aw_valid = in_0_aw_valid & requestAWIO_0_0; // @[LazyModule.scala 173:49]
  assign auto_out_0_aw_bits_id = auto_in_aw_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_0_aw_bits_addr = auto_in_aw_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_0_aw_bits_size = auto_in_aw_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_0_w_valid = in_0_w_valid & requestWIO_0_0; // @[LazyModule.scala 173:49]
  assign auto_out_0_w_bits_data = auto_in_w_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_0_w_bits_strb = auto_in_w_bits_strb; // @[LazyModule.scala 173:49]
  assign auto_out_0_w_bits_last = auto_in_w_bits_last; // @[LazyModule.scala 173:49]
  assign auto_out_0_b_ready = auto_in_b_ready & _T_2427_0; // @[LazyModule.scala 173:49]
  assign auto_out_0_ar_valid = in_0_ar_valid & requestARIO_0_0; // @[LazyModule.scala 173:49]
  assign auto_out_0_ar_bits_id = auto_in_ar_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_0_ar_bits_addr = auto_in_ar_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_0_ar_bits_size = auto_in_ar_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_0_r_ready = auto_in_r_ready & _T_1965_0; // @[LazyModule.scala 173:49]
  assign awIn_0_clock = clock;
  assign awIn_0_reset = reset;
  assign awIn_0_io_enq_valid = auto_in_aw_valid & _T_421; // @[Xbar.scala 140:30]
  assign awIn_0_io_enq_bits = {_T_263,_T_253}; // @[Xbar.scala 64:57]
  assign awIn_0_io_deq_ready = _T_427 & in_0_w_ready; // @[Xbar.scala 147:30]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_360 = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_361 = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_1686 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_1962_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_1962_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_1962_2 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_1962_3 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_1962_4 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_1962_5 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_1962_6 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_1962_7 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_1962_8 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_1962_9 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_1962_10 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_1962_11 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_1962_12 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_1962_13 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_1962_14 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_1962_15 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_1962_16 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_1962_17 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_1962_18 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_1962_19 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_1962_20 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_1962_21 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_1735 = _RAND_25[21:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_414 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T_388 = _RAND_27[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_389 = _RAND_28[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_2148 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_2424_0 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T_2424_1 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _T_2424_2 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _T_2424_3 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _T_2424_4 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _T_2424_5 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _T_2424_6 = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _T_2424_7 = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _T_2424_8 = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _T_2424_9 = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _T_2424_10 = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  _T_2424_11 = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  _T_2424_12 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  _T_2424_13 = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  _T_2424_14 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  _T_2424_15 = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  _T_2424_16 = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  _T_2424_17 = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  _T_2424_18 = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  _T_2424_19 = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  _T_2424_20 = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  _T_2424_21 = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  _T_2197 = _RAND_52[21:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      _T_360 <= 3'h0;
    end else begin
      _T_360 <= _T_365;
    end
    if (_T_355) begin
      _T_361 <= _T_312;
    end
    _T_1686 <= reset | _GEN_94;
    if (reset) begin
      _T_1962_0 <= 1'h0;
    end else if (_T_1686) begin
      _T_1962_0 <= _T_1800;
    end
    if (reset) begin
      _T_1962_1 <= 1'h0;
    end else if (_T_1686) begin
      _T_1962_1 <= _T_1801;
    end
    if (reset) begin
      _T_1962_2 <= 1'h0;
    end else if (_T_1686) begin
      _T_1962_2 <= _T_1802;
    end
    if (reset) begin
      _T_1962_3 <= 1'h0;
    end else if (_T_1686) begin
      _T_1962_3 <= _T_1803;
    end
    if (reset) begin
      _T_1962_4 <= 1'h0;
    end else if (_T_1686) begin
      _T_1962_4 <= _T_1804;
    end
    if (reset) begin
      _T_1962_5 <= 1'h0;
    end else if (_T_1686) begin
      _T_1962_5 <= _T_1805;
    end
    if (reset) begin
      _T_1962_6 <= 1'h0;
    end else if (_T_1686) begin
      _T_1962_6 <= _T_1806;
    end
    if (reset) begin
      _T_1962_7 <= 1'h0;
    end else if (_T_1686) begin
      _T_1962_7 <= _T_1807;
    end
    if (reset) begin
      _T_1962_8 <= 1'h0;
    end else if (_T_1686) begin
      _T_1962_8 <= _T_1808;
    end
    if (reset) begin
      _T_1962_9 <= 1'h0;
    end else if (_T_1686) begin
      _T_1962_9 <= _T_1809;
    end
    if (reset) begin
      _T_1962_10 <= 1'h0;
    end else if (_T_1686) begin
      _T_1962_10 <= _T_1810;
    end
    if (reset) begin
      _T_1962_11 <= 1'h0;
    end else if (_T_1686) begin
      _T_1962_11 <= _T_1811;
    end
    if (reset) begin
      _T_1962_12 <= 1'h0;
    end else if (_T_1686) begin
      _T_1962_12 <= _T_1812;
    end
    if (reset) begin
      _T_1962_13 <= 1'h0;
    end else if (_T_1686) begin
      _T_1962_13 <= _T_1813;
    end
    if (reset) begin
      _T_1962_14 <= 1'h0;
    end else if (_T_1686) begin
      _T_1962_14 <= _T_1814;
    end
    if (reset) begin
      _T_1962_15 <= 1'h0;
    end else if (_T_1686) begin
      _T_1962_15 <= _T_1815;
    end
    if (reset) begin
      _T_1962_16 <= 1'h0;
    end else if (_T_1686) begin
      _T_1962_16 <= _T_1816;
    end
    if (reset) begin
      _T_1962_17 <= 1'h0;
    end else if (_T_1686) begin
      _T_1962_17 <= _T_1817;
    end
    if (reset) begin
      _T_1962_18 <= 1'h0;
    end else if (_T_1686) begin
      _T_1962_18 <= _T_1818;
    end
    if (reset) begin
      _T_1962_19 <= 1'h0;
    end else if (_T_1686) begin
      _T_1962_19 <= _T_1819;
    end
    if (reset) begin
      _T_1962_20 <= 1'h0;
    end else if (_T_1686) begin
      _T_1962_20 <= _T_1820;
    end
    if (reset) begin
      _T_1962_21 <= 1'h0;
    end else if (_T_1686) begin
      _T_1962_21 <= _T_1821;
    end
    if (reset) begin
      _T_1735 <= 22'h3fffff;
    end else if (_T_1758) begin
      _T_1735 <= _T_1774;
    end
    if (reset) begin
      _T_414 <= 1'h0;
    end else if (_T_424) begin
      _T_414 <= 1'h0;
    end else begin
      _T_414 <= _GEN_2;
    end
    if (reset) begin
      _T_388 <= 3'h0;
    end else begin
      _T_388 <= _T_393;
    end
    if (_T_384) begin
      _T_389 <= _T_354;
    end
    _T_2148 <= reset | _GEN_97;
    if (reset) begin
      _T_2424_0 <= 1'h0;
    end else if (_T_2148) begin
      _T_2424_0 <= _T_2262;
    end
    if (reset) begin
      _T_2424_1 <= 1'h0;
    end else if (_T_2148) begin
      _T_2424_1 <= _T_2263;
    end
    if (reset) begin
      _T_2424_2 <= 1'h0;
    end else if (_T_2148) begin
      _T_2424_2 <= _T_2264;
    end
    if (reset) begin
      _T_2424_3 <= 1'h0;
    end else if (_T_2148) begin
      _T_2424_3 <= _T_2265;
    end
    if (reset) begin
      _T_2424_4 <= 1'h0;
    end else if (_T_2148) begin
      _T_2424_4 <= _T_2266;
    end
    if (reset) begin
      _T_2424_5 <= 1'h0;
    end else if (_T_2148) begin
      _T_2424_5 <= _T_2267;
    end
    if (reset) begin
      _T_2424_6 <= 1'h0;
    end else if (_T_2148) begin
      _T_2424_6 <= _T_2268;
    end
    if (reset) begin
      _T_2424_7 <= 1'h0;
    end else if (_T_2148) begin
      _T_2424_7 <= _T_2269;
    end
    if (reset) begin
      _T_2424_8 <= 1'h0;
    end else if (_T_2148) begin
      _T_2424_8 <= _T_2270;
    end
    if (reset) begin
      _T_2424_9 <= 1'h0;
    end else if (_T_2148) begin
      _T_2424_9 <= _T_2271;
    end
    if (reset) begin
      _T_2424_10 <= 1'h0;
    end else if (_T_2148) begin
      _T_2424_10 <= _T_2272;
    end
    if (reset) begin
      _T_2424_11 <= 1'h0;
    end else if (_T_2148) begin
      _T_2424_11 <= _T_2273;
    end
    if (reset) begin
      _T_2424_12 <= 1'h0;
    end else if (_T_2148) begin
      _T_2424_12 <= _T_2274;
    end
    if (reset) begin
      _T_2424_13 <= 1'h0;
    end else if (_T_2148) begin
      _T_2424_13 <= _T_2275;
    end
    if (reset) begin
      _T_2424_14 <= 1'h0;
    end else if (_T_2148) begin
      _T_2424_14 <= _T_2276;
    end
    if (reset) begin
      _T_2424_15 <= 1'h0;
    end else if (_T_2148) begin
      _T_2424_15 <= _T_2277;
    end
    if (reset) begin
      _T_2424_16 <= 1'h0;
    end else if (_T_2148) begin
      _T_2424_16 <= _T_2278;
    end
    if (reset) begin
      _T_2424_17 <= 1'h0;
    end else if (_T_2148) begin
      _T_2424_17 <= _T_2279;
    end
    if (reset) begin
      _T_2424_18 <= 1'h0;
    end else if (_T_2148) begin
      _T_2424_18 <= _T_2280;
    end
    if (reset) begin
      _T_2424_19 <= 1'h0;
    end else if (_T_2148) begin
      _T_2424_19 <= _T_2281;
    end
    if (reset) begin
      _T_2424_20 <= 1'h0;
    end else if (_T_2148) begin
      _T_2424_20 <= _T_2282;
    end
    if (reset) begin
      _T_2424_21 <= 1'h0;
    end else if (_T_2148) begin
      _T_2424_21 <= _T_2283;
    end
    if (reset) begin
      _T_2197 <= 22'h3fffff;
    end else if (_T_2220) begin
      _T_2197 <= _T_2236;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_371) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:107 assert (!resp_fire || count =/= UInt(0))\n"); // @[Xbar.scala 107:22]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_371) begin
          $fatal; // @[Xbar.scala 107:22]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_377) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:108 assert (!req_fire  || count =/= UInt(flight))\n"); // @[Xbar.scala 108:22]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_377) begin
          $fatal; // @[Xbar.scala 108:22]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_399) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:107 assert (!resp_fire || count =/= UInt(0))\n"); // @[Xbar.scala 107:22]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_399) begin
          $fatal; // @[Xbar.scala 107:22]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_405) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:108 assert (!req_fire  || count =/= UInt(flight))\n"); // @[Xbar.scala 108:22]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_405) begin
          $fatal; // @[Xbar.scala 108:22]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_733) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_733) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_754) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_754) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_777) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_777) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_798) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_798) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_821) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_821) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_842) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_842) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_865) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_865) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_886) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_886) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_909) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_909) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_930) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_930) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_953) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_953) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_974) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_974) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_997) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_997) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1018) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1018) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1041) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1041) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1062) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1062) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1085) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1085) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1106) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1106) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1129) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1129) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1150) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1150) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1173) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1173) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1194) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1194) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1217) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1217) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1238) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1238) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1261) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1261) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1282) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1282) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1305) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1305) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1326) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1326) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1349) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1349) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1370) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1370) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1393) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1393) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1414) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1414) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1437) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1437) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1458) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1458) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1481) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1481) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1502) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1502) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1525) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1525) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1546) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1546) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1569) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1569) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1590) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1590) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1613) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1613) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1634) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1634) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1657) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1657) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1678) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1678) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1934) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:256 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n"); // @[Xbar.scala 256:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1934) begin
          $fatal; // @[Xbar.scala 256:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1960) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1960) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2396) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:256 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n"); // @[Xbar.scala 256:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2396) begin
          $fatal; // @[Xbar.scala 256:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2422) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2422) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module Queue_147(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [31:0] io_enq_bits_data,
  input         io_enq_bits_last,
  input         io_deq_ready,
  output        io_deq_valid,
  output [31:0] io_deq_bits_data,
  output        io_deq_bits_last
);
  reg [31:0] _T_data [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_0;
  wire [31:0] _T_data__T_18_data; // @[Decoupled.scala 209:24]
  wire  _T_data__T_18_addr; // @[Decoupled.scala 209:24]
  wire [31:0] _T_data__T_10_data; // @[Decoupled.scala 209:24]
  wire  _T_data__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T_data__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T_data__T_10_en; // @[Decoupled.scala 209:24]
  reg  _T_last [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_1;
  wire  _T_last__T_18_data; // @[Decoupled.scala 209:24]
  wire  _T_last__T_18_addr; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_data; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_en; // @[Decoupled.scala 209:24]
  reg  value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_2;
  reg  value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_3;
  reg  _T_1; // @[Decoupled.scala 212:35]
  reg [31:0] _RAND_4;
  wire  _T_2; // @[Decoupled.scala 214:41]
  wire  _T_3; // @[Decoupled.scala 215:36]
  wire  _T_4; // @[Decoupled.scala 215:33]
  wire  _T_5; // @[Decoupled.scala 216:32]
  wire  _T_6; // @[Decoupled.scala 40:37]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _T_12; // @[Counter.scala 39:22]
  wire  _T_14; // @[Counter.scala 39:22]
  wire  _T_15; // @[Decoupled.scala 227:16]
  assign _T_data__T_18_addr = value_1;
  assign _T_data__T_18_data = _T_data[_T_data__T_18_addr]; // @[Decoupled.scala 209:24]
  assign _T_data__T_10_data = io_enq_bits_data;
  assign _T_data__T_10_addr = value;
  assign _T_data__T_10_mask = 1'h1;
  assign _T_data__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_last__T_18_addr = value_1;
  assign _T_last__T_18_data = _T_last[_T_last__T_18_addr]; // @[Decoupled.scala 209:24]
  assign _T_last__T_10_data = io_enq_bits_last;
  assign _T_last__T_10_addr = value;
  assign _T_last__T_10_mask = 1'h1;
  assign _T_last__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_2 = value == value_1; // @[Decoupled.scala 214:41]
  assign _T_3 = ~_T_1; // @[Decoupled.scala 215:36]
  assign _T_4 = _T_2 & _T_3; // @[Decoupled.scala 215:33]
  assign _T_5 = _T_2 & _T_1; // @[Decoupled.scala 216:32]
  assign _T_6 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  assign _T_8 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  assign _T_12 = value + 1'h1; // @[Counter.scala 39:22]
  assign _T_14 = value_1 + 1'h1; // @[Counter.scala 39:22]
  assign _T_15 = _T_6 != _T_8; // @[Decoupled.scala 227:16]
  assign io_enq_ready = ~_T_5; // @[Decoupled.scala 232:16]
  assign io_deq_valid = ~_T_4; // @[Decoupled.scala 231:16]
  assign io_deq_bits_data = _T_data__T_18_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_last = _T_last__T_18_data; // @[Decoupled.scala 233:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_data[initvar] = _RAND_0[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_last[initvar] = _RAND_1[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  value = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  value_1 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T_data__T_10_en & _T_data__T_10_mask) begin
      _T_data[_T_data__T_10_addr] <= _T_data__T_10_data; // @[Decoupled.scala 209:24]
    end
    if(_T_last__T_10_en & _T_last__T_10_mask) begin
      _T_last[_T_last__T_10_addr] <= _T_last__T_10_data; // @[Decoupled.scala 209:24]
    end
    if (reset) begin
      value <= 1'h0;
    end else if (_T_6) begin
      value <= _T_12;
    end
    if (reset) begin
      value_1 <= 1'h0;
    end else if (_T_8) begin
      value_1 <= _T_14;
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else if (_T_15) begin
      _T_1 <= _T_6;
    end
  end
endmodule
module AXI4StreamBuffer(
  input         clock,
  input         reset,
  output        auto_in_ready,
  input         auto_in_valid,
  input  [31:0] auto_in_bits_data,
  input         auto_in_bits_last,
  input         auto_out_ready,
  output        auto_out_valid,
  output [31:0] auto_out_bits_data,
  output        auto_out_bits_last
);
  wire  Queue_clock; // @[Decoupled.scala 287:21]
  wire  Queue_reset; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_enq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_last; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_deq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_last; // @[Decoupled.scala 287:21]
  Queue_147 Queue ( // @[Decoupled.scala 287:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_last(Queue_io_enq_bits_last),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_last(Queue_io_deq_bits_last)
  );
  assign auto_in_ready = Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_out_valid = Queue_io_deq_valid; // @[LazyModule.scala 173:49]
  assign auto_out_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_bits_last = Queue_io_deq_bits_last; // @[LazyModule.scala 173:49]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_in_valid; // @[Decoupled.scala 288:22]
  assign Queue_io_enq_bits_data = auto_in_bits_data; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_last = auto_in_bits_last; // @[Decoupled.scala 289:21]
  assign Queue_io_deq_ready = auto_out_ready; // @[Decoupled.scala 311:15]
endmodule
module Queue_148(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [31:0] io_enq_bits_data,
  input         io_enq_bits_last,
  input         io_deq_ready,
  output        io_deq_valid,
  output [31:0] io_deq_bits_data,
  output        io_deq_bits_last
);
  reg [31:0] _T_data [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_0;
  wire [31:0] _T_data__T_18_data; // @[Decoupled.scala 209:24]
  wire  _T_data__T_18_addr; // @[Decoupled.scala 209:24]
  wire [31:0] _T_data__T_10_data; // @[Decoupled.scala 209:24]
  wire  _T_data__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T_data__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T_data__T_10_en; // @[Decoupled.scala 209:24]
  reg  _T_last [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_1;
  wire  _T_last__T_18_data; // @[Decoupled.scala 209:24]
  wire  _T_last__T_18_addr; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_data; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_en; // @[Decoupled.scala 209:24]
  reg  value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_2;
  reg  value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_3;
  reg  _T_1; // @[Decoupled.scala 212:35]
  reg [31:0] _RAND_4;
  wire  _T_2; // @[Decoupled.scala 214:41]
  wire  _T_3; // @[Decoupled.scala 215:36]
  wire  _T_4; // @[Decoupled.scala 215:33]
  wire  _T_5; // @[Decoupled.scala 216:32]
  wire  _T_6; // @[Decoupled.scala 40:37]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _T_12; // @[Counter.scala 39:22]
  wire  _T_14; // @[Counter.scala 39:22]
  wire  _T_15; // @[Decoupled.scala 227:16]
  assign _T_data__T_18_addr = value_1;
  assign _T_data__T_18_data = _T_data[_T_data__T_18_addr]; // @[Decoupled.scala 209:24]
  assign _T_data__T_10_data = io_enq_bits_data;
  assign _T_data__T_10_addr = value;
  assign _T_data__T_10_mask = 1'h1;
  assign _T_data__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_last__T_18_addr = value_1;
  assign _T_last__T_18_data = _T_last[_T_last__T_18_addr]; // @[Decoupled.scala 209:24]
  assign _T_last__T_10_data = io_enq_bits_last;
  assign _T_last__T_10_addr = value;
  assign _T_last__T_10_mask = 1'h1;
  assign _T_last__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_2 = value == value_1; // @[Decoupled.scala 214:41]
  assign _T_3 = ~_T_1; // @[Decoupled.scala 215:36]
  assign _T_4 = _T_2 & _T_3; // @[Decoupled.scala 215:33]
  assign _T_5 = _T_2 & _T_1; // @[Decoupled.scala 216:32]
  assign _T_6 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  assign _T_8 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  assign _T_12 = value + 1'h1; // @[Counter.scala 39:22]
  assign _T_14 = value_1 + 1'h1; // @[Counter.scala 39:22]
  assign _T_15 = _T_6 != _T_8; // @[Decoupled.scala 227:16]
  assign io_enq_ready = ~_T_5; // @[Decoupled.scala 232:16]
  assign io_deq_valid = ~_T_4; // @[Decoupled.scala 231:16]
  assign io_deq_bits_data = _T_data__T_18_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_last = _T_last__T_18_data; // @[Decoupled.scala 233:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_data[initvar] = _RAND_0[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_last[initvar] = _RAND_1[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  value = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  value_1 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T_data__T_10_en & _T_data__T_10_mask) begin
      _T_data[_T_data__T_10_addr] <= _T_data__T_10_data; // @[Decoupled.scala 209:24]
    end
    if(_T_last__T_10_en & _T_last__T_10_mask) begin
      _T_last[_T_last__T_10_addr] <= _T_last__T_10_data; // @[Decoupled.scala 209:24]
    end
    if (reset) begin
      value <= 1'h0;
    end else if (_T_6) begin
      value <= _T_12;
    end
    if (reset) begin
      value_1 <= 1'h0;
    end else if (_T_8) begin
      value_1 <= _T_14;
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else if (_T_15) begin
      _T_1 <= _T_6;
    end
  end
endmodule
module AXI4StreamBuffer_1(
  input         clock,
  input         reset,
  output        auto_in_ready,
  input         auto_in_valid,
  input  [31:0] auto_in_bits_data,
  input         auto_in_bits_last,
  input         auto_out_ready,
  output        auto_out_valid,
  output [31:0] auto_out_bits_data,
  output        auto_out_bits_last
);
  wire  Queue_clock; // @[Decoupled.scala 287:21]
  wire  Queue_reset; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_enq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_last; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_deq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_last; // @[Decoupled.scala 287:21]
  Queue_148 Queue ( // @[Decoupled.scala 287:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_last(Queue_io_enq_bits_last),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_last(Queue_io_deq_bits_last)
  );
  assign auto_in_ready = Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_out_valid = Queue_io_deq_valid; // @[LazyModule.scala 173:49]
  assign auto_out_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_bits_last = Queue_io_deq_bits_last; // @[LazyModule.scala 173:49]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_in_valid; // @[Decoupled.scala 288:22]
  assign Queue_io_enq_bits_data = auto_in_bits_data; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_last = auto_in_bits_last; // @[Decoupled.scala 289:21]
  assign Queue_io_deq_ready = auto_out_ready; // @[Decoupled.scala 311:15]
endmodule
module Queue_149(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [31:0] io_enq_bits_data,
  input         io_enq_bits_last,
  input         io_deq_ready,
  output        io_deq_valid,
  output [31:0] io_deq_bits_data,
  output        io_deq_bits_last
);
  reg [31:0] _T_data [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_0;
  wire [31:0] _T_data__T_18_data; // @[Decoupled.scala 209:24]
  wire  _T_data__T_18_addr; // @[Decoupled.scala 209:24]
  wire [31:0] _T_data__T_10_data; // @[Decoupled.scala 209:24]
  wire  _T_data__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T_data__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T_data__T_10_en; // @[Decoupled.scala 209:24]
  reg  _T_last [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_1;
  wire  _T_last__T_18_data; // @[Decoupled.scala 209:24]
  wire  _T_last__T_18_addr; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_data; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_en; // @[Decoupled.scala 209:24]
  reg  value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_2;
  reg  value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_3;
  reg  _T_1; // @[Decoupled.scala 212:35]
  reg [31:0] _RAND_4;
  wire  _T_2; // @[Decoupled.scala 214:41]
  wire  _T_3; // @[Decoupled.scala 215:36]
  wire  _T_4; // @[Decoupled.scala 215:33]
  wire  _T_5; // @[Decoupled.scala 216:32]
  wire  _T_6; // @[Decoupled.scala 40:37]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _T_12; // @[Counter.scala 39:22]
  wire  _T_14; // @[Counter.scala 39:22]
  wire  _T_15; // @[Decoupled.scala 227:16]
  assign _T_data__T_18_addr = value_1;
  assign _T_data__T_18_data = _T_data[_T_data__T_18_addr]; // @[Decoupled.scala 209:24]
  assign _T_data__T_10_data = io_enq_bits_data;
  assign _T_data__T_10_addr = value;
  assign _T_data__T_10_mask = 1'h1;
  assign _T_data__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_last__T_18_addr = value_1;
  assign _T_last__T_18_data = _T_last[_T_last__T_18_addr]; // @[Decoupled.scala 209:24]
  assign _T_last__T_10_data = io_enq_bits_last;
  assign _T_last__T_10_addr = value;
  assign _T_last__T_10_mask = 1'h1;
  assign _T_last__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_2 = value == value_1; // @[Decoupled.scala 214:41]
  assign _T_3 = ~_T_1; // @[Decoupled.scala 215:36]
  assign _T_4 = _T_2 & _T_3; // @[Decoupled.scala 215:33]
  assign _T_5 = _T_2 & _T_1; // @[Decoupled.scala 216:32]
  assign _T_6 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  assign _T_8 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  assign _T_12 = value + 1'h1; // @[Counter.scala 39:22]
  assign _T_14 = value_1 + 1'h1; // @[Counter.scala 39:22]
  assign _T_15 = _T_6 != _T_8; // @[Decoupled.scala 227:16]
  assign io_enq_ready = ~_T_5; // @[Decoupled.scala 232:16]
  assign io_deq_valid = ~_T_4; // @[Decoupled.scala 231:16]
  assign io_deq_bits_data = _T_data__T_18_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_last = _T_last__T_18_data; // @[Decoupled.scala 233:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_data[initvar] = _RAND_0[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_last[initvar] = _RAND_1[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  value = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  value_1 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T_data__T_10_en & _T_data__T_10_mask) begin
      _T_data[_T_data__T_10_addr] <= _T_data__T_10_data; // @[Decoupled.scala 209:24]
    end
    if(_T_last__T_10_en & _T_last__T_10_mask) begin
      _T_last[_T_last__T_10_addr] <= _T_last__T_10_data; // @[Decoupled.scala 209:24]
    end
    if (reset) begin
      value <= 1'h0;
    end else if (_T_6) begin
      value <= _T_12;
    end
    if (reset) begin
      value_1 <= 1'h0;
    end else if (_T_8) begin
      value_1 <= _T_14;
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else if (_T_15) begin
      _T_1 <= _T_6;
    end
  end
endmodule
module AXI4StreamBuffer_2(
  input         clock,
  input         reset,
  output        auto_in_ready,
  input         auto_in_valid,
  input  [31:0] auto_in_bits_data,
  input         auto_in_bits_last,
  input         auto_out_ready,
  output        auto_out_valid,
  output [31:0] auto_out_bits_data,
  output        auto_out_bits_last
);
  wire  Queue_clock; // @[Decoupled.scala 287:21]
  wire  Queue_reset; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_enq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_last; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_deq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_last; // @[Decoupled.scala 287:21]
  Queue_149 Queue ( // @[Decoupled.scala 287:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_last(Queue_io_enq_bits_last),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_last(Queue_io_deq_bits_last)
  );
  assign auto_in_ready = Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_out_valid = Queue_io_deq_valid; // @[LazyModule.scala 173:49]
  assign auto_out_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_bits_last = Queue_io_deq_bits_last; // @[LazyModule.scala 173:49]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_in_valid; // @[Decoupled.scala 288:22]
  assign Queue_io_enq_bits_data = auto_in_bits_data; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_last = auto_in_bits_last; // @[Decoupled.scala 289:21]
  assign Queue_io_deq_ready = auto_out_ready; // @[Decoupled.scala 311:15]
endmodule
module Queue_151(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [31:0] io_enq_bits_data,
  input         io_enq_bits_last,
  input         io_deq_ready,
  output        io_deq_valid,
  output [31:0] io_deq_bits_data,
  output        io_deq_bits_last
);
  reg [31:0] _T_data [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_0;
  wire [31:0] _T_data__T_18_data; // @[Decoupled.scala 209:24]
  wire  _T_data__T_18_addr; // @[Decoupled.scala 209:24]
  wire [31:0] _T_data__T_10_data; // @[Decoupled.scala 209:24]
  wire  _T_data__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T_data__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T_data__T_10_en; // @[Decoupled.scala 209:24]
  reg  _T_last [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_1;
  wire  _T_last__T_18_data; // @[Decoupled.scala 209:24]
  wire  _T_last__T_18_addr; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_data; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_en; // @[Decoupled.scala 209:24]
  reg  value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_2;
  reg  value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_3;
  reg  _T_1; // @[Decoupled.scala 212:35]
  reg [31:0] _RAND_4;
  wire  _T_2; // @[Decoupled.scala 214:41]
  wire  _T_3; // @[Decoupled.scala 215:36]
  wire  _T_4; // @[Decoupled.scala 215:33]
  wire  _T_5; // @[Decoupled.scala 216:32]
  wire  _T_6; // @[Decoupled.scala 40:37]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _T_12; // @[Counter.scala 39:22]
  wire  _T_14; // @[Counter.scala 39:22]
  wire  _T_15; // @[Decoupled.scala 227:16]
  assign _T_data__T_18_addr = value_1;
  assign _T_data__T_18_data = _T_data[_T_data__T_18_addr]; // @[Decoupled.scala 209:24]
  assign _T_data__T_10_data = io_enq_bits_data;
  assign _T_data__T_10_addr = value;
  assign _T_data__T_10_mask = 1'h1;
  assign _T_data__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_last__T_18_addr = value_1;
  assign _T_last__T_18_data = _T_last[_T_last__T_18_addr]; // @[Decoupled.scala 209:24]
  assign _T_last__T_10_data = io_enq_bits_last;
  assign _T_last__T_10_addr = value;
  assign _T_last__T_10_mask = 1'h1;
  assign _T_last__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_2 = value == value_1; // @[Decoupled.scala 214:41]
  assign _T_3 = ~_T_1; // @[Decoupled.scala 215:36]
  assign _T_4 = _T_2 & _T_3; // @[Decoupled.scala 215:33]
  assign _T_5 = _T_2 & _T_1; // @[Decoupled.scala 216:32]
  assign _T_6 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  assign _T_8 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  assign _T_12 = value + 1'h1; // @[Counter.scala 39:22]
  assign _T_14 = value_1 + 1'h1; // @[Counter.scala 39:22]
  assign _T_15 = _T_6 != _T_8; // @[Decoupled.scala 227:16]
  assign io_enq_ready = ~_T_5; // @[Decoupled.scala 232:16]
  assign io_deq_valid = ~_T_4; // @[Decoupled.scala 231:16]
  assign io_deq_bits_data = _T_data__T_18_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_last = _T_last__T_18_data; // @[Decoupled.scala 233:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_data[initvar] = _RAND_0[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_last[initvar] = _RAND_1[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  value = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  value_1 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T_data__T_10_en & _T_data__T_10_mask) begin
      _T_data[_T_data__T_10_addr] <= _T_data__T_10_data; // @[Decoupled.scala 209:24]
    end
    if(_T_last__T_10_en & _T_last__T_10_mask) begin
      _T_last[_T_last__T_10_addr] <= _T_last__T_10_data; // @[Decoupled.scala 209:24]
    end
    if (reset) begin
      value <= 1'h0;
    end else if (_T_6) begin
      value <= _T_12;
    end
    if (reset) begin
      value_1 <= 1'h0;
    end else if (_T_8) begin
      value_1 <= _T_14;
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else if (_T_15) begin
      _T_1 <= _T_6;
    end
  end
endmodule
module AXI4StreamBuffer_4(
  input         clock,
  input         reset,
  output        auto_in_ready,
  input         auto_in_valid,
  input  [31:0] auto_in_bits_data,
  input         auto_in_bits_last,
  input         auto_out_ready,
  output        auto_out_valid,
  output [31:0] auto_out_bits_data,
  output        auto_out_bits_last
);
  wire  Queue_clock; // @[Decoupled.scala 287:21]
  wire  Queue_reset; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_enq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_last; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_deq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_last; // @[Decoupled.scala 287:21]
  Queue_151 Queue ( // @[Decoupled.scala 287:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_last(Queue_io_enq_bits_last),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_last(Queue_io_deq_bits_last)
  );
  assign auto_in_ready = Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_out_valid = Queue_io_deq_valid; // @[LazyModule.scala 173:49]
  assign auto_out_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_bits_last = Queue_io_deq_bits_last; // @[LazyModule.scala 173:49]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_in_valid; // @[Decoupled.scala 288:22]
  assign Queue_io_enq_bits_data = auto_in_bits_data; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_last = auto_in_bits_last; // @[Decoupled.scala 289:21]
  assign Queue_io_deq_ready = auto_out_ready; // @[Decoupled.scala 311:15]
endmodule
module Queue_152(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [31:0] io_enq_bits_data,
  input         io_enq_bits_last,
  input         io_deq_ready,
  output        io_deq_valid,
  output [31:0] io_deq_bits_data,
  output        io_deq_bits_last
);
  reg [31:0] _T_data [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_0;
  wire [31:0] _T_data__T_18_data; // @[Decoupled.scala 209:24]
  wire  _T_data__T_18_addr; // @[Decoupled.scala 209:24]
  wire [31:0] _T_data__T_10_data; // @[Decoupled.scala 209:24]
  wire  _T_data__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T_data__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T_data__T_10_en; // @[Decoupled.scala 209:24]
  reg  _T_last [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_1;
  wire  _T_last__T_18_data; // @[Decoupled.scala 209:24]
  wire  _T_last__T_18_addr; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_data; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_en; // @[Decoupled.scala 209:24]
  reg  value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_2;
  reg  value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_3;
  reg  _T_1; // @[Decoupled.scala 212:35]
  reg [31:0] _RAND_4;
  wire  _T_2; // @[Decoupled.scala 214:41]
  wire  _T_3; // @[Decoupled.scala 215:36]
  wire  _T_4; // @[Decoupled.scala 215:33]
  wire  _T_5; // @[Decoupled.scala 216:32]
  wire  _T_6; // @[Decoupled.scala 40:37]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _T_12; // @[Counter.scala 39:22]
  wire  _T_14; // @[Counter.scala 39:22]
  wire  _T_15; // @[Decoupled.scala 227:16]
  assign _T_data__T_18_addr = value_1;
  assign _T_data__T_18_data = _T_data[_T_data__T_18_addr]; // @[Decoupled.scala 209:24]
  assign _T_data__T_10_data = io_enq_bits_data;
  assign _T_data__T_10_addr = value;
  assign _T_data__T_10_mask = 1'h1;
  assign _T_data__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_last__T_18_addr = value_1;
  assign _T_last__T_18_data = _T_last[_T_last__T_18_addr]; // @[Decoupled.scala 209:24]
  assign _T_last__T_10_data = io_enq_bits_last;
  assign _T_last__T_10_addr = value;
  assign _T_last__T_10_mask = 1'h1;
  assign _T_last__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_2 = value == value_1; // @[Decoupled.scala 214:41]
  assign _T_3 = ~_T_1; // @[Decoupled.scala 215:36]
  assign _T_4 = _T_2 & _T_3; // @[Decoupled.scala 215:33]
  assign _T_5 = _T_2 & _T_1; // @[Decoupled.scala 216:32]
  assign _T_6 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  assign _T_8 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  assign _T_12 = value + 1'h1; // @[Counter.scala 39:22]
  assign _T_14 = value_1 + 1'h1; // @[Counter.scala 39:22]
  assign _T_15 = _T_6 != _T_8; // @[Decoupled.scala 227:16]
  assign io_enq_ready = ~_T_5; // @[Decoupled.scala 232:16]
  assign io_deq_valid = ~_T_4; // @[Decoupled.scala 231:16]
  assign io_deq_bits_data = _T_data__T_18_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_last = _T_last__T_18_data; // @[Decoupled.scala 233:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_data[initvar] = _RAND_0[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_last[initvar] = _RAND_1[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  value = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  value_1 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T_data__T_10_en & _T_data__T_10_mask) begin
      _T_data[_T_data__T_10_addr] <= _T_data__T_10_data; // @[Decoupled.scala 209:24]
    end
    if(_T_last__T_10_en & _T_last__T_10_mask) begin
      _T_last[_T_last__T_10_addr] <= _T_last__T_10_data; // @[Decoupled.scala 209:24]
    end
    if (reset) begin
      value <= 1'h0;
    end else if (_T_6) begin
      value <= _T_12;
    end
    if (reset) begin
      value_1 <= 1'h0;
    end else if (_T_8) begin
      value_1 <= _T_14;
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else if (_T_15) begin
      _T_1 <= _T_6;
    end
  end
endmodule
module AXI4StreamBuffer_5(
  input         clock,
  input         reset,
  output        auto_in_ready,
  input         auto_in_valid,
  input  [31:0] auto_in_bits_data,
  input         auto_in_bits_last,
  input         auto_out_ready,
  output        auto_out_valid,
  output [31:0] auto_out_bits_data,
  output        auto_out_bits_last
);
  wire  Queue_clock; // @[Decoupled.scala 287:21]
  wire  Queue_reset; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_enq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_last; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_deq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_last; // @[Decoupled.scala 287:21]
  Queue_152 Queue ( // @[Decoupled.scala 287:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_last(Queue_io_enq_bits_last),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_last(Queue_io_deq_bits_last)
  );
  assign auto_in_ready = Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_out_valid = Queue_io_deq_valid; // @[LazyModule.scala 173:49]
  assign auto_out_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_bits_last = Queue_io_deq_bits_last; // @[LazyModule.scala 173:49]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_in_valid; // @[Decoupled.scala 288:22]
  assign Queue_io_enq_bits_data = auto_in_bits_data; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_last = auto_in_bits_last; // @[Decoupled.scala 289:21]
  assign Queue_io_deq_ready = auto_out_ready; // @[Decoupled.scala 311:15]
endmodule
module Queue_156(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [31:0] io_enq_bits_data,
  input         io_enq_bits_last,
  input         io_deq_ready,
  output        io_deq_valid,
  output [31:0] io_deq_bits_data,
  output        io_deq_bits_last
);
  reg [31:0] _T_data [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_0;
  wire [31:0] _T_data__T_18_data; // @[Decoupled.scala 209:24]
  wire  _T_data__T_18_addr; // @[Decoupled.scala 209:24]
  wire [31:0] _T_data__T_10_data; // @[Decoupled.scala 209:24]
  wire  _T_data__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T_data__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T_data__T_10_en; // @[Decoupled.scala 209:24]
  reg  _T_last [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_1;
  wire  _T_last__T_18_data; // @[Decoupled.scala 209:24]
  wire  _T_last__T_18_addr; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_data; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_en; // @[Decoupled.scala 209:24]
  reg  value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_2;
  reg  value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_3;
  reg  _T_1; // @[Decoupled.scala 212:35]
  reg [31:0] _RAND_4;
  wire  _T_2; // @[Decoupled.scala 214:41]
  wire  _T_3; // @[Decoupled.scala 215:36]
  wire  _T_4; // @[Decoupled.scala 215:33]
  wire  _T_5; // @[Decoupled.scala 216:32]
  wire  _T_6; // @[Decoupled.scala 40:37]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _T_12; // @[Counter.scala 39:22]
  wire  _T_14; // @[Counter.scala 39:22]
  wire  _T_15; // @[Decoupled.scala 227:16]
  assign _T_data__T_18_addr = value_1;
  assign _T_data__T_18_data = _T_data[_T_data__T_18_addr]; // @[Decoupled.scala 209:24]
  assign _T_data__T_10_data = io_enq_bits_data;
  assign _T_data__T_10_addr = value;
  assign _T_data__T_10_mask = 1'h1;
  assign _T_data__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_last__T_18_addr = value_1;
  assign _T_last__T_18_data = _T_last[_T_last__T_18_addr]; // @[Decoupled.scala 209:24]
  assign _T_last__T_10_data = io_enq_bits_last;
  assign _T_last__T_10_addr = value;
  assign _T_last__T_10_mask = 1'h1;
  assign _T_last__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_2 = value == value_1; // @[Decoupled.scala 214:41]
  assign _T_3 = ~_T_1; // @[Decoupled.scala 215:36]
  assign _T_4 = _T_2 & _T_3; // @[Decoupled.scala 215:33]
  assign _T_5 = _T_2 & _T_1; // @[Decoupled.scala 216:32]
  assign _T_6 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  assign _T_8 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  assign _T_12 = value + 1'h1; // @[Counter.scala 39:22]
  assign _T_14 = value_1 + 1'h1; // @[Counter.scala 39:22]
  assign _T_15 = _T_6 != _T_8; // @[Decoupled.scala 227:16]
  assign io_enq_ready = ~_T_5; // @[Decoupled.scala 232:16]
  assign io_deq_valid = ~_T_4; // @[Decoupled.scala 231:16]
  assign io_deq_bits_data = _T_data__T_18_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_last = _T_last__T_18_data; // @[Decoupled.scala 233:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_data[initvar] = _RAND_0[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_last[initvar] = _RAND_1[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  value = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  value_1 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T_data__T_10_en & _T_data__T_10_mask) begin
      _T_data[_T_data__T_10_addr] <= _T_data__T_10_data; // @[Decoupled.scala 209:24]
    end
    if(_T_last__T_10_en & _T_last__T_10_mask) begin
      _T_last[_T_last__T_10_addr] <= _T_last__T_10_data; // @[Decoupled.scala 209:24]
    end
    if (reset) begin
      value <= 1'h0;
    end else if (_T_6) begin
      value <= _T_12;
    end
    if (reset) begin
      value_1 <= 1'h0;
    end else if (_T_8) begin
      value_1 <= _T_14;
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else if (_T_15) begin
      _T_1 <= _T_6;
    end
  end
endmodule
module AXI4StreamBuffer_9(
  input         clock,
  input         reset,
  output        auto_in_ready,
  input         auto_in_valid,
  input  [31:0] auto_in_bits_data,
  input         auto_in_bits_last,
  input         auto_out_ready,
  output        auto_out_valid,
  output [31:0] auto_out_bits_data,
  output        auto_out_bits_last
);
  wire  Queue_clock; // @[Decoupled.scala 287:21]
  wire  Queue_reset; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_enq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_last; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_deq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_last; // @[Decoupled.scala 287:21]
  Queue_156 Queue ( // @[Decoupled.scala 287:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_last(Queue_io_enq_bits_last),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_last(Queue_io_deq_bits_last)
  );
  assign auto_in_ready = Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_out_valid = Queue_io_deq_valid; // @[LazyModule.scala 173:49]
  assign auto_out_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_bits_last = Queue_io_deq_bits_last; // @[LazyModule.scala 173:49]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_in_valid; // @[Decoupled.scala 288:22]
  assign Queue_io_enq_bits_data = auto_in_bits_data; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_last = auto_in_bits_last; // @[Decoupled.scala 289:21]
  assign Queue_io_deq_ready = auto_out_ready; // @[Decoupled.scala 311:15]
endmodule
module BundleBridgeToAXI4(
  output        auto_in_aw_ready,
  input         auto_in_aw_valid,
  input         auto_in_aw_bits_id,
  input  [31:0] auto_in_aw_bits_addr,
  input  [2:0]  auto_in_aw_bits_size,
  output        auto_in_w_ready,
  input         auto_in_w_valid,
  input  [31:0] auto_in_w_bits_data,
  input  [3:0]  auto_in_w_bits_strb,
  input         auto_in_w_bits_last,
  input         auto_in_b_ready,
  output        auto_in_b_valid,
  output [1:0]  auto_in_b_bits_resp,
  output        auto_in_ar_ready,
  input         auto_in_ar_valid,
  input         auto_in_ar_bits_id,
  input  [31:0] auto_in_ar_bits_addr,
  input  [2:0]  auto_in_ar_bits_size,
  input         auto_in_r_ready,
  output        auto_in_r_valid,
  output [31:0] auto_in_r_bits_data,
  output [1:0]  auto_in_r_bits_resp,
  output        auto_in_r_bits_last,
  input         auto_out_aw_ready,
  output        auto_out_aw_valid,
  output        auto_out_aw_bits_id,
  output [29:0] auto_out_aw_bits_addr,
  output [2:0]  auto_out_aw_bits_size,
  input         auto_out_w_ready,
  output        auto_out_w_valid,
  output [31:0] auto_out_w_bits_data,
  output [3:0]  auto_out_w_bits_strb,
  output        auto_out_w_bits_last,
  output        auto_out_b_ready,
  input         auto_out_b_valid,
  input  [1:0]  auto_out_b_bits_resp,
  input         auto_out_ar_ready,
  output        auto_out_ar_valid,
  output        auto_out_ar_bits_id,
  output [29:0] auto_out_ar_bits_addr,
  output [2:0]  auto_out_ar_bits_size,
  output        auto_out_r_ready,
  input         auto_out_r_valid,
  input  [31:0] auto_out_r_bits_data,
  input  [1:0]  auto_out_r_bits_resp,
  input         auto_out_r_bits_last
);
  assign auto_in_aw_ready = auto_out_aw_ready; // @[LazyModule.scala 173:31]
  assign auto_in_w_ready = auto_out_w_ready; // @[LazyModule.scala 173:31]
  assign auto_in_b_valid = auto_out_b_valid; // @[LazyModule.scala 173:31]
  assign auto_in_b_bits_resp = auto_out_b_bits_resp; // @[LazyModule.scala 173:31]
  assign auto_in_ar_ready = auto_out_ar_ready; // @[LazyModule.scala 173:31]
  assign auto_in_r_valid = auto_out_r_valid; // @[LazyModule.scala 173:31]
  assign auto_in_r_bits_data = auto_out_r_bits_data; // @[LazyModule.scala 173:31]
  assign auto_in_r_bits_resp = auto_out_r_bits_resp; // @[LazyModule.scala 173:31]
  assign auto_in_r_bits_last = auto_out_r_bits_last; // @[LazyModule.scala 173:31]
  assign auto_out_aw_valid = auto_in_aw_valid; // @[LazyModule.scala 173:49]
  assign auto_out_aw_bits_id = auto_in_aw_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_aw_bits_addr = auto_in_aw_bits_addr[29:0]; // @[LazyModule.scala 173:49]
  assign auto_out_aw_bits_size = auto_in_aw_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_w_valid = auto_in_w_valid; // @[LazyModule.scala 173:49]
  assign auto_out_w_bits_data = auto_in_w_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_w_bits_strb = auto_in_w_bits_strb; // @[LazyModule.scala 173:49]
  assign auto_out_w_bits_last = auto_in_w_bits_last; // @[LazyModule.scala 173:49]
  assign auto_out_b_ready = auto_in_b_ready; // @[LazyModule.scala 173:49]
  assign auto_out_ar_valid = auto_in_ar_valid; // @[LazyModule.scala 173:49]
  assign auto_out_ar_bits_id = auto_in_ar_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_ar_bits_addr = auto_in_ar_bits_addr[29:0]; // @[LazyModule.scala 173:49]
  assign auto_out_ar_bits_size = auto_in_ar_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_r_ready = auto_in_r_ready; // @[LazyModule.scala 173:49]
endmodule
module AXI4StreamToBundleBridge(
  output       auto_in_ready,
  input        auto_in_valid,
  input  [7:0] auto_in_bits_data,
  input        auto_in_bits_last,
  input        auto_out_ready,
  output       auto_out_valid,
  output [7:0] auto_out_bits_data,
  output       auto_out_bits_last
);
  assign auto_in_ready = auto_out_ready; // @[LazyModule.scala 173:31]
  assign auto_out_valid = auto_in_valid; // @[LazyModule.scala 173:49]
  assign auto_out_bits_data = auto_in_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_bits_last = auto_in_bits_last; // @[LazyModule.scala 173:49]
endmodule
module SpectrometerTestWithoutLA(
  input         clock,
  input         reset,
  output        ioMem_0_aw_ready,
  input         ioMem_0_aw_valid,
  input         ioMem_0_aw_bits_id,
  input  [31:0] ioMem_0_aw_bits_addr,
  input  [7:0]  ioMem_0_aw_bits_len,
  input  [2:0]  ioMem_0_aw_bits_size,
  input  [1:0]  ioMem_0_aw_bits_burst,
  input         ioMem_0_aw_bits_lock,
  input  [3:0]  ioMem_0_aw_bits_cache,
  input  [2:0]  ioMem_0_aw_bits_prot,
  input  [3:0]  ioMem_0_aw_bits_qos,
  output        ioMem_0_w_ready,
  input         ioMem_0_w_valid,
  input  [31:0] ioMem_0_w_bits_data,
  input  [3:0]  ioMem_0_w_bits_strb,
  input         ioMem_0_w_bits_last,
  input         ioMem_0_b_ready,
  output        ioMem_0_b_valid,
  output        ioMem_0_b_bits_id,
  output [1:0]  ioMem_0_b_bits_resp,
  output        ioMem_0_ar_ready,
  input         ioMem_0_ar_valid,
  input         ioMem_0_ar_bits_id,
  input  [31:0] ioMem_0_ar_bits_addr,
  input  [7:0]  ioMem_0_ar_bits_len,
  input  [2:0]  ioMem_0_ar_bits_size,
  input  [1:0]  ioMem_0_ar_bits_burst,
  input         ioMem_0_ar_bits_lock,
  input  [3:0]  ioMem_0_ar_bits_cache,
  input  [2:0]  ioMem_0_ar_bits_prot,
  input  [3:0]  ioMem_0_ar_bits_qos,
  input         ioMem_0_r_ready,
  output        ioMem_0_r_valid,
  output        ioMem_0_r_bits_id,
  output [31:0] ioMem_0_r_bits_data,
  output [1:0]  ioMem_0_r_bits_resp,
  output        ioMem_0_r_bits_last,
  input         outStream_0_ready,
  output        outStream_0_valid,
  output [7:0]  outStream_0_bits_data,
  output        outStream_0_bits_last,
  output        inStream_0_ready,
  input         inStream_0_valid,
  input  [7:0]  inStream_0_bits_data,
  input         inStream_0_bits_last,
  output        int_0,
  output        uTx,
  input         uRx
);
  wire  widthAdapter_clock; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_reset; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_auto_in_ready; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_auto_in_valid; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire [7:0] widthAdapter_auto_in_bits_data; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_auto_in_bits_last; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_auto_out_ready; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_auto_out_valid; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire [31:0] widthAdapter_auto_out_bits_data; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_auto_out_bits_last; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  in_split_clock; // @[SpectrometerTestWithoutLA.scala 59:29]
  wire  in_split_reset; // @[SpectrometerTestWithoutLA.scala 59:29]
  wire  in_split_auto_mem_in_aw_ready; // @[SpectrometerTestWithoutLA.scala 59:29]
  wire  in_split_auto_mem_in_aw_valid; // @[SpectrometerTestWithoutLA.scala 59:29]
  wire  in_split_auto_mem_in_aw_bits_id; // @[SpectrometerTestWithoutLA.scala 59:29]
  wire [29:0] in_split_auto_mem_in_aw_bits_addr; // @[SpectrometerTestWithoutLA.scala 59:29]
  wire  in_split_auto_mem_in_w_ready; // @[SpectrometerTestWithoutLA.scala 59:29]
  wire  in_split_auto_mem_in_w_valid; // @[SpectrometerTestWithoutLA.scala 59:29]
  wire [31:0] in_split_auto_mem_in_w_bits_data; // @[SpectrometerTestWithoutLA.scala 59:29]
  wire [3:0] in_split_auto_mem_in_w_bits_strb; // @[SpectrometerTestWithoutLA.scala 59:29]
  wire  in_split_auto_mem_in_b_ready; // @[SpectrometerTestWithoutLA.scala 59:29]
  wire  in_split_auto_mem_in_b_valid; // @[SpectrometerTestWithoutLA.scala 59:29]
  wire  in_split_auto_mem_in_b_bits_id; // @[SpectrometerTestWithoutLA.scala 59:29]
  wire  in_split_auto_mem_in_ar_ready; // @[SpectrometerTestWithoutLA.scala 59:29]
  wire  in_split_auto_mem_in_ar_valid; // @[SpectrometerTestWithoutLA.scala 59:29]
  wire  in_split_auto_mem_in_ar_bits_id; // @[SpectrometerTestWithoutLA.scala 59:29]
  wire [29:0] in_split_auto_mem_in_ar_bits_addr; // @[SpectrometerTestWithoutLA.scala 59:29]
  wire [2:0] in_split_auto_mem_in_ar_bits_size; // @[SpectrometerTestWithoutLA.scala 59:29]
  wire  in_split_auto_mem_in_r_ready; // @[SpectrometerTestWithoutLA.scala 59:29]
  wire  in_split_auto_mem_in_r_valid; // @[SpectrometerTestWithoutLA.scala 59:29]
  wire  in_split_auto_mem_in_r_bits_id; // @[SpectrometerTestWithoutLA.scala 59:29]
  wire [31:0] in_split_auto_mem_in_r_bits_data; // @[SpectrometerTestWithoutLA.scala 59:29]
  wire  in_split_auto_stream_in_ready; // @[SpectrometerTestWithoutLA.scala 59:29]
  wire  in_split_auto_stream_in_valid; // @[SpectrometerTestWithoutLA.scala 59:29]
  wire [31:0] in_split_auto_stream_in_bits_data; // @[SpectrometerTestWithoutLA.scala 59:29]
  wire  in_split_auto_stream_in_bits_last; // @[SpectrometerTestWithoutLA.scala 59:29]
  wire  in_split_auto_stream_out_4_ready; // @[SpectrometerTestWithoutLA.scala 59:29]
  wire  in_split_auto_stream_out_4_valid; // @[SpectrometerTestWithoutLA.scala 59:29]
  wire [31:0] in_split_auto_stream_out_4_bits_data; // @[SpectrometerTestWithoutLA.scala 59:29]
  wire  in_split_auto_stream_out_4_bits_last; // @[SpectrometerTestWithoutLA.scala 59:29]
  wire  in_split_auto_stream_out_3_ready; // @[SpectrometerTestWithoutLA.scala 59:29]
  wire  in_split_auto_stream_out_3_valid; // @[SpectrometerTestWithoutLA.scala 59:29]
  wire [31:0] in_split_auto_stream_out_3_bits_data; // @[SpectrometerTestWithoutLA.scala 59:29]
  wire  in_split_auto_stream_out_3_bits_last; // @[SpectrometerTestWithoutLA.scala 59:29]
  wire  in_split_auto_stream_out_2_ready; // @[SpectrometerTestWithoutLA.scala 59:29]
  wire  in_split_auto_stream_out_2_valid; // @[SpectrometerTestWithoutLA.scala 59:29]
  wire [31:0] in_split_auto_stream_out_2_bits_data; // @[SpectrometerTestWithoutLA.scala 59:29]
  wire  in_split_auto_stream_out_2_bits_last; // @[SpectrometerTestWithoutLA.scala 59:29]
  wire  in_split_auto_stream_out_1_ready; // @[SpectrometerTestWithoutLA.scala 59:29]
  wire  in_split_auto_stream_out_1_valid; // @[SpectrometerTestWithoutLA.scala 59:29]
  wire [31:0] in_split_auto_stream_out_1_bits_data; // @[SpectrometerTestWithoutLA.scala 59:29]
  wire  in_split_auto_stream_out_1_bits_last; // @[SpectrometerTestWithoutLA.scala 59:29]
  wire  in_split_auto_stream_out_0_ready; // @[SpectrometerTestWithoutLA.scala 59:29]
  wire  in_split_auto_stream_out_0_valid; // @[SpectrometerTestWithoutLA.scala 59:29]
  wire [31:0] in_split_auto_stream_out_0_bits_data; // @[SpectrometerTestWithoutLA.scala 59:29]
  wire  in_split_auto_stream_out_0_bits_last; // @[SpectrometerTestWithoutLA.scala 59:29]
  wire  in_queue_clock; // @[SpectrometerTestWithoutLA.scala 60:29]
  wire  in_queue_reset; // @[SpectrometerTestWithoutLA.scala 60:29]
  wire  in_queue_auto_out_out_ready; // @[SpectrometerTestWithoutLA.scala 60:29]
  wire  in_queue_auto_out_out_valid; // @[SpectrometerTestWithoutLA.scala 60:29]
  wire [7:0] in_queue_auto_out_out_bits_data; // @[SpectrometerTestWithoutLA.scala 60:29]
  wire  in_queue_auto_out_out_bits_last; // @[SpectrometerTestWithoutLA.scala 60:29]
  wire  in_queue_auto_in_in_ready; // @[SpectrometerTestWithoutLA.scala 60:29]
  wire  in_queue_auto_in_in_valid; // @[SpectrometerTestWithoutLA.scala 60:29]
  wire [7:0] in_queue_auto_in_in_bits_data; // @[SpectrometerTestWithoutLA.scala 60:29]
  wire  in_queue_auto_in_in_bits_last; // @[SpectrometerTestWithoutLA.scala 60:29]
  wire  plfg_clock; // @[SpectrometerTestWithoutLA.scala 62:30]
  wire  plfg_reset; // @[SpectrometerTestWithoutLA.scala 62:30]
  wire  plfg_auto_mem_in_aw_ready; // @[SpectrometerTestWithoutLA.scala 62:30]
  wire  plfg_auto_mem_in_aw_valid; // @[SpectrometerTestWithoutLA.scala 62:30]
  wire  plfg_auto_mem_in_aw_bits_id; // @[SpectrometerTestWithoutLA.scala 62:30]
  wire [29:0] plfg_auto_mem_in_aw_bits_addr; // @[SpectrometerTestWithoutLA.scala 62:30]
  wire  plfg_auto_mem_in_w_ready; // @[SpectrometerTestWithoutLA.scala 62:30]
  wire  plfg_auto_mem_in_w_valid; // @[SpectrometerTestWithoutLA.scala 62:30]
  wire [31:0] plfg_auto_mem_in_w_bits_data; // @[SpectrometerTestWithoutLA.scala 62:30]
  wire [3:0] plfg_auto_mem_in_w_bits_strb; // @[SpectrometerTestWithoutLA.scala 62:30]
  wire  plfg_auto_mem_in_w_bits_last; // @[SpectrometerTestWithoutLA.scala 62:30]
  wire  plfg_auto_mem_in_b_ready; // @[SpectrometerTestWithoutLA.scala 62:30]
  wire  plfg_auto_mem_in_b_valid; // @[SpectrometerTestWithoutLA.scala 62:30]
  wire [1:0] plfg_auto_mem_in_b_bits_resp; // @[SpectrometerTestWithoutLA.scala 62:30]
  wire  plfg_auto_mem_in_ar_ready; // @[SpectrometerTestWithoutLA.scala 62:30]
  wire  plfg_auto_mem_in_ar_valid; // @[SpectrometerTestWithoutLA.scala 62:30]
  wire  plfg_auto_mem_in_ar_bits_id; // @[SpectrometerTestWithoutLA.scala 62:30]
  wire [29:0] plfg_auto_mem_in_ar_bits_addr; // @[SpectrometerTestWithoutLA.scala 62:30]
  wire [2:0] plfg_auto_mem_in_ar_bits_size; // @[SpectrometerTestWithoutLA.scala 62:30]
  wire  plfg_auto_mem_in_r_ready; // @[SpectrometerTestWithoutLA.scala 62:30]
  wire  plfg_auto_mem_in_r_valid; // @[SpectrometerTestWithoutLA.scala 62:30]
  wire [31:0] plfg_auto_mem_in_r_bits_data; // @[SpectrometerTestWithoutLA.scala 62:30]
  wire [1:0] plfg_auto_mem_in_r_bits_resp; // @[SpectrometerTestWithoutLA.scala 62:30]
  wire  plfg_auto_mem_in_r_bits_last; // @[SpectrometerTestWithoutLA.scala 62:30]
  wire  plfg_auto_stream_out_ready; // @[SpectrometerTestWithoutLA.scala 62:30]
  wire  plfg_auto_stream_out_valid; // @[SpectrometerTestWithoutLA.scala 62:30]
  wire [31:0] plfg_auto_stream_out_bits_data; // @[SpectrometerTestWithoutLA.scala 62:30]
  wire  plfg_auto_stream_out_bits_last; // @[SpectrometerTestWithoutLA.scala 62:30]
  wire  plfg_split_clock; // @[SpectrometerTestWithoutLA.scala 63:30]
  wire  plfg_split_reset; // @[SpectrometerTestWithoutLA.scala 63:30]
  wire  plfg_split_auto_mem_in_aw_ready; // @[SpectrometerTestWithoutLA.scala 63:30]
  wire  plfg_split_auto_mem_in_aw_valid; // @[SpectrometerTestWithoutLA.scala 63:30]
  wire  plfg_split_auto_mem_in_aw_bits_id; // @[SpectrometerTestWithoutLA.scala 63:30]
  wire [29:0] plfg_split_auto_mem_in_aw_bits_addr; // @[SpectrometerTestWithoutLA.scala 63:30]
  wire  plfg_split_auto_mem_in_w_ready; // @[SpectrometerTestWithoutLA.scala 63:30]
  wire  plfg_split_auto_mem_in_w_valid; // @[SpectrometerTestWithoutLA.scala 63:30]
  wire [31:0] plfg_split_auto_mem_in_w_bits_data; // @[SpectrometerTestWithoutLA.scala 63:30]
  wire [3:0] plfg_split_auto_mem_in_w_bits_strb; // @[SpectrometerTestWithoutLA.scala 63:30]
  wire  plfg_split_auto_mem_in_b_ready; // @[SpectrometerTestWithoutLA.scala 63:30]
  wire  plfg_split_auto_mem_in_b_valid; // @[SpectrometerTestWithoutLA.scala 63:30]
  wire  plfg_split_auto_mem_in_b_bits_id; // @[SpectrometerTestWithoutLA.scala 63:30]
  wire  plfg_split_auto_mem_in_ar_ready; // @[SpectrometerTestWithoutLA.scala 63:30]
  wire  plfg_split_auto_mem_in_ar_valid; // @[SpectrometerTestWithoutLA.scala 63:30]
  wire  plfg_split_auto_mem_in_ar_bits_id; // @[SpectrometerTestWithoutLA.scala 63:30]
  wire [29:0] plfg_split_auto_mem_in_ar_bits_addr; // @[SpectrometerTestWithoutLA.scala 63:30]
  wire [2:0] plfg_split_auto_mem_in_ar_bits_size; // @[SpectrometerTestWithoutLA.scala 63:30]
  wire  plfg_split_auto_mem_in_r_ready; // @[SpectrometerTestWithoutLA.scala 63:30]
  wire  plfg_split_auto_mem_in_r_valid; // @[SpectrometerTestWithoutLA.scala 63:30]
  wire  plfg_split_auto_mem_in_r_bits_id; // @[SpectrometerTestWithoutLA.scala 63:30]
  wire [31:0] plfg_split_auto_mem_in_r_bits_data; // @[SpectrometerTestWithoutLA.scala 63:30]
  wire  plfg_split_auto_stream_in_ready; // @[SpectrometerTestWithoutLA.scala 63:30]
  wire  plfg_split_auto_stream_in_valid; // @[SpectrometerTestWithoutLA.scala 63:30]
  wire [31:0] plfg_split_auto_stream_in_bits_data; // @[SpectrometerTestWithoutLA.scala 63:30]
  wire  plfg_split_auto_stream_in_bits_last; // @[SpectrometerTestWithoutLA.scala 63:30]
  wire  plfg_split_auto_stream_out_1_ready; // @[SpectrometerTestWithoutLA.scala 63:30]
  wire  plfg_split_auto_stream_out_1_valid; // @[SpectrometerTestWithoutLA.scala 63:30]
  wire [31:0] plfg_split_auto_stream_out_1_bits_data; // @[SpectrometerTestWithoutLA.scala 63:30]
  wire  plfg_split_auto_stream_out_1_bits_last; // @[SpectrometerTestWithoutLA.scala 63:30]
  wire  plfg_split_auto_stream_out_0_ready; // @[SpectrometerTestWithoutLA.scala 63:30]
  wire  plfg_split_auto_stream_out_0_valid; // @[SpectrometerTestWithoutLA.scala 63:30]
  wire [31:0] plfg_split_auto_stream_out_0_bits_data; // @[SpectrometerTestWithoutLA.scala 63:30]
  wire  plfg_split_auto_stream_out_0_bits_last; // @[SpectrometerTestWithoutLA.scala 63:30]
  wire  plfg_mux_0_clock; // @[SpectrometerTestWithoutLA.scala 64:30]
  wire  plfg_mux_0_reset; // @[SpectrometerTestWithoutLA.scala 64:30]
  wire  plfg_mux_0_auto_register_in_aw_ready; // @[SpectrometerTestWithoutLA.scala 64:30]
  wire  plfg_mux_0_auto_register_in_aw_valid; // @[SpectrometerTestWithoutLA.scala 64:30]
  wire  plfg_mux_0_auto_register_in_aw_bits_id; // @[SpectrometerTestWithoutLA.scala 64:30]
  wire [29:0] plfg_mux_0_auto_register_in_aw_bits_addr; // @[SpectrometerTestWithoutLA.scala 64:30]
  wire  plfg_mux_0_auto_register_in_w_ready; // @[SpectrometerTestWithoutLA.scala 64:30]
  wire  plfg_mux_0_auto_register_in_w_valid; // @[SpectrometerTestWithoutLA.scala 64:30]
  wire [31:0] plfg_mux_0_auto_register_in_w_bits_data; // @[SpectrometerTestWithoutLA.scala 64:30]
  wire [3:0] plfg_mux_0_auto_register_in_w_bits_strb; // @[SpectrometerTestWithoutLA.scala 64:30]
  wire  plfg_mux_0_auto_register_in_b_ready; // @[SpectrometerTestWithoutLA.scala 64:30]
  wire  plfg_mux_0_auto_register_in_b_valid; // @[SpectrometerTestWithoutLA.scala 64:30]
  wire  plfg_mux_0_auto_register_in_b_bits_id; // @[SpectrometerTestWithoutLA.scala 64:30]
  wire  plfg_mux_0_auto_register_in_ar_ready; // @[SpectrometerTestWithoutLA.scala 64:30]
  wire  plfg_mux_0_auto_register_in_ar_valid; // @[SpectrometerTestWithoutLA.scala 64:30]
  wire  plfg_mux_0_auto_register_in_ar_bits_id; // @[SpectrometerTestWithoutLA.scala 64:30]
  wire [29:0] plfg_mux_0_auto_register_in_ar_bits_addr; // @[SpectrometerTestWithoutLA.scala 64:30]
  wire [2:0] plfg_mux_0_auto_register_in_ar_bits_size; // @[SpectrometerTestWithoutLA.scala 64:30]
  wire  plfg_mux_0_auto_register_in_r_ready; // @[SpectrometerTestWithoutLA.scala 64:30]
  wire  plfg_mux_0_auto_register_in_r_valid; // @[SpectrometerTestWithoutLA.scala 64:30]
  wire  plfg_mux_0_auto_register_in_r_bits_id; // @[SpectrometerTestWithoutLA.scala 64:30]
  wire [31:0] plfg_mux_0_auto_register_in_r_bits_data; // @[SpectrometerTestWithoutLA.scala 64:30]
  wire  plfg_mux_0_auto_stream_in_2_ready; // @[SpectrometerTestWithoutLA.scala 64:30]
  wire  plfg_mux_0_auto_stream_in_2_valid; // @[SpectrometerTestWithoutLA.scala 64:30]
  wire [31:0] plfg_mux_0_auto_stream_in_2_bits_data; // @[SpectrometerTestWithoutLA.scala 64:30]
  wire  plfg_mux_0_auto_stream_in_2_bits_last; // @[SpectrometerTestWithoutLA.scala 64:30]
  wire  plfg_mux_0_auto_stream_in_1_ready; // @[SpectrometerTestWithoutLA.scala 64:30]
  wire  plfg_mux_0_auto_stream_in_1_valid; // @[SpectrometerTestWithoutLA.scala 64:30]
  wire [31:0] plfg_mux_0_auto_stream_in_1_bits_data; // @[SpectrometerTestWithoutLA.scala 64:30]
  wire  plfg_mux_0_auto_stream_in_1_bits_last; // @[SpectrometerTestWithoutLA.scala 64:30]
  wire  plfg_mux_0_auto_stream_in_0_ready; // @[SpectrometerTestWithoutLA.scala 64:30]
  wire  plfg_mux_0_auto_stream_in_0_valid; // @[SpectrometerTestWithoutLA.scala 64:30]
  wire [31:0] plfg_mux_0_auto_stream_in_0_bits_data; // @[SpectrometerTestWithoutLA.scala 64:30]
  wire  plfg_mux_0_auto_stream_in_0_bits_last; // @[SpectrometerTestWithoutLA.scala 64:30]
  wire  plfg_mux_0_auto_stream_out_0_ready; // @[SpectrometerTestWithoutLA.scala 64:30]
  wire  plfg_mux_0_auto_stream_out_0_valid; // @[SpectrometerTestWithoutLA.scala 64:30]
  wire [31:0] plfg_mux_0_auto_stream_out_0_bits_data; // @[SpectrometerTestWithoutLA.scala 64:30]
  wire  plfg_mux_0_auto_stream_out_0_bits_last; // @[SpectrometerTestWithoutLA.scala 64:30]
  wire  plfg_mux_1_clock; // @[SpectrometerTestWithoutLA.scala 65:30]
  wire  plfg_mux_1_reset; // @[SpectrometerTestWithoutLA.scala 65:30]
  wire  plfg_mux_1_auto_register_in_aw_ready; // @[SpectrometerTestWithoutLA.scala 65:30]
  wire  plfg_mux_1_auto_register_in_aw_valid; // @[SpectrometerTestWithoutLA.scala 65:30]
  wire  plfg_mux_1_auto_register_in_aw_bits_id; // @[SpectrometerTestWithoutLA.scala 65:30]
  wire [29:0] plfg_mux_1_auto_register_in_aw_bits_addr; // @[SpectrometerTestWithoutLA.scala 65:30]
  wire  plfg_mux_1_auto_register_in_w_ready; // @[SpectrometerTestWithoutLA.scala 65:30]
  wire  plfg_mux_1_auto_register_in_w_valid; // @[SpectrometerTestWithoutLA.scala 65:30]
  wire [31:0] plfg_mux_1_auto_register_in_w_bits_data; // @[SpectrometerTestWithoutLA.scala 65:30]
  wire [3:0] plfg_mux_1_auto_register_in_w_bits_strb; // @[SpectrometerTestWithoutLA.scala 65:30]
  wire  plfg_mux_1_auto_register_in_b_ready; // @[SpectrometerTestWithoutLA.scala 65:30]
  wire  plfg_mux_1_auto_register_in_b_valid; // @[SpectrometerTestWithoutLA.scala 65:30]
  wire  plfg_mux_1_auto_register_in_b_bits_id; // @[SpectrometerTestWithoutLA.scala 65:30]
  wire  plfg_mux_1_auto_register_in_ar_ready; // @[SpectrometerTestWithoutLA.scala 65:30]
  wire  plfg_mux_1_auto_register_in_ar_valid; // @[SpectrometerTestWithoutLA.scala 65:30]
  wire  plfg_mux_1_auto_register_in_ar_bits_id; // @[SpectrometerTestWithoutLA.scala 65:30]
  wire [29:0] plfg_mux_1_auto_register_in_ar_bits_addr; // @[SpectrometerTestWithoutLA.scala 65:30]
  wire [2:0] plfg_mux_1_auto_register_in_ar_bits_size; // @[SpectrometerTestWithoutLA.scala 65:30]
  wire  plfg_mux_1_auto_register_in_r_ready; // @[SpectrometerTestWithoutLA.scala 65:30]
  wire  plfg_mux_1_auto_register_in_r_valid; // @[SpectrometerTestWithoutLA.scala 65:30]
  wire  plfg_mux_1_auto_register_in_r_bits_id; // @[SpectrometerTestWithoutLA.scala 65:30]
  wire [31:0] plfg_mux_1_auto_register_in_r_bits_data; // @[SpectrometerTestWithoutLA.scala 65:30]
  wire  plfg_mux_1_auto_stream_in_ready; // @[SpectrometerTestWithoutLA.scala 65:30]
  wire  plfg_mux_1_auto_stream_in_valid; // @[SpectrometerTestWithoutLA.scala 65:30]
  wire [31:0] plfg_mux_1_auto_stream_in_bits_data; // @[SpectrometerTestWithoutLA.scala 65:30]
  wire  plfg_mux_1_auto_stream_in_bits_last; // @[SpectrometerTestWithoutLA.scala 65:30]
  wire  plfg_mux_1_auto_stream_out_1_ready; // @[SpectrometerTestWithoutLA.scala 65:30]
  wire  plfg_mux_1_auto_stream_out_1_valid; // @[SpectrometerTestWithoutLA.scala 65:30]
  wire [31:0] plfg_mux_1_auto_stream_out_1_bits_data; // @[SpectrometerTestWithoutLA.scala 65:30]
  wire  plfg_mux_1_auto_stream_out_1_bits_last; // @[SpectrometerTestWithoutLA.scala 65:30]
  wire  nco_clock; // @[SpectrometerTestWithoutLA.scala 71:29]
  wire  nco_reset; // @[SpectrometerTestWithoutLA.scala 71:29]
  wire  nco_auto_stream_out_ready; // @[SpectrometerTestWithoutLA.scala 71:29]
  wire  nco_auto_stream_out_valid; // @[SpectrometerTestWithoutLA.scala 71:29]
  wire [31:0] nco_auto_stream_out_bits_data; // @[SpectrometerTestWithoutLA.scala 71:29]
  wire  nco_auto_stream_out_bits_last; // @[SpectrometerTestWithoutLA.scala 71:29]
  wire  nco_auto_freq_in_ready; // @[SpectrometerTestWithoutLA.scala 71:29]
  wire  nco_auto_freq_in_valid; // @[SpectrometerTestWithoutLA.scala 71:29]
  wire [31:0] nco_auto_freq_in_bits_data; // @[SpectrometerTestWithoutLA.scala 71:29]
  wire  nco_auto_freq_in_bits_last; // @[SpectrometerTestWithoutLA.scala 71:29]
  wire  nco_split_clock; // @[SpectrometerTestWithoutLA.scala 72:29]
  wire  nco_split_reset; // @[SpectrometerTestWithoutLA.scala 72:29]
  wire  nco_split_auto_mem_in_aw_ready; // @[SpectrometerTestWithoutLA.scala 72:29]
  wire  nco_split_auto_mem_in_aw_valid; // @[SpectrometerTestWithoutLA.scala 72:29]
  wire  nco_split_auto_mem_in_aw_bits_id; // @[SpectrometerTestWithoutLA.scala 72:29]
  wire [29:0] nco_split_auto_mem_in_aw_bits_addr; // @[SpectrometerTestWithoutLA.scala 72:29]
  wire  nco_split_auto_mem_in_w_ready; // @[SpectrometerTestWithoutLA.scala 72:29]
  wire  nco_split_auto_mem_in_w_valid; // @[SpectrometerTestWithoutLA.scala 72:29]
  wire [31:0] nco_split_auto_mem_in_w_bits_data; // @[SpectrometerTestWithoutLA.scala 72:29]
  wire [3:0] nco_split_auto_mem_in_w_bits_strb; // @[SpectrometerTestWithoutLA.scala 72:29]
  wire  nco_split_auto_mem_in_b_ready; // @[SpectrometerTestWithoutLA.scala 72:29]
  wire  nco_split_auto_mem_in_b_valid; // @[SpectrometerTestWithoutLA.scala 72:29]
  wire  nco_split_auto_mem_in_b_bits_id; // @[SpectrometerTestWithoutLA.scala 72:29]
  wire  nco_split_auto_mem_in_ar_ready; // @[SpectrometerTestWithoutLA.scala 72:29]
  wire  nco_split_auto_mem_in_ar_valid; // @[SpectrometerTestWithoutLA.scala 72:29]
  wire  nco_split_auto_mem_in_ar_bits_id; // @[SpectrometerTestWithoutLA.scala 72:29]
  wire [29:0] nco_split_auto_mem_in_ar_bits_addr; // @[SpectrometerTestWithoutLA.scala 72:29]
  wire [2:0] nco_split_auto_mem_in_ar_bits_size; // @[SpectrometerTestWithoutLA.scala 72:29]
  wire  nco_split_auto_mem_in_r_ready; // @[SpectrometerTestWithoutLA.scala 72:29]
  wire  nco_split_auto_mem_in_r_valid; // @[SpectrometerTestWithoutLA.scala 72:29]
  wire  nco_split_auto_mem_in_r_bits_id; // @[SpectrometerTestWithoutLA.scala 72:29]
  wire [31:0] nco_split_auto_mem_in_r_bits_data; // @[SpectrometerTestWithoutLA.scala 72:29]
  wire  nco_split_auto_stream_in_ready; // @[SpectrometerTestWithoutLA.scala 72:29]
  wire  nco_split_auto_stream_in_valid; // @[SpectrometerTestWithoutLA.scala 72:29]
  wire [31:0] nco_split_auto_stream_in_bits_data; // @[SpectrometerTestWithoutLA.scala 72:29]
  wire  nco_split_auto_stream_in_bits_last; // @[SpectrometerTestWithoutLA.scala 72:29]
  wire  nco_split_auto_stream_out_1_ready; // @[SpectrometerTestWithoutLA.scala 72:29]
  wire  nco_split_auto_stream_out_1_valid; // @[SpectrometerTestWithoutLA.scala 72:29]
  wire [31:0] nco_split_auto_stream_out_1_bits_data; // @[SpectrometerTestWithoutLA.scala 72:29]
  wire  nco_split_auto_stream_out_1_bits_last; // @[SpectrometerTestWithoutLA.scala 72:29]
  wire  nco_split_auto_stream_out_0_ready; // @[SpectrometerTestWithoutLA.scala 72:29]
  wire  nco_split_auto_stream_out_0_valid; // @[SpectrometerTestWithoutLA.scala 72:29]
  wire [31:0] nco_split_auto_stream_out_0_bits_data; // @[SpectrometerTestWithoutLA.scala 72:29]
  wire  nco_split_auto_stream_out_0_bits_last; // @[SpectrometerTestWithoutLA.scala 72:29]
  wire  nco_mux_0_clock; // @[SpectrometerTestWithoutLA.scala 73:29]
  wire  nco_mux_0_reset; // @[SpectrometerTestWithoutLA.scala 73:29]
  wire  nco_mux_0_auto_register_in_aw_ready; // @[SpectrometerTestWithoutLA.scala 73:29]
  wire  nco_mux_0_auto_register_in_aw_valid; // @[SpectrometerTestWithoutLA.scala 73:29]
  wire  nco_mux_0_auto_register_in_aw_bits_id; // @[SpectrometerTestWithoutLA.scala 73:29]
  wire [29:0] nco_mux_0_auto_register_in_aw_bits_addr; // @[SpectrometerTestWithoutLA.scala 73:29]
  wire  nco_mux_0_auto_register_in_w_ready; // @[SpectrometerTestWithoutLA.scala 73:29]
  wire  nco_mux_0_auto_register_in_w_valid; // @[SpectrometerTestWithoutLA.scala 73:29]
  wire [31:0] nco_mux_0_auto_register_in_w_bits_data; // @[SpectrometerTestWithoutLA.scala 73:29]
  wire [3:0] nco_mux_0_auto_register_in_w_bits_strb; // @[SpectrometerTestWithoutLA.scala 73:29]
  wire  nco_mux_0_auto_register_in_b_ready; // @[SpectrometerTestWithoutLA.scala 73:29]
  wire  nco_mux_0_auto_register_in_b_valid; // @[SpectrometerTestWithoutLA.scala 73:29]
  wire  nco_mux_0_auto_register_in_b_bits_id; // @[SpectrometerTestWithoutLA.scala 73:29]
  wire  nco_mux_0_auto_register_in_ar_ready; // @[SpectrometerTestWithoutLA.scala 73:29]
  wire  nco_mux_0_auto_register_in_ar_valid; // @[SpectrometerTestWithoutLA.scala 73:29]
  wire  nco_mux_0_auto_register_in_ar_bits_id; // @[SpectrometerTestWithoutLA.scala 73:29]
  wire [29:0] nco_mux_0_auto_register_in_ar_bits_addr; // @[SpectrometerTestWithoutLA.scala 73:29]
  wire [2:0] nco_mux_0_auto_register_in_ar_bits_size; // @[SpectrometerTestWithoutLA.scala 73:29]
  wire  nco_mux_0_auto_register_in_r_ready; // @[SpectrometerTestWithoutLA.scala 73:29]
  wire  nco_mux_0_auto_register_in_r_valid; // @[SpectrometerTestWithoutLA.scala 73:29]
  wire  nco_mux_0_auto_register_in_r_bits_id; // @[SpectrometerTestWithoutLA.scala 73:29]
  wire [31:0] nco_mux_0_auto_register_in_r_bits_data; // @[SpectrometerTestWithoutLA.scala 73:29]
  wire  nco_mux_0_auto_stream_in_2_ready; // @[SpectrometerTestWithoutLA.scala 73:29]
  wire  nco_mux_0_auto_stream_in_2_valid; // @[SpectrometerTestWithoutLA.scala 73:29]
  wire [31:0] nco_mux_0_auto_stream_in_2_bits_data; // @[SpectrometerTestWithoutLA.scala 73:29]
  wire  nco_mux_0_auto_stream_in_2_bits_last; // @[SpectrometerTestWithoutLA.scala 73:29]
  wire  nco_mux_0_auto_stream_in_1_ready; // @[SpectrometerTestWithoutLA.scala 73:29]
  wire  nco_mux_0_auto_stream_in_1_valid; // @[SpectrometerTestWithoutLA.scala 73:29]
  wire [31:0] nco_mux_0_auto_stream_in_1_bits_data; // @[SpectrometerTestWithoutLA.scala 73:29]
  wire  nco_mux_0_auto_stream_in_1_bits_last; // @[SpectrometerTestWithoutLA.scala 73:29]
  wire  nco_mux_0_auto_stream_in_0_ready; // @[SpectrometerTestWithoutLA.scala 73:29]
  wire  nco_mux_0_auto_stream_in_0_valid; // @[SpectrometerTestWithoutLA.scala 73:29]
  wire [31:0] nco_mux_0_auto_stream_in_0_bits_data; // @[SpectrometerTestWithoutLA.scala 73:29]
  wire  nco_mux_0_auto_stream_in_0_bits_last; // @[SpectrometerTestWithoutLA.scala 73:29]
  wire  nco_mux_0_auto_stream_out_0_ready; // @[SpectrometerTestWithoutLA.scala 73:29]
  wire  nco_mux_0_auto_stream_out_0_valid; // @[SpectrometerTestWithoutLA.scala 73:29]
  wire [31:0] nco_mux_0_auto_stream_out_0_bits_data; // @[SpectrometerTestWithoutLA.scala 73:29]
  wire  nco_mux_0_auto_stream_out_0_bits_last; // @[SpectrometerTestWithoutLA.scala 73:29]
  wire  nco_mux_1_clock; // @[SpectrometerTestWithoutLA.scala 74:29]
  wire  nco_mux_1_reset; // @[SpectrometerTestWithoutLA.scala 74:29]
  wire  nco_mux_1_auto_register_in_aw_ready; // @[SpectrometerTestWithoutLA.scala 74:29]
  wire  nco_mux_1_auto_register_in_aw_valid; // @[SpectrometerTestWithoutLA.scala 74:29]
  wire  nco_mux_1_auto_register_in_aw_bits_id; // @[SpectrometerTestWithoutLA.scala 74:29]
  wire [29:0] nco_mux_1_auto_register_in_aw_bits_addr; // @[SpectrometerTestWithoutLA.scala 74:29]
  wire  nco_mux_1_auto_register_in_w_ready; // @[SpectrometerTestWithoutLA.scala 74:29]
  wire  nco_mux_1_auto_register_in_w_valid; // @[SpectrometerTestWithoutLA.scala 74:29]
  wire [31:0] nco_mux_1_auto_register_in_w_bits_data; // @[SpectrometerTestWithoutLA.scala 74:29]
  wire [3:0] nco_mux_1_auto_register_in_w_bits_strb; // @[SpectrometerTestWithoutLA.scala 74:29]
  wire  nco_mux_1_auto_register_in_b_ready; // @[SpectrometerTestWithoutLA.scala 74:29]
  wire  nco_mux_1_auto_register_in_b_valid; // @[SpectrometerTestWithoutLA.scala 74:29]
  wire  nco_mux_1_auto_register_in_b_bits_id; // @[SpectrometerTestWithoutLA.scala 74:29]
  wire  nco_mux_1_auto_register_in_ar_ready; // @[SpectrometerTestWithoutLA.scala 74:29]
  wire  nco_mux_1_auto_register_in_ar_valid; // @[SpectrometerTestWithoutLA.scala 74:29]
  wire  nco_mux_1_auto_register_in_ar_bits_id; // @[SpectrometerTestWithoutLA.scala 74:29]
  wire [29:0] nco_mux_1_auto_register_in_ar_bits_addr; // @[SpectrometerTestWithoutLA.scala 74:29]
  wire [2:0] nco_mux_1_auto_register_in_ar_bits_size; // @[SpectrometerTestWithoutLA.scala 74:29]
  wire  nco_mux_1_auto_register_in_r_ready; // @[SpectrometerTestWithoutLA.scala 74:29]
  wire  nco_mux_1_auto_register_in_r_valid; // @[SpectrometerTestWithoutLA.scala 74:29]
  wire  nco_mux_1_auto_register_in_r_bits_id; // @[SpectrometerTestWithoutLA.scala 74:29]
  wire [31:0] nco_mux_1_auto_register_in_r_bits_data; // @[SpectrometerTestWithoutLA.scala 74:29]
  wire  nco_mux_1_auto_stream_in_ready; // @[SpectrometerTestWithoutLA.scala 74:29]
  wire  nco_mux_1_auto_stream_in_valid; // @[SpectrometerTestWithoutLA.scala 74:29]
  wire [31:0] nco_mux_1_auto_stream_in_bits_data; // @[SpectrometerTestWithoutLA.scala 74:29]
  wire  nco_mux_1_auto_stream_in_bits_last; // @[SpectrometerTestWithoutLA.scala 74:29]
  wire  nco_mux_1_auto_stream_out_1_ready; // @[SpectrometerTestWithoutLA.scala 74:29]
  wire  nco_mux_1_auto_stream_out_1_valid; // @[SpectrometerTestWithoutLA.scala 74:29]
  wire [31:0] nco_mux_1_auto_stream_out_1_bits_data; // @[SpectrometerTestWithoutLA.scala 74:29]
  wire  nco_mux_1_auto_stream_out_1_bits_last; // @[SpectrometerTestWithoutLA.scala 74:29]
  wire  fft_clock; // @[SpectrometerTestWithoutLA.scala 80:29]
  wire  fft_reset; // @[SpectrometerTestWithoutLA.scala 80:29]
  wire  fft_auto_mem_in_aw_ready; // @[SpectrometerTestWithoutLA.scala 80:29]
  wire  fft_auto_mem_in_aw_valid; // @[SpectrometerTestWithoutLA.scala 80:29]
  wire  fft_auto_mem_in_aw_bits_id; // @[SpectrometerTestWithoutLA.scala 80:29]
  wire [29:0] fft_auto_mem_in_aw_bits_addr; // @[SpectrometerTestWithoutLA.scala 80:29]
  wire  fft_auto_mem_in_w_ready; // @[SpectrometerTestWithoutLA.scala 80:29]
  wire  fft_auto_mem_in_w_valid; // @[SpectrometerTestWithoutLA.scala 80:29]
  wire [31:0] fft_auto_mem_in_w_bits_data; // @[SpectrometerTestWithoutLA.scala 80:29]
  wire [3:0] fft_auto_mem_in_w_bits_strb; // @[SpectrometerTestWithoutLA.scala 80:29]
  wire  fft_auto_mem_in_b_ready; // @[SpectrometerTestWithoutLA.scala 80:29]
  wire  fft_auto_mem_in_b_valid; // @[SpectrometerTestWithoutLA.scala 80:29]
  wire  fft_auto_mem_in_b_bits_id; // @[SpectrometerTestWithoutLA.scala 80:29]
  wire  fft_auto_mem_in_ar_ready; // @[SpectrometerTestWithoutLA.scala 80:29]
  wire  fft_auto_mem_in_ar_valid; // @[SpectrometerTestWithoutLA.scala 80:29]
  wire  fft_auto_mem_in_ar_bits_id; // @[SpectrometerTestWithoutLA.scala 80:29]
  wire [29:0] fft_auto_mem_in_ar_bits_addr; // @[SpectrometerTestWithoutLA.scala 80:29]
  wire [2:0] fft_auto_mem_in_ar_bits_size; // @[SpectrometerTestWithoutLA.scala 80:29]
  wire  fft_auto_mem_in_r_ready; // @[SpectrometerTestWithoutLA.scala 80:29]
  wire  fft_auto_mem_in_r_valid; // @[SpectrometerTestWithoutLA.scala 80:29]
  wire  fft_auto_mem_in_r_bits_id; // @[SpectrometerTestWithoutLA.scala 80:29]
  wire [31:0] fft_auto_mem_in_r_bits_data; // @[SpectrometerTestWithoutLA.scala 80:29]
  wire  fft_auto_stream_in_ready; // @[SpectrometerTestWithoutLA.scala 80:29]
  wire  fft_auto_stream_in_valid; // @[SpectrometerTestWithoutLA.scala 80:29]
  wire [31:0] fft_auto_stream_in_bits_data; // @[SpectrometerTestWithoutLA.scala 80:29]
  wire  fft_auto_stream_in_bits_last; // @[SpectrometerTestWithoutLA.scala 80:29]
  wire  fft_auto_stream_out_ready; // @[SpectrometerTestWithoutLA.scala 80:29]
  wire  fft_auto_stream_out_valid; // @[SpectrometerTestWithoutLA.scala 80:29]
  wire [31:0] fft_auto_stream_out_bits_data; // @[SpectrometerTestWithoutLA.scala 80:29]
  wire  fft_auto_stream_out_bits_last; // @[SpectrometerTestWithoutLA.scala 80:29]
  wire  fft_split_clock; // @[SpectrometerTestWithoutLA.scala 81:29]
  wire  fft_split_reset; // @[SpectrometerTestWithoutLA.scala 81:29]
  wire  fft_split_auto_mem_in_aw_ready; // @[SpectrometerTestWithoutLA.scala 81:29]
  wire  fft_split_auto_mem_in_aw_valid; // @[SpectrometerTestWithoutLA.scala 81:29]
  wire  fft_split_auto_mem_in_aw_bits_id; // @[SpectrometerTestWithoutLA.scala 81:29]
  wire [29:0] fft_split_auto_mem_in_aw_bits_addr; // @[SpectrometerTestWithoutLA.scala 81:29]
  wire  fft_split_auto_mem_in_w_ready; // @[SpectrometerTestWithoutLA.scala 81:29]
  wire  fft_split_auto_mem_in_w_valid; // @[SpectrometerTestWithoutLA.scala 81:29]
  wire [31:0] fft_split_auto_mem_in_w_bits_data; // @[SpectrometerTestWithoutLA.scala 81:29]
  wire [3:0] fft_split_auto_mem_in_w_bits_strb; // @[SpectrometerTestWithoutLA.scala 81:29]
  wire  fft_split_auto_mem_in_b_ready; // @[SpectrometerTestWithoutLA.scala 81:29]
  wire  fft_split_auto_mem_in_b_valid; // @[SpectrometerTestWithoutLA.scala 81:29]
  wire  fft_split_auto_mem_in_b_bits_id; // @[SpectrometerTestWithoutLA.scala 81:29]
  wire  fft_split_auto_mem_in_ar_ready; // @[SpectrometerTestWithoutLA.scala 81:29]
  wire  fft_split_auto_mem_in_ar_valid; // @[SpectrometerTestWithoutLA.scala 81:29]
  wire  fft_split_auto_mem_in_ar_bits_id; // @[SpectrometerTestWithoutLA.scala 81:29]
  wire [29:0] fft_split_auto_mem_in_ar_bits_addr; // @[SpectrometerTestWithoutLA.scala 81:29]
  wire [2:0] fft_split_auto_mem_in_ar_bits_size; // @[SpectrometerTestWithoutLA.scala 81:29]
  wire  fft_split_auto_mem_in_r_ready; // @[SpectrometerTestWithoutLA.scala 81:29]
  wire  fft_split_auto_mem_in_r_valid; // @[SpectrometerTestWithoutLA.scala 81:29]
  wire  fft_split_auto_mem_in_r_bits_id; // @[SpectrometerTestWithoutLA.scala 81:29]
  wire [31:0] fft_split_auto_mem_in_r_bits_data; // @[SpectrometerTestWithoutLA.scala 81:29]
  wire  fft_split_auto_stream_in_ready; // @[SpectrometerTestWithoutLA.scala 81:29]
  wire  fft_split_auto_stream_in_valid; // @[SpectrometerTestWithoutLA.scala 81:29]
  wire [31:0] fft_split_auto_stream_in_bits_data; // @[SpectrometerTestWithoutLA.scala 81:29]
  wire  fft_split_auto_stream_in_bits_last; // @[SpectrometerTestWithoutLA.scala 81:29]
  wire  fft_split_auto_stream_out_1_ready; // @[SpectrometerTestWithoutLA.scala 81:29]
  wire  fft_split_auto_stream_out_1_valid; // @[SpectrometerTestWithoutLA.scala 81:29]
  wire [31:0] fft_split_auto_stream_out_1_bits_data; // @[SpectrometerTestWithoutLA.scala 81:29]
  wire  fft_split_auto_stream_out_1_bits_last; // @[SpectrometerTestWithoutLA.scala 81:29]
  wire  fft_split_auto_stream_out_0_ready; // @[SpectrometerTestWithoutLA.scala 81:29]
  wire  fft_split_auto_stream_out_0_valid; // @[SpectrometerTestWithoutLA.scala 81:29]
  wire [31:0] fft_split_auto_stream_out_0_bits_data; // @[SpectrometerTestWithoutLA.scala 81:29]
  wire  fft_split_auto_stream_out_0_bits_last; // @[SpectrometerTestWithoutLA.scala 81:29]
  wire  fft_mux_0_clock; // @[SpectrometerTestWithoutLA.scala 82:29]
  wire  fft_mux_0_reset; // @[SpectrometerTestWithoutLA.scala 82:29]
  wire  fft_mux_0_auto_register_in_aw_ready; // @[SpectrometerTestWithoutLA.scala 82:29]
  wire  fft_mux_0_auto_register_in_aw_valid; // @[SpectrometerTestWithoutLA.scala 82:29]
  wire  fft_mux_0_auto_register_in_aw_bits_id; // @[SpectrometerTestWithoutLA.scala 82:29]
  wire [29:0] fft_mux_0_auto_register_in_aw_bits_addr; // @[SpectrometerTestWithoutLA.scala 82:29]
  wire  fft_mux_0_auto_register_in_w_ready; // @[SpectrometerTestWithoutLA.scala 82:29]
  wire  fft_mux_0_auto_register_in_w_valid; // @[SpectrometerTestWithoutLA.scala 82:29]
  wire [31:0] fft_mux_0_auto_register_in_w_bits_data; // @[SpectrometerTestWithoutLA.scala 82:29]
  wire [3:0] fft_mux_0_auto_register_in_w_bits_strb; // @[SpectrometerTestWithoutLA.scala 82:29]
  wire  fft_mux_0_auto_register_in_b_ready; // @[SpectrometerTestWithoutLA.scala 82:29]
  wire  fft_mux_0_auto_register_in_b_valid; // @[SpectrometerTestWithoutLA.scala 82:29]
  wire  fft_mux_0_auto_register_in_b_bits_id; // @[SpectrometerTestWithoutLA.scala 82:29]
  wire  fft_mux_0_auto_register_in_ar_ready; // @[SpectrometerTestWithoutLA.scala 82:29]
  wire  fft_mux_0_auto_register_in_ar_valid; // @[SpectrometerTestWithoutLA.scala 82:29]
  wire  fft_mux_0_auto_register_in_ar_bits_id; // @[SpectrometerTestWithoutLA.scala 82:29]
  wire [29:0] fft_mux_0_auto_register_in_ar_bits_addr; // @[SpectrometerTestWithoutLA.scala 82:29]
  wire [2:0] fft_mux_0_auto_register_in_ar_bits_size; // @[SpectrometerTestWithoutLA.scala 82:29]
  wire  fft_mux_0_auto_register_in_r_ready; // @[SpectrometerTestWithoutLA.scala 82:29]
  wire  fft_mux_0_auto_register_in_r_valid; // @[SpectrometerTestWithoutLA.scala 82:29]
  wire  fft_mux_0_auto_register_in_r_bits_id; // @[SpectrometerTestWithoutLA.scala 82:29]
  wire [31:0] fft_mux_0_auto_register_in_r_bits_data; // @[SpectrometerTestWithoutLA.scala 82:29]
  wire  fft_mux_0_auto_stream_in_2_ready; // @[SpectrometerTestWithoutLA.scala 82:29]
  wire  fft_mux_0_auto_stream_in_2_valid; // @[SpectrometerTestWithoutLA.scala 82:29]
  wire [31:0] fft_mux_0_auto_stream_in_2_bits_data; // @[SpectrometerTestWithoutLA.scala 82:29]
  wire  fft_mux_0_auto_stream_in_2_bits_last; // @[SpectrometerTestWithoutLA.scala 82:29]
  wire  fft_mux_0_auto_stream_in_1_ready; // @[SpectrometerTestWithoutLA.scala 82:29]
  wire  fft_mux_0_auto_stream_in_1_valid; // @[SpectrometerTestWithoutLA.scala 82:29]
  wire [31:0] fft_mux_0_auto_stream_in_1_bits_data; // @[SpectrometerTestWithoutLA.scala 82:29]
  wire  fft_mux_0_auto_stream_in_1_bits_last; // @[SpectrometerTestWithoutLA.scala 82:29]
  wire  fft_mux_0_auto_stream_in_0_ready; // @[SpectrometerTestWithoutLA.scala 82:29]
  wire  fft_mux_0_auto_stream_in_0_valid; // @[SpectrometerTestWithoutLA.scala 82:29]
  wire [31:0] fft_mux_0_auto_stream_in_0_bits_data; // @[SpectrometerTestWithoutLA.scala 82:29]
  wire  fft_mux_0_auto_stream_in_0_bits_last; // @[SpectrometerTestWithoutLA.scala 82:29]
  wire  fft_mux_0_auto_stream_out_0_ready; // @[SpectrometerTestWithoutLA.scala 82:29]
  wire  fft_mux_0_auto_stream_out_0_valid; // @[SpectrometerTestWithoutLA.scala 82:29]
  wire [31:0] fft_mux_0_auto_stream_out_0_bits_data; // @[SpectrometerTestWithoutLA.scala 82:29]
  wire  fft_mux_0_auto_stream_out_0_bits_last; // @[SpectrometerTestWithoutLA.scala 82:29]
  wire  fft_mux_1_clock; // @[SpectrometerTestWithoutLA.scala 83:29]
  wire  fft_mux_1_reset; // @[SpectrometerTestWithoutLA.scala 83:29]
  wire  fft_mux_1_auto_register_in_aw_ready; // @[SpectrometerTestWithoutLA.scala 83:29]
  wire  fft_mux_1_auto_register_in_aw_valid; // @[SpectrometerTestWithoutLA.scala 83:29]
  wire  fft_mux_1_auto_register_in_aw_bits_id; // @[SpectrometerTestWithoutLA.scala 83:29]
  wire [29:0] fft_mux_1_auto_register_in_aw_bits_addr; // @[SpectrometerTestWithoutLA.scala 83:29]
  wire  fft_mux_1_auto_register_in_w_ready; // @[SpectrometerTestWithoutLA.scala 83:29]
  wire  fft_mux_1_auto_register_in_w_valid; // @[SpectrometerTestWithoutLA.scala 83:29]
  wire [31:0] fft_mux_1_auto_register_in_w_bits_data; // @[SpectrometerTestWithoutLA.scala 83:29]
  wire [3:0] fft_mux_1_auto_register_in_w_bits_strb; // @[SpectrometerTestWithoutLA.scala 83:29]
  wire  fft_mux_1_auto_register_in_b_ready; // @[SpectrometerTestWithoutLA.scala 83:29]
  wire  fft_mux_1_auto_register_in_b_valid; // @[SpectrometerTestWithoutLA.scala 83:29]
  wire  fft_mux_1_auto_register_in_b_bits_id; // @[SpectrometerTestWithoutLA.scala 83:29]
  wire  fft_mux_1_auto_register_in_ar_ready; // @[SpectrometerTestWithoutLA.scala 83:29]
  wire  fft_mux_1_auto_register_in_ar_valid; // @[SpectrometerTestWithoutLA.scala 83:29]
  wire  fft_mux_1_auto_register_in_ar_bits_id; // @[SpectrometerTestWithoutLA.scala 83:29]
  wire [29:0] fft_mux_1_auto_register_in_ar_bits_addr; // @[SpectrometerTestWithoutLA.scala 83:29]
  wire [2:0] fft_mux_1_auto_register_in_ar_bits_size; // @[SpectrometerTestWithoutLA.scala 83:29]
  wire  fft_mux_1_auto_register_in_r_ready; // @[SpectrometerTestWithoutLA.scala 83:29]
  wire  fft_mux_1_auto_register_in_r_valid; // @[SpectrometerTestWithoutLA.scala 83:29]
  wire  fft_mux_1_auto_register_in_r_bits_id; // @[SpectrometerTestWithoutLA.scala 83:29]
  wire [31:0] fft_mux_1_auto_register_in_r_bits_data; // @[SpectrometerTestWithoutLA.scala 83:29]
  wire  fft_mux_1_auto_stream_in_ready; // @[SpectrometerTestWithoutLA.scala 83:29]
  wire  fft_mux_1_auto_stream_in_valid; // @[SpectrometerTestWithoutLA.scala 83:29]
  wire [31:0] fft_mux_1_auto_stream_in_bits_data; // @[SpectrometerTestWithoutLA.scala 83:29]
  wire  fft_mux_1_auto_stream_in_bits_last; // @[SpectrometerTestWithoutLA.scala 83:29]
  wire  fft_mux_1_auto_stream_out_1_ready; // @[SpectrometerTestWithoutLA.scala 83:29]
  wire  fft_mux_1_auto_stream_out_1_valid; // @[SpectrometerTestWithoutLA.scala 83:29]
  wire [31:0] fft_mux_1_auto_stream_out_1_bits_data; // @[SpectrometerTestWithoutLA.scala 83:29]
  wire  fft_mux_1_auto_stream_out_1_bits_last; // @[SpectrometerTestWithoutLA.scala 83:29]
  wire  mag_clock; // @[SpectrometerTestWithoutLA.scala 89:29]
  wire  mag_reset; // @[SpectrometerTestWithoutLA.scala 89:29]
  wire  mag_auto_mem_in_aw_ready; // @[SpectrometerTestWithoutLA.scala 89:29]
  wire  mag_auto_mem_in_aw_valid; // @[SpectrometerTestWithoutLA.scala 89:29]
  wire  mag_auto_mem_in_aw_bits_id; // @[SpectrometerTestWithoutLA.scala 89:29]
  wire [29:0] mag_auto_mem_in_aw_bits_addr; // @[SpectrometerTestWithoutLA.scala 89:29]
  wire  mag_auto_mem_in_w_ready; // @[SpectrometerTestWithoutLA.scala 89:29]
  wire  mag_auto_mem_in_w_valid; // @[SpectrometerTestWithoutLA.scala 89:29]
  wire [31:0] mag_auto_mem_in_w_bits_data; // @[SpectrometerTestWithoutLA.scala 89:29]
  wire [3:0] mag_auto_mem_in_w_bits_strb; // @[SpectrometerTestWithoutLA.scala 89:29]
  wire  mag_auto_mem_in_b_ready; // @[SpectrometerTestWithoutLA.scala 89:29]
  wire  mag_auto_mem_in_b_valid; // @[SpectrometerTestWithoutLA.scala 89:29]
  wire  mag_auto_mem_in_b_bits_id; // @[SpectrometerTestWithoutLA.scala 89:29]
  wire  mag_auto_mem_in_ar_ready; // @[SpectrometerTestWithoutLA.scala 89:29]
  wire  mag_auto_mem_in_ar_valid; // @[SpectrometerTestWithoutLA.scala 89:29]
  wire  mag_auto_mem_in_ar_bits_id; // @[SpectrometerTestWithoutLA.scala 89:29]
  wire [29:0] mag_auto_mem_in_ar_bits_addr; // @[SpectrometerTestWithoutLA.scala 89:29]
  wire [2:0] mag_auto_mem_in_ar_bits_size; // @[SpectrometerTestWithoutLA.scala 89:29]
  wire  mag_auto_mem_in_r_ready; // @[SpectrometerTestWithoutLA.scala 89:29]
  wire  mag_auto_mem_in_r_valid; // @[SpectrometerTestWithoutLA.scala 89:29]
  wire  mag_auto_mem_in_r_bits_id; // @[SpectrometerTestWithoutLA.scala 89:29]
  wire [31:0] mag_auto_mem_in_r_bits_data; // @[SpectrometerTestWithoutLA.scala 89:29]
  wire  mag_auto_stream_in_ready; // @[SpectrometerTestWithoutLA.scala 89:29]
  wire  mag_auto_stream_in_valid; // @[SpectrometerTestWithoutLA.scala 89:29]
  wire [31:0] mag_auto_stream_in_bits_data; // @[SpectrometerTestWithoutLA.scala 89:29]
  wire  mag_auto_stream_in_bits_last; // @[SpectrometerTestWithoutLA.scala 89:29]
  wire  mag_auto_stream_out_ready; // @[SpectrometerTestWithoutLA.scala 89:29]
  wire  mag_auto_stream_out_valid; // @[SpectrometerTestWithoutLA.scala 89:29]
  wire [31:0] mag_auto_stream_out_bits_data; // @[SpectrometerTestWithoutLA.scala 89:29]
  wire  mag_auto_stream_out_bits_last; // @[SpectrometerTestWithoutLA.scala 89:29]
  wire  mag_split_clock; // @[SpectrometerTestWithoutLA.scala 90:29]
  wire  mag_split_reset; // @[SpectrometerTestWithoutLA.scala 90:29]
  wire  mag_split_auto_mem_in_aw_ready; // @[SpectrometerTestWithoutLA.scala 90:29]
  wire  mag_split_auto_mem_in_aw_valid; // @[SpectrometerTestWithoutLA.scala 90:29]
  wire  mag_split_auto_mem_in_aw_bits_id; // @[SpectrometerTestWithoutLA.scala 90:29]
  wire [29:0] mag_split_auto_mem_in_aw_bits_addr; // @[SpectrometerTestWithoutLA.scala 90:29]
  wire  mag_split_auto_mem_in_w_ready; // @[SpectrometerTestWithoutLA.scala 90:29]
  wire  mag_split_auto_mem_in_w_valid; // @[SpectrometerTestWithoutLA.scala 90:29]
  wire [31:0] mag_split_auto_mem_in_w_bits_data; // @[SpectrometerTestWithoutLA.scala 90:29]
  wire [3:0] mag_split_auto_mem_in_w_bits_strb; // @[SpectrometerTestWithoutLA.scala 90:29]
  wire  mag_split_auto_mem_in_b_ready; // @[SpectrometerTestWithoutLA.scala 90:29]
  wire  mag_split_auto_mem_in_b_valid; // @[SpectrometerTestWithoutLA.scala 90:29]
  wire  mag_split_auto_mem_in_b_bits_id; // @[SpectrometerTestWithoutLA.scala 90:29]
  wire  mag_split_auto_mem_in_ar_ready; // @[SpectrometerTestWithoutLA.scala 90:29]
  wire  mag_split_auto_mem_in_ar_valid; // @[SpectrometerTestWithoutLA.scala 90:29]
  wire  mag_split_auto_mem_in_ar_bits_id; // @[SpectrometerTestWithoutLA.scala 90:29]
  wire [29:0] mag_split_auto_mem_in_ar_bits_addr; // @[SpectrometerTestWithoutLA.scala 90:29]
  wire [2:0] mag_split_auto_mem_in_ar_bits_size; // @[SpectrometerTestWithoutLA.scala 90:29]
  wire  mag_split_auto_mem_in_r_ready; // @[SpectrometerTestWithoutLA.scala 90:29]
  wire  mag_split_auto_mem_in_r_valid; // @[SpectrometerTestWithoutLA.scala 90:29]
  wire  mag_split_auto_mem_in_r_bits_id; // @[SpectrometerTestWithoutLA.scala 90:29]
  wire [31:0] mag_split_auto_mem_in_r_bits_data; // @[SpectrometerTestWithoutLA.scala 90:29]
  wire  mag_split_auto_stream_in_ready; // @[SpectrometerTestWithoutLA.scala 90:29]
  wire  mag_split_auto_stream_in_valid; // @[SpectrometerTestWithoutLA.scala 90:29]
  wire [31:0] mag_split_auto_stream_in_bits_data; // @[SpectrometerTestWithoutLA.scala 90:29]
  wire  mag_split_auto_stream_in_bits_last; // @[SpectrometerTestWithoutLA.scala 90:29]
  wire  mag_split_auto_stream_out_1_ready; // @[SpectrometerTestWithoutLA.scala 90:29]
  wire  mag_split_auto_stream_out_1_valid; // @[SpectrometerTestWithoutLA.scala 90:29]
  wire [31:0] mag_split_auto_stream_out_1_bits_data; // @[SpectrometerTestWithoutLA.scala 90:29]
  wire  mag_split_auto_stream_out_1_bits_last; // @[SpectrometerTestWithoutLA.scala 90:29]
  wire  mag_split_auto_stream_out_0_ready; // @[SpectrometerTestWithoutLA.scala 90:29]
  wire  mag_split_auto_stream_out_0_valid; // @[SpectrometerTestWithoutLA.scala 90:29]
  wire [31:0] mag_split_auto_stream_out_0_bits_data; // @[SpectrometerTestWithoutLA.scala 90:29]
  wire  mag_split_auto_stream_out_0_bits_last; // @[SpectrometerTestWithoutLA.scala 90:29]
  wire  mag_mux_0_clock; // @[SpectrometerTestWithoutLA.scala 91:29]
  wire  mag_mux_0_reset; // @[SpectrometerTestWithoutLA.scala 91:29]
  wire  mag_mux_0_auto_register_in_aw_ready; // @[SpectrometerTestWithoutLA.scala 91:29]
  wire  mag_mux_0_auto_register_in_aw_valid; // @[SpectrometerTestWithoutLA.scala 91:29]
  wire  mag_mux_0_auto_register_in_aw_bits_id; // @[SpectrometerTestWithoutLA.scala 91:29]
  wire [29:0] mag_mux_0_auto_register_in_aw_bits_addr; // @[SpectrometerTestWithoutLA.scala 91:29]
  wire  mag_mux_0_auto_register_in_w_ready; // @[SpectrometerTestWithoutLA.scala 91:29]
  wire  mag_mux_0_auto_register_in_w_valid; // @[SpectrometerTestWithoutLA.scala 91:29]
  wire [31:0] mag_mux_0_auto_register_in_w_bits_data; // @[SpectrometerTestWithoutLA.scala 91:29]
  wire [3:0] mag_mux_0_auto_register_in_w_bits_strb; // @[SpectrometerTestWithoutLA.scala 91:29]
  wire  mag_mux_0_auto_register_in_b_ready; // @[SpectrometerTestWithoutLA.scala 91:29]
  wire  mag_mux_0_auto_register_in_b_valid; // @[SpectrometerTestWithoutLA.scala 91:29]
  wire  mag_mux_0_auto_register_in_b_bits_id; // @[SpectrometerTestWithoutLA.scala 91:29]
  wire  mag_mux_0_auto_register_in_ar_ready; // @[SpectrometerTestWithoutLA.scala 91:29]
  wire  mag_mux_0_auto_register_in_ar_valid; // @[SpectrometerTestWithoutLA.scala 91:29]
  wire  mag_mux_0_auto_register_in_ar_bits_id; // @[SpectrometerTestWithoutLA.scala 91:29]
  wire [29:0] mag_mux_0_auto_register_in_ar_bits_addr; // @[SpectrometerTestWithoutLA.scala 91:29]
  wire [2:0] mag_mux_0_auto_register_in_ar_bits_size; // @[SpectrometerTestWithoutLA.scala 91:29]
  wire  mag_mux_0_auto_register_in_r_ready; // @[SpectrometerTestWithoutLA.scala 91:29]
  wire  mag_mux_0_auto_register_in_r_valid; // @[SpectrometerTestWithoutLA.scala 91:29]
  wire  mag_mux_0_auto_register_in_r_bits_id; // @[SpectrometerTestWithoutLA.scala 91:29]
  wire [31:0] mag_mux_0_auto_register_in_r_bits_data; // @[SpectrometerTestWithoutLA.scala 91:29]
  wire  mag_mux_0_auto_stream_in_2_ready; // @[SpectrometerTestWithoutLA.scala 91:29]
  wire  mag_mux_0_auto_stream_in_2_valid; // @[SpectrometerTestWithoutLA.scala 91:29]
  wire [31:0] mag_mux_0_auto_stream_in_2_bits_data; // @[SpectrometerTestWithoutLA.scala 91:29]
  wire  mag_mux_0_auto_stream_in_2_bits_last; // @[SpectrometerTestWithoutLA.scala 91:29]
  wire  mag_mux_0_auto_stream_in_1_ready; // @[SpectrometerTestWithoutLA.scala 91:29]
  wire  mag_mux_0_auto_stream_in_1_valid; // @[SpectrometerTestWithoutLA.scala 91:29]
  wire [31:0] mag_mux_0_auto_stream_in_1_bits_data; // @[SpectrometerTestWithoutLA.scala 91:29]
  wire  mag_mux_0_auto_stream_in_1_bits_last; // @[SpectrometerTestWithoutLA.scala 91:29]
  wire  mag_mux_0_auto_stream_in_0_ready; // @[SpectrometerTestWithoutLA.scala 91:29]
  wire  mag_mux_0_auto_stream_in_0_valid; // @[SpectrometerTestWithoutLA.scala 91:29]
  wire [31:0] mag_mux_0_auto_stream_in_0_bits_data; // @[SpectrometerTestWithoutLA.scala 91:29]
  wire  mag_mux_0_auto_stream_in_0_bits_last; // @[SpectrometerTestWithoutLA.scala 91:29]
  wire  mag_mux_0_auto_stream_out_0_ready; // @[SpectrometerTestWithoutLA.scala 91:29]
  wire  mag_mux_0_auto_stream_out_0_valid; // @[SpectrometerTestWithoutLA.scala 91:29]
  wire [31:0] mag_mux_0_auto_stream_out_0_bits_data; // @[SpectrometerTestWithoutLA.scala 91:29]
  wire  mag_mux_0_auto_stream_out_0_bits_last; // @[SpectrometerTestWithoutLA.scala 91:29]
  wire  mag_mux_1_clock; // @[SpectrometerTestWithoutLA.scala 92:29]
  wire  mag_mux_1_reset; // @[SpectrometerTestWithoutLA.scala 92:29]
  wire  mag_mux_1_auto_register_in_aw_ready; // @[SpectrometerTestWithoutLA.scala 92:29]
  wire  mag_mux_1_auto_register_in_aw_valid; // @[SpectrometerTestWithoutLA.scala 92:29]
  wire  mag_mux_1_auto_register_in_aw_bits_id; // @[SpectrometerTestWithoutLA.scala 92:29]
  wire [29:0] mag_mux_1_auto_register_in_aw_bits_addr; // @[SpectrometerTestWithoutLA.scala 92:29]
  wire  mag_mux_1_auto_register_in_w_ready; // @[SpectrometerTestWithoutLA.scala 92:29]
  wire  mag_mux_1_auto_register_in_w_valid; // @[SpectrometerTestWithoutLA.scala 92:29]
  wire [31:0] mag_mux_1_auto_register_in_w_bits_data; // @[SpectrometerTestWithoutLA.scala 92:29]
  wire [3:0] mag_mux_1_auto_register_in_w_bits_strb; // @[SpectrometerTestWithoutLA.scala 92:29]
  wire  mag_mux_1_auto_register_in_b_ready; // @[SpectrometerTestWithoutLA.scala 92:29]
  wire  mag_mux_1_auto_register_in_b_valid; // @[SpectrometerTestWithoutLA.scala 92:29]
  wire  mag_mux_1_auto_register_in_b_bits_id; // @[SpectrometerTestWithoutLA.scala 92:29]
  wire  mag_mux_1_auto_register_in_ar_ready; // @[SpectrometerTestWithoutLA.scala 92:29]
  wire  mag_mux_1_auto_register_in_ar_valid; // @[SpectrometerTestWithoutLA.scala 92:29]
  wire  mag_mux_1_auto_register_in_ar_bits_id; // @[SpectrometerTestWithoutLA.scala 92:29]
  wire [29:0] mag_mux_1_auto_register_in_ar_bits_addr; // @[SpectrometerTestWithoutLA.scala 92:29]
  wire [2:0] mag_mux_1_auto_register_in_ar_bits_size; // @[SpectrometerTestWithoutLA.scala 92:29]
  wire  mag_mux_1_auto_register_in_r_ready; // @[SpectrometerTestWithoutLA.scala 92:29]
  wire  mag_mux_1_auto_register_in_r_valid; // @[SpectrometerTestWithoutLA.scala 92:29]
  wire  mag_mux_1_auto_register_in_r_bits_id; // @[SpectrometerTestWithoutLA.scala 92:29]
  wire [31:0] mag_mux_1_auto_register_in_r_bits_data; // @[SpectrometerTestWithoutLA.scala 92:29]
  wire  mag_mux_1_auto_stream_in_ready; // @[SpectrometerTestWithoutLA.scala 92:29]
  wire  mag_mux_1_auto_stream_in_valid; // @[SpectrometerTestWithoutLA.scala 92:29]
  wire [31:0] mag_mux_1_auto_stream_in_bits_data; // @[SpectrometerTestWithoutLA.scala 92:29]
  wire  mag_mux_1_auto_stream_in_bits_last; // @[SpectrometerTestWithoutLA.scala 92:29]
  wire  mag_mux_1_auto_stream_out_1_ready; // @[SpectrometerTestWithoutLA.scala 92:29]
  wire  mag_mux_1_auto_stream_out_1_valid; // @[SpectrometerTestWithoutLA.scala 92:29]
  wire [31:0] mag_mux_1_auto_stream_out_1_bits_data; // @[SpectrometerTestWithoutLA.scala 92:29]
  wire  mag_mux_1_auto_stream_out_1_bits_last; // @[SpectrometerTestWithoutLA.scala 92:29]
  wire  acc_clock; // @[SpectrometerTestWithoutLA.scala 98:29]
  wire  acc_reset; // @[SpectrometerTestWithoutLA.scala 98:29]
  wire  acc_auto_bus_in_aw_ready; // @[SpectrometerTestWithoutLA.scala 98:29]
  wire  acc_auto_bus_in_aw_valid; // @[SpectrometerTestWithoutLA.scala 98:29]
  wire  acc_auto_bus_in_aw_bits_id; // @[SpectrometerTestWithoutLA.scala 98:29]
  wire [29:0] acc_auto_bus_in_aw_bits_addr; // @[SpectrometerTestWithoutLA.scala 98:29]
  wire [2:0] acc_auto_bus_in_aw_bits_size; // @[SpectrometerTestWithoutLA.scala 98:29]
  wire  acc_auto_bus_in_w_ready; // @[SpectrometerTestWithoutLA.scala 98:29]
  wire  acc_auto_bus_in_w_valid; // @[SpectrometerTestWithoutLA.scala 98:29]
  wire [31:0] acc_auto_bus_in_w_bits_data; // @[SpectrometerTestWithoutLA.scala 98:29]
  wire [3:0] acc_auto_bus_in_w_bits_strb; // @[SpectrometerTestWithoutLA.scala 98:29]
  wire  acc_auto_bus_in_w_bits_last; // @[SpectrometerTestWithoutLA.scala 98:29]
  wire  acc_auto_bus_in_b_ready; // @[SpectrometerTestWithoutLA.scala 98:29]
  wire  acc_auto_bus_in_b_valid; // @[SpectrometerTestWithoutLA.scala 98:29]
  wire [1:0] acc_auto_bus_in_b_bits_resp; // @[SpectrometerTestWithoutLA.scala 98:29]
  wire  acc_auto_bus_in_ar_ready; // @[SpectrometerTestWithoutLA.scala 98:29]
  wire  acc_auto_bus_in_ar_valid; // @[SpectrometerTestWithoutLA.scala 98:29]
  wire  acc_auto_bus_in_ar_bits_id; // @[SpectrometerTestWithoutLA.scala 98:29]
  wire [29:0] acc_auto_bus_in_ar_bits_addr; // @[SpectrometerTestWithoutLA.scala 98:29]
  wire [2:0] acc_auto_bus_in_ar_bits_size; // @[SpectrometerTestWithoutLA.scala 98:29]
  wire  acc_auto_bus_in_r_ready; // @[SpectrometerTestWithoutLA.scala 98:29]
  wire  acc_auto_bus_in_r_valid; // @[SpectrometerTestWithoutLA.scala 98:29]
  wire [31:0] acc_auto_bus_in_r_bits_data; // @[SpectrometerTestWithoutLA.scala 98:29]
  wire [1:0] acc_auto_bus_in_r_bits_resp; // @[SpectrometerTestWithoutLA.scala 98:29]
  wire  acc_auto_bus_in_r_bits_last; // @[SpectrometerTestWithoutLA.scala 98:29]
  wire  acc_auto_dspQueue_stream_out_ready; // @[SpectrometerTestWithoutLA.scala 98:29]
  wire  acc_auto_dspQueue_stream_out_valid; // @[SpectrometerTestWithoutLA.scala 98:29]
  wire [15:0] acc_auto_dspQueue_stream_out_bits_data; // @[SpectrometerTestWithoutLA.scala 98:29]
  wire  acc_auto_dspQueue_stream_out_bits_last; // @[SpectrometerTestWithoutLA.scala 98:29]
  wire  acc_auto_accumulator_slave_in_ready; // @[SpectrometerTestWithoutLA.scala 98:29]
  wire  acc_auto_accumulator_slave_in_valid; // @[SpectrometerTestWithoutLA.scala 98:29]
  wire [31:0] acc_auto_accumulator_slave_in_bits_data; // @[SpectrometerTestWithoutLA.scala 98:29]
  wire  acc_auto_accumulator_slave_in_bits_last; // @[SpectrometerTestWithoutLA.scala 98:29]
  wire  widthAdapter_1_clock; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_1_reset; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_1_auto_in_ready; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_1_auto_in_valid; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire [15:0] widthAdapter_1_auto_in_bits_data; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_1_auto_in_bits_last; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_1_auto_out_ready; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_1_auto_out_valid; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire [31:0] widthAdapter_1_auto_out_bits_data; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_1_auto_out_bits_last; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  acc_queue_clock; // @[SpectrometerTestWithoutLA.scala 100:29]
  wire  acc_queue_reset; // @[SpectrometerTestWithoutLA.scala 100:29]
  wire  acc_queue_auto_out_out_ready; // @[SpectrometerTestWithoutLA.scala 100:29]
  wire  acc_queue_auto_out_out_valid; // @[SpectrometerTestWithoutLA.scala 100:29]
  wire [31:0] acc_queue_auto_out_out_bits_data; // @[SpectrometerTestWithoutLA.scala 100:29]
  wire  acc_queue_auto_out_out_bits_last; // @[SpectrometerTestWithoutLA.scala 100:29]
  wire  acc_queue_auto_in_in_ready; // @[SpectrometerTestWithoutLA.scala 100:29]
  wire  acc_queue_auto_in_in_valid; // @[SpectrometerTestWithoutLA.scala 100:29]
  wire [31:0] acc_queue_auto_in_in_bits_data; // @[SpectrometerTestWithoutLA.scala 100:29]
  wire  acc_queue_auto_in_in_bits_last; // @[SpectrometerTestWithoutLA.scala 100:29]
  wire  out_mux_clock; // @[SpectrometerTestWithoutLA.scala 102:29]
  wire  out_mux_reset; // @[SpectrometerTestWithoutLA.scala 102:29]
  wire  out_mux_auto_register_in_aw_ready; // @[SpectrometerTestWithoutLA.scala 102:29]
  wire  out_mux_auto_register_in_aw_valid; // @[SpectrometerTestWithoutLA.scala 102:29]
  wire  out_mux_auto_register_in_aw_bits_id; // @[SpectrometerTestWithoutLA.scala 102:29]
  wire [29:0] out_mux_auto_register_in_aw_bits_addr; // @[SpectrometerTestWithoutLA.scala 102:29]
  wire  out_mux_auto_register_in_w_ready; // @[SpectrometerTestWithoutLA.scala 102:29]
  wire  out_mux_auto_register_in_w_valid; // @[SpectrometerTestWithoutLA.scala 102:29]
  wire [31:0] out_mux_auto_register_in_w_bits_data; // @[SpectrometerTestWithoutLA.scala 102:29]
  wire [3:0] out_mux_auto_register_in_w_bits_strb; // @[SpectrometerTestWithoutLA.scala 102:29]
  wire  out_mux_auto_register_in_b_ready; // @[SpectrometerTestWithoutLA.scala 102:29]
  wire  out_mux_auto_register_in_b_valid; // @[SpectrometerTestWithoutLA.scala 102:29]
  wire  out_mux_auto_register_in_b_bits_id; // @[SpectrometerTestWithoutLA.scala 102:29]
  wire  out_mux_auto_register_in_ar_ready; // @[SpectrometerTestWithoutLA.scala 102:29]
  wire  out_mux_auto_register_in_ar_valid; // @[SpectrometerTestWithoutLA.scala 102:29]
  wire  out_mux_auto_register_in_ar_bits_id; // @[SpectrometerTestWithoutLA.scala 102:29]
  wire [29:0] out_mux_auto_register_in_ar_bits_addr; // @[SpectrometerTestWithoutLA.scala 102:29]
  wire [2:0] out_mux_auto_register_in_ar_bits_size; // @[SpectrometerTestWithoutLA.scala 102:29]
  wire  out_mux_auto_register_in_r_ready; // @[SpectrometerTestWithoutLA.scala 102:29]
  wire  out_mux_auto_register_in_r_valid; // @[SpectrometerTestWithoutLA.scala 102:29]
  wire  out_mux_auto_register_in_r_bits_id; // @[SpectrometerTestWithoutLA.scala 102:29]
  wire [31:0] out_mux_auto_register_in_r_bits_data; // @[SpectrometerTestWithoutLA.scala 102:29]
  wire  out_mux_auto_stream_in_6_ready; // @[SpectrometerTestWithoutLA.scala 102:29]
  wire  out_mux_auto_stream_in_6_valid; // @[SpectrometerTestWithoutLA.scala 102:29]
  wire [31:0] out_mux_auto_stream_in_6_bits_data; // @[SpectrometerTestWithoutLA.scala 102:29]
  wire  out_mux_auto_stream_in_6_bits_last; // @[SpectrometerTestWithoutLA.scala 102:29]
  wire  out_mux_auto_stream_in_5_ready; // @[SpectrometerTestWithoutLA.scala 102:29]
  wire  out_mux_auto_stream_in_5_valid; // @[SpectrometerTestWithoutLA.scala 102:29]
  wire [31:0] out_mux_auto_stream_in_5_bits_data; // @[SpectrometerTestWithoutLA.scala 102:29]
  wire  out_mux_auto_stream_in_5_bits_last; // @[SpectrometerTestWithoutLA.scala 102:29]
  wire  out_mux_auto_stream_in_4_ready; // @[SpectrometerTestWithoutLA.scala 102:29]
  wire  out_mux_auto_stream_in_4_valid; // @[SpectrometerTestWithoutLA.scala 102:29]
  wire [31:0] out_mux_auto_stream_in_4_bits_data; // @[SpectrometerTestWithoutLA.scala 102:29]
  wire  out_mux_auto_stream_in_4_bits_last; // @[SpectrometerTestWithoutLA.scala 102:29]
  wire  out_mux_auto_stream_in_3_ready; // @[SpectrometerTestWithoutLA.scala 102:29]
  wire  out_mux_auto_stream_in_3_valid; // @[SpectrometerTestWithoutLA.scala 102:29]
  wire [31:0] out_mux_auto_stream_in_3_bits_data; // @[SpectrometerTestWithoutLA.scala 102:29]
  wire  out_mux_auto_stream_in_3_bits_last; // @[SpectrometerTestWithoutLA.scala 102:29]
  wire  out_mux_auto_stream_in_2_ready; // @[SpectrometerTestWithoutLA.scala 102:29]
  wire  out_mux_auto_stream_in_2_valid; // @[SpectrometerTestWithoutLA.scala 102:29]
  wire [31:0] out_mux_auto_stream_in_2_bits_data; // @[SpectrometerTestWithoutLA.scala 102:29]
  wire  out_mux_auto_stream_in_2_bits_last; // @[SpectrometerTestWithoutLA.scala 102:29]
  wire  out_mux_auto_stream_in_1_ready; // @[SpectrometerTestWithoutLA.scala 102:29]
  wire  out_mux_auto_stream_in_1_valid; // @[SpectrometerTestWithoutLA.scala 102:29]
  wire [31:0] out_mux_auto_stream_in_1_bits_data; // @[SpectrometerTestWithoutLA.scala 102:29]
  wire  out_mux_auto_stream_in_1_bits_last; // @[SpectrometerTestWithoutLA.scala 102:29]
  wire  out_mux_auto_stream_in_0_ready; // @[SpectrometerTestWithoutLA.scala 102:29]
  wire  out_mux_auto_stream_in_0_valid; // @[SpectrometerTestWithoutLA.scala 102:29]
  wire [31:0] out_mux_auto_stream_in_0_bits_data; // @[SpectrometerTestWithoutLA.scala 102:29]
  wire  out_mux_auto_stream_in_0_bits_last; // @[SpectrometerTestWithoutLA.scala 102:29]
  wire  out_mux_auto_stream_out_1_ready; // @[SpectrometerTestWithoutLA.scala 102:29]
  wire  out_mux_auto_stream_out_1_valid; // @[SpectrometerTestWithoutLA.scala 102:29]
  wire [31:0] out_mux_auto_stream_out_1_bits_data; // @[SpectrometerTestWithoutLA.scala 102:29]
  wire  out_mux_auto_stream_out_1_bits_last; // @[SpectrometerTestWithoutLA.scala 102:29]
  wire  out_mux_auto_stream_out_0_ready; // @[SpectrometerTestWithoutLA.scala 102:29]
  wire  out_mux_auto_stream_out_0_valid; // @[SpectrometerTestWithoutLA.scala 102:29]
  wire [31:0] out_mux_auto_stream_out_0_bits_data; // @[SpectrometerTestWithoutLA.scala 102:29]
  wire  out_mux_auto_stream_out_0_bits_last; // @[SpectrometerTestWithoutLA.scala 102:29]
  wire  out_split_clock; // @[SpectrometerTestWithoutLA.scala 103:29]
  wire  out_split_reset; // @[SpectrometerTestWithoutLA.scala 103:29]
  wire  out_split_auto_mem_in_aw_ready; // @[SpectrometerTestWithoutLA.scala 103:29]
  wire  out_split_auto_mem_in_aw_valid; // @[SpectrometerTestWithoutLA.scala 103:29]
  wire  out_split_auto_mem_in_aw_bits_id; // @[SpectrometerTestWithoutLA.scala 103:29]
  wire [29:0] out_split_auto_mem_in_aw_bits_addr; // @[SpectrometerTestWithoutLA.scala 103:29]
  wire  out_split_auto_mem_in_w_ready; // @[SpectrometerTestWithoutLA.scala 103:29]
  wire  out_split_auto_mem_in_w_valid; // @[SpectrometerTestWithoutLA.scala 103:29]
  wire [31:0] out_split_auto_mem_in_w_bits_data; // @[SpectrometerTestWithoutLA.scala 103:29]
  wire [3:0] out_split_auto_mem_in_w_bits_strb; // @[SpectrometerTestWithoutLA.scala 103:29]
  wire  out_split_auto_mem_in_b_ready; // @[SpectrometerTestWithoutLA.scala 103:29]
  wire  out_split_auto_mem_in_b_valid; // @[SpectrometerTestWithoutLA.scala 103:29]
  wire  out_split_auto_mem_in_b_bits_id; // @[SpectrometerTestWithoutLA.scala 103:29]
  wire  out_split_auto_mem_in_ar_ready; // @[SpectrometerTestWithoutLA.scala 103:29]
  wire  out_split_auto_mem_in_ar_valid; // @[SpectrometerTestWithoutLA.scala 103:29]
  wire  out_split_auto_mem_in_ar_bits_id; // @[SpectrometerTestWithoutLA.scala 103:29]
  wire [29:0] out_split_auto_mem_in_ar_bits_addr; // @[SpectrometerTestWithoutLA.scala 103:29]
  wire [2:0] out_split_auto_mem_in_ar_bits_size; // @[SpectrometerTestWithoutLA.scala 103:29]
  wire  out_split_auto_mem_in_r_ready; // @[SpectrometerTestWithoutLA.scala 103:29]
  wire  out_split_auto_mem_in_r_valid; // @[SpectrometerTestWithoutLA.scala 103:29]
  wire  out_split_auto_mem_in_r_bits_id; // @[SpectrometerTestWithoutLA.scala 103:29]
  wire [31:0] out_split_auto_mem_in_r_bits_data; // @[SpectrometerTestWithoutLA.scala 103:29]
  wire  out_split_auto_stream_in_ready; // @[SpectrometerTestWithoutLA.scala 103:29]
  wire  out_split_auto_stream_in_valid; // @[SpectrometerTestWithoutLA.scala 103:29]
  wire [31:0] out_split_auto_stream_in_bits_data; // @[SpectrometerTestWithoutLA.scala 103:29]
  wire  out_split_auto_stream_in_bits_last; // @[SpectrometerTestWithoutLA.scala 103:29]
  wire  out_split_auto_stream_out_ready; // @[SpectrometerTestWithoutLA.scala 103:29]
  wire  out_split_auto_stream_out_valid; // @[SpectrometerTestWithoutLA.scala 103:29]
  wire [31:0] out_split_auto_stream_out_bits_data; // @[SpectrometerTestWithoutLA.scala 103:29]
  wire  out_split_auto_stream_out_bits_last; // @[SpectrometerTestWithoutLA.scala 103:29]
  wire  out_queue_clock; // @[SpectrometerTestWithoutLA.scala 104:29]
  wire  out_queue_reset; // @[SpectrometerTestWithoutLA.scala 104:29]
  wire  out_queue_auto_out_out_ready; // @[SpectrometerTestWithoutLA.scala 104:29]
  wire  out_queue_auto_out_out_valid; // @[SpectrometerTestWithoutLA.scala 104:29]
  wire [31:0] out_queue_auto_out_out_bits_data; // @[SpectrometerTestWithoutLA.scala 104:29]
  wire  out_queue_auto_out_out_bits_last; // @[SpectrometerTestWithoutLA.scala 104:29]
  wire  out_queue_auto_in_in_ready; // @[SpectrometerTestWithoutLA.scala 104:29]
  wire  out_queue_auto_in_in_valid; // @[SpectrometerTestWithoutLA.scala 104:29]
  wire [31:0] out_queue_auto_in_in_bits_data; // @[SpectrometerTestWithoutLA.scala 104:29]
  wire  out_queue_auto_in_in_bits_last; // @[SpectrometerTestWithoutLA.scala 104:29]
  wire  widthAdapter_2_clock; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_2_reset; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_2_auto_in_ready; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_2_auto_in_valid; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire [31:0] widthAdapter_2_auto_in_bits_data; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_2_auto_in_bits_last; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_2_auto_out_ready; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_2_auto_out_valid; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire [7:0] widthAdapter_2_auto_out_bits_data; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_2_auto_out_bits_last; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  uTx_queue_clock; // @[SpectrometerTestWithoutLA.scala 108:29]
  wire  uTx_queue_reset; // @[SpectrometerTestWithoutLA.scala 108:29]
  wire  uTx_queue_auto_out_out_ready; // @[SpectrometerTestWithoutLA.scala 108:29]
  wire  uTx_queue_auto_out_out_valid; // @[SpectrometerTestWithoutLA.scala 108:29]
  wire [31:0] uTx_queue_auto_out_out_bits_data; // @[SpectrometerTestWithoutLA.scala 108:29]
  wire  uTx_queue_auto_out_out_bits_last; // @[SpectrometerTestWithoutLA.scala 108:29]
  wire  uTx_queue_auto_in_in_ready; // @[SpectrometerTestWithoutLA.scala 108:29]
  wire  uTx_queue_auto_in_in_valid; // @[SpectrometerTestWithoutLA.scala 108:29]
  wire [31:0] uTx_queue_auto_in_in_bits_data; // @[SpectrometerTestWithoutLA.scala 108:29]
  wire  uTx_queue_auto_in_in_bits_last; // @[SpectrometerTestWithoutLA.scala 108:29]
  wire  widthAdapter_3_clock; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_3_reset; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_3_auto_in_ready; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_3_auto_in_valid; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire [31:0] widthAdapter_3_auto_in_bits_data; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_3_auto_in_bits_last; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_3_auto_out_ready; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_3_auto_out_valid; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire [7:0] widthAdapter_3_auto_out_bits_data; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_3_auto_out_bits_last; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_4_clock; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_4_reset; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_4_auto_in_ready; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_4_auto_in_valid; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire [7:0] widthAdapter_4_auto_in_bits_data; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_4_auto_in_bits_last; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_4_auto_out_ready; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_4_auto_out_valid; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire [31:0] widthAdapter_4_auto_out_bits_data; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_4_auto_out_bits_last; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  uRx_split_clock; // @[SpectrometerTestWithoutLA.scala 111:29]
  wire  uRx_split_reset; // @[SpectrometerTestWithoutLA.scala 111:29]
  wire  uRx_split_auto_mem_in_aw_ready; // @[SpectrometerTestWithoutLA.scala 111:29]
  wire  uRx_split_auto_mem_in_aw_valid; // @[SpectrometerTestWithoutLA.scala 111:29]
  wire  uRx_split_auto_mem_in_aw_bits_id; // @[SpectrometerTestWithoutLA.scala 111:29]
  wire [29:0] uRx_split_auto_mem_in_aw_bits_addr; // @[SpectrometerTestWithoutLA.scala 111:29]
  wire  uRx_split_auto_mem_in_w_ready; // @[SpectrometerTestWithoutLA.scala 111:29]
  wire  uRx_split_auto_mem_in_w_valid; // @[SpectrometerTestWithoutLA.scala 111:29]
  wire [31:0] uRx_split_auto_mem_in_w_bits_data; // @[SpectrometerTestWithoutLA.scala 111:29]
  wire [3:0] uRx_split_auto_mem_in_w_bits_strb; // @[SpectrometerTestWithoutLA.scala 111:29]
  wire  uRx_split_auto_mem_in_b_ready; // @[SpectrometerTestWithoutLA.scala 111:29]
  wire  uRx_split_auto_mem_in_b_valid; // @[SpectrometerTestWithoutLA.scala 111:29]
  wire  uRx_split_auto_mem_in_b_bits_id; // @[SpectrometerTestWithoutLA.scala 111:29]
  wire  uRx_split_auto_mem_in_ar_ready; // @[SpectrometerTestWithoutLA.scala 111:29]
  wire  uRx_split_auto_mem_in_ar_valid; // @[SpectrometerTestWithoutLA.scala 111:29]
  wire  uRx_split_auto_mem_in_ar_bits_id; // @[SpectrometerTestWithoutLA.scala 111:29]
  wire [29:0] uRx_split_auto_mem_in_ar_bits_addr; // @[SpectrometerTestWithoutLA.scala 111:29]
  wire [2:0] uRx_split_auto_mem_in_ar_bits_size; // @[SpectrometerTestWithoutLA.scala 111:29]
  wire  uRx_split_auto_mem_in_r_ready; // @[SpectrometerTestWithoutLA.scala 111:29]
  wire  uRx_split_auto_mem_in_r_valid; // @[SpectrometerTestWithoutLA.scala 111:29]
  wire  uRx_split_auto_mem_in_r_bits_id; // @[SpectrometerTestWithoutLA.scala 111:29]
  wire [31:0] uRx_split_auto_mem_in_r_bits_data; // @[SpectrometerTestWithoutLA.scala 111:29]
  wire  uRx_split_auto_stream_in_ready; // @[SpectrometerTestWithoutLA.scala 111:29]
  wire  uRx_split_auto_stream_in_valid; // @[SpectrometerTestWithoutLA.scala 111:29]
  wire [31:0] uRx_split_auto_stream_in_bits_data; // @[SpectrometerTestWithoutLA.scala 111:29]
  wire  uRx_split_auto_stream_in_bits_last; // @[SpectrometerTestWithoutLA.scala 111:29]
  wire  uRx_split_auto_stream_out_4_ready; // @[SpectrometerTestWithoutLA.scala 111:29]
  wire  uRx_split_auto_stream_out_4_valid; // @[SpectrometerTestWithoutLA.scala 111:29]
  wire [31:0] uRx_split_auto_stream_out_4_bits_data; // @[SpectrometerTestWithoutLA.scala 111:29]
  wire  uRx_split_auto_stream_out_4_bits_last; // @[SpectrometerTestWithoutLA.scala 111:29]
  wire  uRx_split_auto_stream_out_3_ready; // @[SpectrometerTestWithoutLA.scala 111:29]
  wire  uRx_split_auto_stream_out_3_valid; // @[SpectrometerTestWithoutLA.scala 111:29]
  wire [31:0] uRx_split_auto_stream_out_3_bits_data; // @[SpectrometerTestWithoutLA.scala 111:29]
  wire  uRx_split_auto_stream_out_3_bits_last; // @[SpectrometerTestWithoutLA.scala 111:29]
  wire  uRx_split_auto_stream_out_2_ready; // @[SpectrometerTestWithoutLA.scala 111:29]
  wire  uRx_split_auto_stream_out_2_valid; // @[SpectrometerTestWithoutLA.scala 111:29]
  wire [31:0] uRx_split_auto_stream_out_2_bits_data; // @[SpectrometerTestWithoutLA.scala 111:29]
  wire  uRx_split_auto_stream_out_2_bits_last; // @[SpectrometerTestWithoutLA.scala 111:29]
  wire  uRx_split_auto_stream_out_1_ready; // @[SpectrometerTestWithoutLA.scala 111:29]
  wire  uRx_split_auto_stream_out_1_valid; // @[SpectrometerTestWithoutLA.scala 111:29]
  wire [31:0] uRx_split_auto_stream_out_1_bits_data; // @[SpectrometerTestWithoutLA.scala 111:29]
  wire  uRx_split_auto_stream_out_1_bits_last; // @[SpectrometerTestWithoutLA.scala 111:29]
  wire  uRx_split_auto_stream_out_0_ready; // @[SpectrometerTestWithoutLA.scala 111:29]
  wire  uRx_split_auto_stream_out_0_valid; // @[SpectrometerTestWithoutLA.scala 111:29]
  wire [31:0] uRx_split_auto_stream_out_0_bits_data; // @[SpectrometerTestWithoutLA.scala 111:29]
  wire  uRx_split_auto_stream_out_0_bits_last; // @[SpectrometerTestWithoutLA.scala 111:29]
  wire  uart_clock; // @[SpectrometerTestWithoutLA.scala 112:29]
  wire  uart_reset; // @[SpectrometerTestWithoutLA.scala 112:29]
  wire  uart_auto_mem_in_aw_ready; // @[SpectrometerTestWithoutLA.scala 112:29]
  wire  uart_auto_mem_in_aw_valid; // @[SpectrometerTestWithoutLA.scala 112:29]
  wire  uart_auto_mem_in_aw_bits_id; // @[SpectrometerTestWithoutLA.scala 112:29]
  wire [29:0] uart_auto_mem_in_aw_bits_addr; // @[SpectrometerTestWithoutLA.scala 112:29]
  wire  uart_auto_mem_in_w_ready; // @[SpectrometerTestWithoutLA.scala 112:29]
  wire  uart_auto_mem_in_w_valid; // @[SpectrometerTestWithoutLA.scala 112:29]
  wire [31:0] uart_auto_mem_in_w_bits_data; // @[SpectrometerTestWithoutLA.scala 112:29]
  wire [3:0] uart_auto_mem_in_w_bits_strb; // @[SpectrometerTestWithoutLA.scala 112:29]
  wire  uart_auto_mem_in_b_ready; // @[SpectrometerTestWithoutLA.scala 112:29]
  wire  uart_auto_mem_in_b_valid; // @[SpectrometerTestWithoutLA.scala 112:29]
  wire  uart_auto_mem_in_b_bits_id; // @[SpectrometerTestWithoutLA.scala 112:29]
  wire  uart_auto_mem_in_ar_ready; // @[SpectrometerTestWithoutLA.scala 112:29]
  wire  uart_auto_mem_in_ar_valid; // @[SpectrometerTestWithoutLA.scala 112:29]
  wire  uart_auto_mem_in_ar_bits_id; // @[SpectrometerTestWithoutLA.scala 112:29]
  wire [29:0] uart_auto_mem_in_ar_bits_addr; // @[SpectrometerTestWithoutLA.scala 112:29]
  wire [2:0] uart_auto_mem_in_ar_bits_size; // @[SpectrometerTestWithoutLA.scala 112:29]
  wire  uart_auto_mem_in_r_ready; // @[SpectrometerTestWithoutLA.scala 112:29]
  wire  uart_auto_mem_in_r_valid; // @[SpectrometerTestWithoutLA.scala 112:29]
  wire  uart_auto_mem_in_r_bits_id; // @[SpectrometerTestWithoutLA.scala 112:29]
  wire [31:0] uart_auto_mem_in_r_bits_data; // @[SpectrometerTestWithoutLA.scala 112:29]
  wire  uart_auto_in_in_ready; // @[SpectrometerTestWithoutLA.scala 112:29]
  wire  uart_auto_in_in_valid; // @[SpectrometerTestWithoutLA.scala 112:29]
  wire [7:0] uart_auto_in_in_bits_data; // @[SpectrometerTestWithoutLA.scala 112:29]
  wire  uart_auto_out_out_ready; // @[SpectrometerTestWithoutLA.scala 112:29]
  wire  uart_auto_out_out_valid; // @[SpectrometerTestWithoutLA.scala 112:29]
  wire [7:0] uart_auto_out_out_bits_data; // @[SpectrometerTestWithoutLA.scala 112:29]
  wire  uart_int_0; // @[SpectrometerTestWithoutLA.scala 112:29]
  wire  uart_io_txd; // @[SpectrometerTestWithoutLA.scala 112:29]
  wire  uart_io_rxd; // @[SpectrometerTestWithoutLA.scala 112:29]
  wire  bus_clock; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_reset; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_in_aw_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_in_aw_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_in_aw_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [29:0] bus_auto_in_aw_bits_addr; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [2:0] bus_auto_in_aw_bits_size; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_in_w_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_in_w_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [31:0] bus_auto_in_w_bits_data; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [3:0] bus_auto_in_w_bits_strb; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_in_w_bits_last; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_in_b_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_in_b_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [1:0] bus_auto_in_b_bits_resp; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_in_ar_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_in_ar_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_in_ar_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [29:0] bus_auto_in_ar_bits_addr; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [2:0] bus_auto_in_ar_bits_size; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_in_r_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_in_r_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [31:0] bus_auto_in_r_bits_data; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [1:0] bus_auto_in_r_bits_resp; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_in_r_bits_last; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_21_aw_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_21_aw_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_21_aw_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [29:0] bus_auto_out_21_aw_bits_addr; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [2:0] bus_auto_out_21_aw_bits_size; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_21_w_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_21_w_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [31:0] bus_auto_out_21_w_bits_data; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [3:0] bus_auto_out_21_w_bits_strb; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_21_w_bits_last; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_21_b_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_21_b_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [1:0] bus_auto_out_21_b_bits_resp; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_21_ar_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_21_ar_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_21_ar_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [29:0] bus_auto_out_21_ar_bits_addr; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [2:0] bus_auto_out_21_ar_bits_size; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_21_r_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_21_r_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [31:0] bus_auto_out_21_r_bits_data; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [1:0] bus_auto_out_21_r_bits_resp; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_21_r_bits_last; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_20_aw_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_20_aw_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_20_aw_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [29:0] bus_auto_out_20_aw_bits_addr; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [2:0] bus_auto_out_20_aw_bits_size; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_20_w_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_20_w_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [31:0] bus_auto_out_20_w_bits_data; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [3:0] bus_auto_out_20_w_bits_strb; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_20_w_bits_last; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_20_b_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_20_b_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_20_b_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [1:0] bus_auto_out_20_b_bits_resp; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_20_ar_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_20_ar_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_20_ar_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [29:0] bus_auto_out_20_ar_bits_addr; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [2:0] bus_auto_out_20_ar_bits_size; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_20_r_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_20_r_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_20_r_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [31:0] bus_auto_out_20_r_bits_data; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [1:0] bus_auto_out_20_r_bits_resp; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_20_r_bits_last; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_19_aw_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_19_aw_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_19_aw_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [29:0] bus_auto_out_19_aw_bits_addr; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [2:0] bus_auto_out_19_aw_bits_size; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_19_w_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_19_w_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [31:0] bus_auto_out_19_w_bits_data; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [3:0] bus_auto_out_19_w_bits_strb; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_19_w_bits_last; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_19_b_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_19_b_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_19_b_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [1:0] bus_auto_out_19_b_bits_resp; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_19_ar_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_19_ar_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_19_ar_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [29:0] bus_auto_out_19_ar_bits_addr; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [2:0] bus_auto_out_19_ar_bits_size; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_19_r_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_19_r_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_19_r_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [31:0] bus_auto_out_19_r_bits_data; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [1:0] bus_auto_out_19_r_bits_resp; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_19_r_bits_last; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_18_aw_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_18_aw_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_18_aw_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [29:0] bus_auto_out_18_aw_bits_addr; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [2:0] bus_auto_out_18_aw_bits_size; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_18_w_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_18_w_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [31:0] bus_auto_out_18_w_bits_data; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [3:0] bus_auto_out_18_w_bits_strb; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_18_w_bits_last; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_18_b_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_18_b_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_18_b_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [1:0] bus_auto_out_18_b_bits_resp; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_18_ar_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_18_ar_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_18_ar_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [29:0] bus_auto_out_18_ar_bits_addr; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [2:0] bus_auto_out_18_ar_bits_size; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_18_r_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_18_r_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_18_r_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [31:0] bus_auto_out_18_r_bits_data; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [1:0] bus_auto_out_18_r_bits_resp; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_18_r_bits_last; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_17_aw_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_17_aw_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_17_aw_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [29:0] bus_auto_out_17_aw_bits_addr; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [2:0] bus_auto_out_17_aw_bits_size; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_17_w_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_17_w_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [31:0] bus_auto_out_17_w_bits_data; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [3:0] bus_auto_out_17_w_bits_strb; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_17_w_bits_last; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_17_b_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_17_b_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_17_b_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [1:0] bus_auto_out_17_b_bits_resp; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_17_ar_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_17_ar_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_17_ar_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [29:0] bus_auto_out_17_ar_bits_addr; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [2:0] bus_auto_out_17_ar_bits_size; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_17_r_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_17_r_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_17_r_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [31:0] bus_auto_out_17_r_bits_data; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [1:0] bus_auto_out_17_r_bits_resp; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_17_r_bits_last; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_16_aw_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_16_aw_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_16_aw_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [29:0] bus_auto_out_16_aw_bits_addr; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [2:0] bus_auto_out_16_aw_bits_size; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_16_w_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_16_w_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [31:0] bus_auto_out_16_w_bits_data; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [3:0] bus_auto_out_16_w_bits_strb; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_16_w_bits_last; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_16_b_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_16_b_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_16_b_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [1:0] bus_auto_out_16_b_bits_resp; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_16_ar_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_16_ar_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_16_ar_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [29:0] bus_auto_out_16_ar_bits_addr; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [2:0] bus_auto_out_16_ar_bits_size; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_16_r_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_16_r_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_16_r_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [31:0] bus_auto_out_16_r_bits_data; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [1:0] bus_auto_out_16_r_bits_resp; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_16_r_bits_last; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_15_aw_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_15_aw_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_15_aw_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [29:0] bus_auto_out_15_aw_bits_addr; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [2:0] bus_auto_out_15_aw_bits_size; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_15_w_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_15_w_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [31:0] bus_auto_out_15_w_bits_data; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [3:0] bus_auto_out_15_w_bits_strb; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_15_w_bits_last; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_15_b_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_15_b_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_15_b_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [1:0] bus_auto_out_15_b_bits_resp; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_15_ar_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_15_ar_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_15_ar_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [29:0] bus_auto_out_15_ar_bits_addr; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [2:0] bus_auto_out_15_ar_bits_size; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_15_r_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_15_r_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_15_r_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [31:0] bus_auto_out_15_r_bits_data; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [1:0] bus_auto_out_15_r_bits_resp; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_15_r_bits_last; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_14_aw_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_14_aw_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_14_aw_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [29:0] bus_auto_out_14_aw_bits_addr; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [2:0] bus_auto_out_14_aw_bits_size; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_14_w_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_14_w_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [31:0] bus_auto_out_14_w_bits_data; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [3:0] bus_auto_out_14_w_bits_strb; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_14_w_bits_last; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_14_b_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_14_b_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_14_b_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [1:0] bus_auto_out_14_b_bits_resp; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_14_ar_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_14_ar_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_14_ar_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [29:0] bus_auto_out_14_ar_bits_addr; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [2:0] bus_auto_out_14_ar_bits_size; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_14_r_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_14_r_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_14_r_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [31:0] bus_auto_out_14_r_bits_data; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [1:0] bus_auto_out_14_r_bits_resp; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_14_r_bits_last; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_13_aw_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_13_aw_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_13_aw_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [29:0] bus_auto_out_13_aw_bits_addr; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [2:0] bus_auto_out_13_aw_bits_size; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_13_w_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_13_w_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [31:0] bus_auto_out_13_w_bits_data; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [3:0] bus_auto_out_13_w_bits_strb; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_13_w_bits_last; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_13_b_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_13_b_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_13_b_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [1:0] bus_auto_out_13_b_bits_resp; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_13_ar_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_13_ar_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_13_ar_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [29:0] bus_auto_out_13_ar_bits_addr; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [2:0] bus_auto_out_13_ar_bits_size; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_13_r_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_13_r_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_13_r_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [31:0] bus_auto_out_13_r_bits_data; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [1:0] bus_auto_out_13_r_bits_resp; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_13_r_bits_last; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_12_aw_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_12_aw_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_12_aw_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [29:0] bus_auto_out_12_aw_bits_addr; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [2:0] bus_auto_out_12_aw_bits_size; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_12_w_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_12_w_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [31:0] bus_auto_out_12_w_bits_data; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [3:0] bus_auto_out_12_w_bits_strb; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_12_w_bits_last; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_12_b_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_12_b_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_12_b_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [1:0] bus_auto_out_12_b_bits_resp; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_12_ar_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_12_ar_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_12_ar_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [29:0] bus_auto_out_12_ar_bits_addr; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [2:0] bus_auto_out_12_ar_bits_size; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_12_r_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_12_r_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_12_r_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [31:0] bus_auto_out_12_r_bits_data; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [1:0] bus_auto_out_12_r_bits_resp; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_12_r_bits_last; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_11_aw_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_11_aw_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_11_aw_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [29:0] bus_auto_out_11_aw_bits_addr; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [2:0] bus_auto_out_11_aw_bits_size; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_11_w_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_11_w_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [31:0] bus_auto_out_11_w_bits_data; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [3:0] bus_auto_out_11_w_bits_strb; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_11_w_bits_last; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_11_b_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_11_b_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_11_b_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [1:0] bus_auto_out_11_b_bits_resp; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_11_ar_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_11_ar_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_11_ar_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [29:0] bus_auto_out_11_ar_bits_addr; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [2:0] bus_auto_out_11_ar_bits_size; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_11_r_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_11_r_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_11_r_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [31:0] bus_auto_out_11_r_bits_data; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [1:0] bus_auto_out_11_r_bits_resp; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_11_r_bits_last; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_10_aw_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_10_aw_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_10_aw_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [29:0] bus_auto_out_10_aw_bits_addr; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [2:0] bus_auto_out_10_aw_bits_size; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_10_w_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_10_w_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [31:0] bus_auto_out_10_w_bits_data; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [3:0] bus_auto_out_10_w_bits_strb; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_10_w_bits_last; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_10_b_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_10_b_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_10_b_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [1:0] bus_auto_out_10_b_bits_resp; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_10_ar_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_10_ar_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_10_ar_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [29:0] bus_auto_out_10_ar_bits_addr; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [2:0] bus_auto_out_10_ar_bits_size; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_10_r_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_10_r_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_10_r_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [31:0] bus_auto_out_10_r_bits_data; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [1:0] bus_auto_out_10_r_bits_resp; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_10_r_bits_last; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_9_aw_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_9_aw_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_9_aw_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [29:0] bus_auto_out_9_aw_bits_addr; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [2:0] bus_auto_out_9_aw_bits_size; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_9_w_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_9_w_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [31:0] bus_auto_out_9_w_bits_data; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [3:0] bus_auto_out_9_w_bits_strb; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_9_w_bits_last; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_9_b_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_9_b_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_9_b_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [1:0] bus_auto_out_9_b_bits_resp; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_9_ar_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_9_ar_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_9_ar_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [29:0] bus_auto_out_9_ar_bits_addr; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [2:0] bus_auto_out_9_ar_bits_size; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_9_r_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_9_r_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_9_r_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [31:0] bus_auto_out_9_r_bits_data; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [1:0] bus_auto_out_9_r_bits_resp; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_9_r_bits_last; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_8_aw_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_8_aw_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_8_aw_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [29:0] bus_auto_out_8_aw_bits_addr; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [2:0] bus_auto_out_8_aw_bits_size; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_8_w_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_8_w_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [31:0] bus_auto_out_8_w_bits_data; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [3:0] bus_auto_out_8_w_bits_strb; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_8_w_bits_last; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_8_b_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_8_b_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_8_b_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [1:0] bus_auto_out_8_b_bits_resp; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_8_ar_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_8_ar_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_8_ar_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [29:0] bus_auto_out_8_ar_bits_addr; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [2:0] bus_auto_out_8_ar_bits_size; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_8_r_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_8_r_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_8_r_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [31:0] bus_auto_out_8_r_bits_data; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [1:0] bus_auto_out_8_r_bits_resp; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_8_r_bits_last; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_7_aw_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_7_aw_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_7_aw_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [29:0] bus_auto_out_7_aw_bits_addr; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [2:0] bus_auto_out_7_aw_bits_size; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_7_w_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_7_w_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [31:0] bus_auto_out_7_w_bits_data; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [3:0] bus_auto_out_7_w_bits_strb; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_7_w_bits_last; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_7_b_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_7_b_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_7_b_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [1:0] bus_auto_out_7_b_bits_resp; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_7_ar_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_7_ar_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_7_ar_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [29:0] bus_auto_out_7_ar_bits_addr; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [2:0] bus_auto_out_7_ar_bits_size; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_7_r_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_7_r_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_7_r_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [31:0] bus_auto_out_7_r_bits_data; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [1:0] bus_auto_out_7_r_bits_resp; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_7_r_bits_last; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_6_aw_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_6_aw_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_6_aw_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [29:0] bus_auto_out_6_aw_bits_addr; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [2:0] bus_auto_out_6_aw_bits_size; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_6_w_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_6_w_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [31:0] bus_auto_out_6_w_bits_data; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [3:0] bus_auto_out_6_w_bits_strb; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_6_w_bits_last; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_6_b_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_6_b_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_6_b_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [1:0] bus_auto_out_6_b_bits_resp; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_6_ar_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_6_ar_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_6_ar_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [29:0] bus_auto_out_6_ar_bits_addr; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [2:0] bus_auto_out_6_ar_bits_size; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_6_r_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_6_r_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_6_r_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [31:0] bus_auto_out_6_r_bits_data; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [1:0] bus_auto_out_6_r_bits_resp; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_6_r_bits_last; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_5_aw_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_5_aw_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_5_aw_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [29:0] bus_auto_out_5_aw_bits_addr; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [2:0] bus_auto_out_5_aw_bits_size; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_5_w_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_5_w_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [31:0] bus_auto_out_5_w_bits_data; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [3:0] bus_auto_out_5_w_bits_strb; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_5_w_bits_last; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_5_b_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_5_b_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_5_b_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [1:0] bus_auto_out_5_b_bits_resp; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_5_ar_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_5_ar_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_5_ar_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [29:0] bus_auto_out_5_ar_bits_addr; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [2:0] bus_auto_out_5_ar_bits_size; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_5_r_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_5_r_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_5_r_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [31:0] bus_auto_out_5_r_bits_data; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [1:0] bus_auto_out_5_r_bits_resp; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_5_r_bits_last; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_4_aw_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_4_aw_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_4_aw_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [29:0] bus_auto_out_4_aw_bits_addr; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [2:0] bus_auto_out_4_aw_bits_size; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_4_w_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_4_w_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [31:0] bus_auto_out_4_w_bits_data; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [3:0] bus_auto_out_4_w_bits_strb; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_4_w_bits_last; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_4_b_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_4_b_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_4_b_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [1:0] bus_auto_out_4_b_bits_resp; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_4_ar_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_4_ar_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_4_ar_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [29:0] bus_auto_out_4_ar_bits_addr; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [2:0] bus_auto_out_4_ar_bits_size; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_4_r_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_4_r_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_4_r_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [31:0] bus_auto_out_4_r_bits_data; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [1:0] bus_auto_out_4_r_bits_resp; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_4_r_bits_last; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_3_aw_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_3_aw_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_3_aw_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [29:0] bus_auto_out_3_aw_bits_addr; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [2:0] bus_auto_out_3_aw_bits_size; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_3_w_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_3_w_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [31:0] bus_auto_out_3_w_bits_data; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [3:0] bus_auto_out_3_w_bits_strb; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_3_w_bits_last; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_3_b_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_3_b_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_3_b_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [1:0] bus_auto_out_3_b_bits_resp; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_3_ar_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_3_ar_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_3_ar_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [29:0] bus_auto_out_3_ar_bits_addr; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [2:0] bus_auto_out_3_ar_bits_size; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_3_r_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_3_r_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_3_r_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [31:0] bus_auto_out_3_r_bits_data; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [1:0] bus_auto_out_3_r_bits_resp; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_3_r_bits_last; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_2_aw_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_2_aw_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_2_aw_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [29:0] bus_auto_out_2_aw_bits_addr; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [2:0] bus_auto_out_2_aw_bits_size; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_2_w_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_2_w_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [31:0] bus_auto_out_2_w_bits_data; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [3:0] bus_auto_out_2_w_bits_strb; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_2_w_bits_last; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_2_b_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_2_b_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_2_b_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [1:0] bus_auto_out_2_b_bits_resp; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_2_ar_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_2_ar_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_2_ar_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [29:0] bus_auto_out_2_ar_bits_addr; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [2:0] bus_auto_out_2_ar_bits_size; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_2_r_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_2_r_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_2_r_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [31:0] bus_auto_out_2_r_bits_data; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [1:0] bus_auto_out_2_r_bits_resp; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_2_r_bits_last; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_1_aw_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_1_aw_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_1_aw_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [29:0] bus_auto_out_1_aw_bits_addr; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [2:0] bus_auto_out_1_aw_bits_size; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_1_w_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_1_w_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [31:0] bus_auto_out_1_w_bits_data; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [3:0] bus_auto_out_1_w_bits_strb; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_1_w_bits_last; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_1_b_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_1_b_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_1_b_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [1:0] bus_auto_out_1_b_bits_resp; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_1_ar_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_1_ar_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_1_ar_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [29:0] bus_auto_out_1_ar_bits_addr; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [2:0] bus_auto_out_1_ar_bits_size; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_1_r_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_1_r_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_1_r_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [31:0] bus_auto_out_1_r_bits_data; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [1:0] bus_auto_out_1_r_bits_resp; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_1_r_bits_last; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_0_aw_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_0_aw_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_0_aw_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [29:0] bus_auto_out_0_aw_bits_addr; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [2:0] bus_auto_out_0_aw_bits_size; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_0_w_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_0_w_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [31:0] bus_auto_out_0_w_bits_data; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [3:0] bus_auto_out_0_w_bits_strb; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_0_w_bits_last; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_0_b_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_0_b_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_0_b_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [1:0] bus_auto_out_0_b_bits_resp; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_0_ar_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_0_ar_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_0_ar_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [29:0] bus_auto_out_0_ar_bits_addr; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [2:0] bus_auto_out_0_ar_bits_size; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_0_r_ready; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_0_r_valid; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_0_r_bits_id; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [31:0] bus_auto_out_0_r_bits_data; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire [1:0] bus_auto_out_0_r_bits_resp; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  bus_auto_out_0_r_bits_last; // @[SpectrometerTestWithoutLA.scala 126:23]
  wire  axi4buf_clock; // @[Buffer.scala 58:29]
  wire  axi4buf_reset; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_in_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_in_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_in_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_auto_in_aw_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_auto_in_aw_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_in_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_in_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_auto_in_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_auto_in_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_in_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_in_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_in_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_in_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_auto_in_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_in_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_in_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_in_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_auto_in_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_auto_in_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_in_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_in_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_in_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_auto_in_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_auto_in_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_in_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_out_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_out_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_out_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_auto_out_aw_bits_addr; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_out_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_out_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_auto_out_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_auto_out_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_out_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_out_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_out_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_out_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_auto_out_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_out_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_out_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_out_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_auto_out_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_auto_out_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_out_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_out_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_out_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_auto_out_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_auto_out_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_out_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_1_clock; // @[Buffer.scala 58:29]
  wire  axi4buf_1_reset; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_in_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_in_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_in_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_1_auto_in_aw_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_1_auto_in_aw_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_in_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_in_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_1_auto_in_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_1_auto_in_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_in_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_in_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_in_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_in_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_1_auto_in_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_in_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_in_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_in_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_1_auto_in_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_1_auto_in_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_in_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_in_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_in_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_1_auto_in_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_1_auto_in_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_in_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_out_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_out_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_out_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_1_auto_out_aw_bits_addr; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_out_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_out_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_1_auto_out_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_1_auto_out_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_out_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_out_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_out_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_out_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_1_auto_out_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_out_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_out_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_out_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_1_auto_out_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_1_auto_out_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_out_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_out_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_out_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_1_auto_out_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_1_auto_out_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_out_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_2_clock; // @[Buffer.scala 58:29]
  wire  axi4buf_2_reset; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_in_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_in_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_in_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_2_auto_in_aw_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_2_auto_in_aw_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_in_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_in_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_2_auto_in_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_2_auto_in_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_in_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_in_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_in_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_in_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_2_auto_in_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_in_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_in_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_in_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_2_auto_in_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_2_auto_in_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_in_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_in_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_in_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_2_auto_in_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_2_auto_in_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_in_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_out_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_out_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_out_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_2_auto_out_aw_bits_addr; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_out_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_out_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_2_auto_out_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_2_auto_out_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_out_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_out_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_out_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_out_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_2_auto_out_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_out_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_out_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_out_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_2_auto_out_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_2_auto_out_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_out_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_out_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_out_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_2_auto_out_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_2_auto_out_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_out_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_3_clock; // @[Buffer.scala 58:29]
  wire  axi4buf_3_reset; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_in_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_in_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_in_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_3_auto_in_aw_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_3_auto_in_aw_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_in_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_in_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_3_auto_in_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_3_auto_in_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_in_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_in_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_in_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_in_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_3_auto_in_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_in_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_in_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_in_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_3_auto_in_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_3_auto_in_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_in_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_in_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_in_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_3_auto_in_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_3_auto_in_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_in_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_out_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_out_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_out_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_3_auto_out_aw_bits_addr; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_out_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_out_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_3_auto_out_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_3_auto_out_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_out_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_out_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_out_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_out_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_3_auto_out_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_out_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_out_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_out_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_3_auto_out_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_3_auto_out_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_out_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_out_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_out_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_3_auto_out_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_3_auto_out_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_out_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_4_clock; // @[Buffer.scala 58:29]
  wire  axi4buf_4_reset; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_in_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_in_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_in_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_4_auto_in_aw_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_4_auto_in_aw_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_in_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_in_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_4_auto_in_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_4_auto_in_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_in_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_in_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_in_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_in_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_4_auto_in_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_in_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_in_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_in_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_4_auto_in_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_4_auto_in_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_in_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_in_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_in_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_4_auto_in_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_4_auto_in_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_in_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_out_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_out_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_out_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_4_auto_out_aw_bits_addr; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_out_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_out_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_4_auto_out_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_4_auto_out_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_out_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_out_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_out_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_out_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_4_auto_out_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_out_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_out_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_out_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_4_auto_out_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_4_auto_out_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_out_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_out_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_out_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_4_auto_out_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_4_auto_out_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_out_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_5_clock; // @[Buffer.scala 58:29]
  wire  axi4buf_5_reset; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_in_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_in_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_in_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_5_auto_in_aw_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_5_auto_in_aw_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_in_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_in_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_5_auto_in_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_5_auto_in_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_in_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_in_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_in_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_in_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_5_auto_in_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_in_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_in_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_in_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_5_auto_in_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_5_auto_in_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_in_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_in_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_in_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_5_auto_in_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_5_auto_in_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_in_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_out_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_out_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_out_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_5_auto_out_aw_bits_addr; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_out_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_out_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_5_auto_out_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_5_auto_out_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_out_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_out_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_out_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_out_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_5_auto_out_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_out_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_out_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_out_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_5_auto_out_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_5_auto_out_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_out_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_out_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_out_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_5_auto_out_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_5_auto_out_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_out_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_6_clock; // @[Buffer.scala 58:29]
  wire  axi4buf_6_reset; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_in_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_in_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_in_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_6_auto_in_aw_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_6_auto_in_aw_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_in_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_in_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_6_auto_in_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_6_auto_in_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_in_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_in_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_in_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_in_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_6_auto_in_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_in_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_in_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_in_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_6_auto_in_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_6_auto_in_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_in_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_in_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_in_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_6_auto_in_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_6_auto_in_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_in_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_out_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_out_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_out_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_6_auto_out_aw_bits_addr; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_out_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_out_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_6_auto_out_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_6_auto_out_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_out_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_out_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_out_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_out_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_6_auto_out_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_out_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_out_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_out_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_6_auto_out_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_6_auto_out_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_out_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_out_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_out_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_6_auto_out_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_6_auto_out_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_out_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_7_clock; // @[Buffer.scala 58:29]
  wire  axi4buf_7_reset; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_in_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_in_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_in_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_7_auto_in_aw_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_7_auto_in_aw_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_in_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_in_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_7_auto_in_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_7_auto_in_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_in_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_in_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_in_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_in_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_7_auto_in_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_in_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_in_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_in_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_7_auto_in_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_7_auto_in_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_in_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_in_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_in_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_7_auto_in_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_7_auto_in_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_in_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_out_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_out_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_out_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_7_auto_out_aw_bits_addr; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_out_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_out_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_7_auto_out_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_7_auto_out_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_out_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_out_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_out_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_out_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_7_auto_out_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_out_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_out_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_out_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_7_auto_out_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_7_auto_out_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_out_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_out_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_out_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_7_auto_out_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_7_auto_out_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_out_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_8_clock; // @[Buffer.scala 58:29]
  wire  axi4buf_8_reset; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_in_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_in_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_in_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_8_auto_in_aw_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_8_auto_in_aw_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_in_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_in_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_8_auto_in_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_8_auto_in_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_in_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_in_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_in_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_in_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_8_auto_in_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_in_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_in_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_in_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_8_auto_in_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_8_auto_in_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_in_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_in_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_in_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_8_auto_in_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_8_auto_in_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_in_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_out_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_out_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_out_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_8_auto_out_aw_bits_addr; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_out_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_out_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_8_auto_out_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_8_auto_out_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_out_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_out_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_out_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_out_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_8_auto_out_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_out_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_out_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_out_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_8_auto_out_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_8_auto_out_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_out_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_out_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_out_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_8_auto_out_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_8_auto_out_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_out_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_9_clock; // @[Buffer.scala 58:29]
  wire  axi4buf_9_reset; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_in_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_in_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_in_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_9_auto_in_aw_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_9_auto_in_aw_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_in_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_in_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_9_auto_in_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_9_auto_in_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_in_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_in_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_in_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_in_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_9_auto_in_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_in_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_in_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_in_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_9_auto_in_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_9_auto_in_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_in_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_in_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_in_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_9_auto_in_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_9_auto_in_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_in_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_out_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_out_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_out_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_9_auto_out_aw_bits_addr; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_out_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_out_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_9_auto_out_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_9_auto_out_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_out_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_out_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_out_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_out_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_9_auto_out_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_out_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_out_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_out_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_9_auto_out_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_9_auto_out_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_out_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_out_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_out_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_9_auto_out_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_9_auto_out_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_out_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_10_clock; // @[Buffer.scala 58:29]
  wire  axi4buf_10_reset; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_in_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_in_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_in_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_10_auto_in_aw_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_10_auto_in_aw_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_in_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_in_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_10_auto_in_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_10_auto_in_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_in_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_in_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_in_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_in_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_10_auto_in_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_in_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_in_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_in_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_10_auto_in_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_10_auto_in_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_in_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_in_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_in_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_10_auto_in_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_10_auto_in_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_in_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_out_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_out_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_out_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_10_auto_out_aw_bits_addr; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_out_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_out_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_10_auto_out_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_10_auto_out_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_out_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_out_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_out_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_out_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_10_auto_out_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_out_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_out_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_out_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_10_auto_out_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_10_auto_out_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_out_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_out_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_out_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_10_auto_out_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_10_auto_out_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_out_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_11_clock; // @[Buffer.scala 58:29]
  wire  axi4buf_11_reset; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_in_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_in_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_in_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_11_auto_in_aw_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_11_auto_in_aw_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_in_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_in_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_11_auto_in_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_11_auto_in_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_in_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_in_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_in_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_in_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_11_auto_in_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_in_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_in_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_in_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_11_auto_in_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_11_auto_in_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_in_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_in_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_in_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_11_auto_in_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_11_auto_in_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_in_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_out_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_out_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_out_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_11_auto_out_aw_bits_addr; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_out_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_out_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_11_auto_out_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_11_auto_out_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_out_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_out_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_out_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_out_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_11_auto_out_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_out_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_out_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_out_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_11_auto_out_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_11_auto_out_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_out_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_out_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_out_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_11_auto_out_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_11_auto_out_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_out_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_12_clock; // @[Buffer.scala 58:29]
  wire  axi4buf_12_reset; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_in_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_in_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_in_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_12_auto_in_aw_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_12_auto_in_aw_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_in_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_in_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_12_auto_in_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_12_auto_in_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_in_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_in_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_in_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_in_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_12_auto_in_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_in_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_in_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_in_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_12_auto_in_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_12_auto_in_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_in_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_in_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_in_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_12_auto_in_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_12_auto_in_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_in_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_out_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_out_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_out_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_12_auto_out_aw_bits_addr; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_out_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_out_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_12_auto_out_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_12_auto_out_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_out_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_out_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_out_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_out_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_12_auto_out_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_out_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_out_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_out_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_12_auto_out_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_12_auto_out_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_out_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_out_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_out_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_12_auto_out_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_12_auto_out_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_out_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_13_clock; // @[Buffer.scala 58:29]
  wire  axi4buf_13_reset; // @[Buffer.scala 58:29]
  wire  axi4buf_13_auto_in_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_13_auto_in_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_13_auto_in_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_13_auto_in_aw_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_13_auto_in_aw_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_13_auto_in_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_13_auto_in_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_13_auto_in_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_13_auto_in_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_13_auto_in_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_13_auto_in_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_13_auto_in_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_13_auto_in_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_13_auto_in_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_13_auto_in_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_13_auto_in_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_13_auto_in_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_13_auto_in_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_13_auto_in_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_13_auto_in_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_13_auto_in_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_13_auto_in_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_13_auto_in_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_13_auto_in_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_13_auto_in_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_13_auto_out_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_13_auto_out_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_13_auto_out_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_13_auto_out_aw_bits_addr; // @[Buffer.scala 58:29]
  wire  axi4buf_13_auto_out_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_13_auto_out_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_13_auto_out_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_13_auto_out_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_13_auto_out_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_13_auto_out_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_13_auto_out_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_13_auto_out_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_13_auto_out_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_13_auto_out_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_13_auto_out_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_13_auto_out_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_13_auto_out_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_13_auto_out_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_13_auto_out_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_13_auto_out_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_13_auto_out_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_13_auto_out_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_13_auto_out_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_13_auto_out_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_14_clock; // @[Buffer.scala 58:29]
  wire  axi4buf_14_reset; // @[Buffer.scala 58:29]
  wire  axi4buf_14_auto_in_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_14_auto_in_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_14_auto_in_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_14_auto_in_aw_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_14_auto_in_aw_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_14_auto_in_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_14_auto_in_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_14_auto_in_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_14_auto_in_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_14_auto_in_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_14_auto_in_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_14_auto_in_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_14_auto_in_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_14_auto_in_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_14_auto_in_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_14_auto_in_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_14_auto_in_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_14_auto_in_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_14_auto_in_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_14_auto_in_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_14_auto_in_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_14_auto_in_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_14_auto_in_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_14_auto_in_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_14_auto_in_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_14_auto_out_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_14_auto_out_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_14_auto_out_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_14_auto_out_aw_bits_addr; // @[Buffer.scala 58:29]
  wire  axi4buf_14_auto_out_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_14_auto_out_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_14_auto_out_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_14_auto_out_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_14_auto_out_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_14_auto_out_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_14_auto_out_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_14_auto_out_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_14_auto_out_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_14_auto_out_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_14_auto_out_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_14_auto_out_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_14_auto_out_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_14_auto_out_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_14_auto_out_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_14_auto_out_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_14_auto_out_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_14_auto_out_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_14_auto_out_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_14_auto_out_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_15_clock; // @[Buffer.scala 58:29]
  wire  axi4buf_15_reset; // @[Buffer.scala 58:29]
  wire  axi4buf_15_auto_in_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_15_auto_in_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_15_auto_in_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_15_auto_in_aw_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_15_auto_in_aw_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_15_auto_in_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_15_auto_in_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_15_auto_in_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_15_auto_in_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_15_auto_in_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_15_auto_in_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_15_auto_in_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_15_auto_in_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_15_auto_in_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_15_auto_in_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_15_auto_in_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_15_auto_in_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_15_auto_in_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_15_auto_in_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_15_auto_in_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_15_auto_in_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_15_auto_in_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_15_auto_in_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_15_auto_in_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_15_auto_in_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_15_auto_out_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_15_auto_out_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_15_auto_out_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_15_auto_out_aw_bits_addr; // @[Buffer.scala 58:29]
  wire  axi4buf_15_auto_out_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_15_auto_out_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_15_auto_out_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_15_auto_out_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_15_auto_out_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_15_auto_out_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_15_auto_out_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_15_auto_out_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_15_auto_out_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_15_auto_out_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_15_auto_out_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_15_auto_out_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_15_auto_out_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_15_auto_out_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_15_auto_out_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_15_auto_out_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_15_auto_out_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_15_auto_out_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_15_auto_out_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_15_auto_out_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_16_clock; // @[Buffer.scala 58:29]
  wire  axi4buf_16_reset; // @[Buffer.scala 58:29]
  wire  axi4buf_16_auto_in_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_16_auto_in_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_16_auto_in_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_16_auto_in_aw_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_16_auto_in_aw_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_16_auto_in_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_16_auto_in_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_16_auto_in_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_16_auto_in_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_16_auto_in_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_16_auto_in_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_16_auto_in_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_16_auto_in_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_16_auto_in_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_16_auto_in_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_16_auto_in_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_16_auto_in_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_16_auto_in_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_16_auto_in_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_16_auto_in_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_16_auto_in_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_16_auto_in_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_16_auto_in_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_16_auto_in_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_16_auto_in_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_16_auto_out_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_16_auto_out_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_16_auto_out_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_16_auto_out_aw_bits_addr; // @[Buffer.scala 58:29]
  wire  axi4buf_16_auto_out_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_16_auto_out_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_16_auto_out_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_16_auto_out_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_16_auto_out_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_16_auto_out_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_16_auto_out_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_16_auto_out_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_16_auto_out_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_16_auto_out_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_16_auto_out_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_16_auto_out_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_16_auto_out_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_16_auto_out_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_16_auto_out_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_16_auto_out_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_16_auto_out_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_16_auto_out_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_16_auto_out_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_16_auto_out_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_17_clock; // @[Buffer.scala 58:29]
  wire  axi4buf_17_reset; // @[Buffer.scala 58:29]
  wire  axi4buf_17_auto_in_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_17_auto_in_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_17_auto_in_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_17_auto_in_aw_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_17_auto_in_aw_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_17_auto_in_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_17_auto_in_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_17_auto_in_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_17_auto_in_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_17_auto_in_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_17_auto_in_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_17_auto_in_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_17_auto_in_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_17_auto_in_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_17_auto_in_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_17_auto_in_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_17_auto_in_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_17_auto_in_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_17_auto_in_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_17_auto_in_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_17_auto_in_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_17_auto_in_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_17_auto_in_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_17_auto_in_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_17_auto_in_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_17_auto_out_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_17_auto_out_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_17_auto_out_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_17_auto_out_aw_bits_addr; // @[Buffer.scala 58:29]
  wire  axi4buf_17_auto_out_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_17_auto_out_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_17_auto_out_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_17_auto_out_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_17_auto_out_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_17_auto_out_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_17_auto_out_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_17_auto_out_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_17_auto_out_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_17_auto_out_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_17_auto_out_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_17_auto_out_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_17_auto_out_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_17_auto_out_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_17_auto_out_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_17_auto_out_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_17_auto_out_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_17_auto_out_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_17_auto_out_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_17_auto_out_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_18_clock; // @[Buffer.scala 58:29]
  wire  axi4buf_18_reset; // @[Buffer.scala 58:29]
  wire  axi4buf_18_auto_in_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_18_auto_in_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_18_auto_in_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_18_auto_in_aw_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_18_auto_in_aw_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_18_auto_in_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_18_auto_in_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_18_auto_in_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_18_auto_in_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_18_auto_in_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_18_auto_in_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_18_auto_in_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_18_auto_in_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_18_auto_in_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_18_auto_in_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_18_auto_in_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_18_auto_in_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_18_auto_in_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_18_auto_in_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_18_auto_in_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_18_auto_in_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_18_auto_in_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_18_auto_in_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_18_auto_in_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_18_auto_in_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_18_auto_out_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_18_auto_out_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_18_auto_out_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_18_auto_out_aw_bits_addr; // @[Buffer.scala 58:29]
  wire  axi4buf_18_auto_out_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_18_auto_out_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_18_auto_out_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_18_auto_out_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_18_auto_out_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_18_auto_out_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_18_auto_out_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_18_auto_out_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_18_auto_out_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_18_auto_out_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_18_auto_out_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_18_auto_out_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_18_auto_out_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_18_auto_out_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_18_auto_out_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_18_auto_out_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_18_auto_out_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_18_auto_out_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_18_auto_out_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_18_auto_out_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_19_clock; // @[Buffer.scala 58:29]
  wire  axi4buf_19_reset; // @[Buffer.scala 58:29]
  wire  axi4buf_19_auto_in_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_19_auto_in_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_19_auto_in_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_19_auto_in_aw_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_19_auto_in_aw_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_19_auto_in_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_19_auto_in_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_19_auto_in_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_19_auto_in_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_19_auto_in_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_19_auto_in_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_19_auto_in_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_19_auto_in_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_19_auto_in_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_19_auto_in_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_19_auto_in_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_19_auto_in_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_19_auto_in_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_19_auto_in_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_19_auto_in_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_19_auto_in_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_19_auto_in_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_19_auto_in_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_19_auto_in_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_19_auto_in_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_19_auto_out_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_19_auto_out_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_19_auto_out_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_19_auto_out_aw_bits_addr; // @[Buffer.scala 58:29]
  wire  axi4buf_19_auto_out_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_19_auto_out_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_19_auto_out_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_19_auto_out_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_19_auto_out_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_19_auto_out_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_19_auto_out_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_19_auto_out_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_19_auto_out_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_19_auto_out_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_19_auto_out_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_19_auto_out_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_19_auto_out_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_19_auto_out_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_19_auto_out_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_19_auto_out_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_19_auto_out_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_19_auto_out_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_19_auto_out_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_19_auto_out_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_20_clock; // @[Buffer.scala 58:29]
  wire  axi4buf_20_reset; // @[Buffer.scala 58:29]
  wire  axi4buf_20_auto_in_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_20_auto_in_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_20_auto_in_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_20_auto_in_aw_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_20_auto_in_aw_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_20_auto_in_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_20_auto_in_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_20_auto_in_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_20_auto_in_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_20_auto_in_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_20_auto_in_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_20_auto_in_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_20_auto_in_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_20_auto_in_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_20_auto_in_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_20_auto_in_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_20_auto_in_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_20_auto_in_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_20_auto_in_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_20_auto_in_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_20_auto_in_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_20_auto_in_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_20_auto_in_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_20_auto_in_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_20_auto_in_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_20_auto_out_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_20_auto_out_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_20_auto_out_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_20_auto_out_aw_bits_addr; // @[Buffer.scala 58:29]
  wire  axi4buf_20_auto_out_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_20_auto_out_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_20_auto_out_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_20_auto_out_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_20_auto_out_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_20_auto_out_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_20_auto_out_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_20_auto_out_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_20_auto_out_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_20_auto_out_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_20_auto_out_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_20_auto_out_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_20_auto_out_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_20_auto_out_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_20_auto_out_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_20_auto_out_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_20_auto_out_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_20_auto_out_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_20_auto_out_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_20_auto_out_r_bits_last; // @[Buffer.scala 58:29]
  wire  buffer_clock; // @[Buffer.scala 29:28]
  wire  buffer_reset; // @[Buffer.scala 29:28]
  wire  buffer_auto_in_ready; // @[Buffer.scala 29:28]
  wire  buffer_auto_in_valid; // @[Buffer.scala 29:28]
  wire [31:0] buffer_auto_in_bits_data; // @[Buffer.scala 29:28]
  wire  buffer_auto_in_bits_last; // @[Buffer.scala 29:28]
  wire  buffer_auto_out_ready; // @[Buffer.scala 29:28]
  wire  buffer_auto_out_valid; // @[Buffer.scala 29:28]
  wire [31:0] buffer_auto_out_bits_data; // @[Buffer.scala 29:28]
  wire  buffer_auto_out_bits_last; // @[Buffer.scala 29:28]
  wire  buffer_1_clock; // @[Buffer.scala 29:28]
  wire  buffer_1_reset; // @[Buffer.scala 29:28]
  wire  buffer_1_auto_in_ready; // @[Buffer.scala 29:28]
  wire  buffer_1_auto_in_valid; // @[Buffer.scala 29:28]
  wire [31:0] buffer_1_auto_in_bits_data; // @[Buffer.scala 29:28]
  wire  buffer_1_auto_in_bits_last; // @[Buffer.scala 29:28]
  wire  buffer_1_auto_out_ready; // @[Buffer.scala 29:28]
  wire  buffer_1_auto_out_valid; // @[Buffer.scala 29:28]
  wire [31:0] buffer_1_auto_out_bits_data; // @[Buffer.scala 29:28]
  wire  buffer_1_auto_out_bits_last; // @[Buffer.scala 29:28]
  wire  buffer_2_clock; // @[Buffer.scala 29:28]
  wire  buffer_2_reset; // @[Buffer.scala 29:28]
  wire  buffer_2_auto_in_ready; // @[Buffer.scala 29:28]
  wire  buffer_2_auto_in_valid; // @[Buffer.scala 29:28]
  wire [31:0] buffer_2_auto_in_bits_data; // @[Buffer.scala 29:28]
  wire  buffer_2_auto_in_bits_last; // @[Buffer.scala 29:28]
  wire  buffer_2_auto_out_ready; // @[Buffer.scala 29:28]
  wire  buffer_2_auto_out_valid; // @[Buffer.scala 29:28]
  wire [31:0] buffer_2_auto_out_bits_data; // @[Buffer.scala 29:28]
  wire  buffer_2_auto_out_bits_last; // @[Buffer.scala 29:28]
  wire  buffer_3_clock; // @[Buffer.scala 29:28]
  wire  buffer_3_reset; // @[Buffer.scala 29:28]
  wire  buffer_3_auto_in_ready; // @[Buffer.scala 29:28]
  wire  buffer_3_auto_in_valid; // @[Buffer.scala 29:28]
  wire [31:0] buffer_3_auto_in_bits_data; // @[Buffer.scala 29:28]
  wire  buffer_3_auto_in_bits_last; // @[Buffer.scala 29:28]
  wire  buffer_3_auto_out_ready; // @[Buffer.scala 29:28]
  wire  buffer_3_auto_out_valid; // @[Buffer.scala 29:28]
  wire [31:0] buffer_3_auto_out_bits_data; // @[Buffer.scala 29:28]
  wire  buffer_3_auto_out_bits_last; // @[Buffer.scala 29:28]
  wire  buffer_4_clock; // @[Buffer.scala 29:28]
  wire  buffer_4_reset; // @[Buffer.scala 29:28]
  wire  buffer_4_auto_in_ready; // @[Buffer.scala 29:28]
  wire  buffer_4_auto_in_valid; // @[Buffer.scala 29:28]
  wire [31:0] buffer_4_auto_in_bits_data; // @[Buffer.scala 29:28]
  wire  buffer_4_auto_in_bits_last; // @[Buffer.scala 29:28]
  wire  buffer_4_auto_out_ready; // @[Buffer.scala 29:28]
  wire  buffer_4_auto_out_valid; // @[Buffer.scala 29:28]
  wire [31:0] buffer_4_auto_out_bits_data; // @[Buffer.scala 29:28]
  wire  buffer_4_auto_out_bits_last; // @[Buffer.scala 29:28]
  wire  buffer_5_clock; // @[Buffer.scala 29:28]
  wire  buffer_5_reset; // @[Buffer.scala 29:28]
  wire  buffer_5_auto_in_ready; // @[Buffer.scala 29:28]
  wire  buffer_5_auto_in_valid; // @[Buffer.scala 29:28]
  wire [31:0] buffer_5_auto_in_bits_data; // @[Buffer.scala 29:28]
  wire  buffer_5_auto_in_bits_last; // @[Buffer.scala 29:28]
  wire  buffer_5_auto_out_ready; // @[Buffer.scala 29:28]
  wire  buffer_5_auto_out_valid; // @[Buffer.scala 29:28]
  wire [31:0] buffer_5_auto_out_bits_data; // @[Buffer.scala 29:28]
  wire  buffer_5_auto_out_bits_last; // @[Buffer.scala 29:28]
  wire  buffer_6_clock; // @[Buffer.scala 29:28]
  wire  buffer_6_reset; // @[Buffer.scala 29:28]
  wire  buffer_6_auto_in_ready; // @[Buffer.scala 29:28]
  wire  buffer_6_auto_in_valid; // @[Buffer.scala 29:28]
  wire [31:0] buffer_6_auto_in_bits_data; // @[Buffer.scala 29:28]
  wire  buffer_6_auto_in_bits_last; // @[Buffer.scala 29:28]
  wire  buffer_6_auto_out_ready; // @[Buffer.scala 29:28]
  wire  buffer_6_auto_out_valid; // @[Buffer.scala 29:28]
  wire [31:0] buffer_6_auto_out_bits_data; // @[Buffer.scala 29:28]
  wire  buffer_6_auto_out_bits_last; // @[Buffer.scala 29:28]
  wire  buffer_7_clock; // @[Buffer.scala 29:28]
  wire  buffer_7_reset; // @[Buffer.scala 29:28]
  wire  buffer_7_auto_in_ready; // @[Buffer.scala 29:28]
  wire  buffer_7_auto_in_valid; // @[Buffer.scala 29:28]
  wire [31:0] buffer_7_auto_in_bits_data; // @[Buffer.scala 29:28]
  wire  buffer_7_auto_in_bits_last; // @[Buffer.scala 29:28]
  wire  buffer_7_auto_out_ready; // @[Buffer.scala 29:28]
  wire  buffer_7_auto_out_valid; // @[Buffer.scala 29:28]
  wire [31:0] buffer_7_auto_out_bits_data; // @[Buffer.scala 29:28]
  wire  buffer_7_auto_out_bits_last; // @[Buffer.scala 29:28]
  wire  buffer_8_clock; // @[Buffer.scala 29:28]
  wire  buffer_8_reset; // @[Buffer.scala 29:28]
  wire  buffer_8_auto_in_ready; // @[Buffer.scala 29:28]
  wire  buffer_8_auto_in_valid; // @[Buffer.scala 29:28]
  wire [31:0] buffer_8_auto_in_bits_data; // @[Buffer.scala 29:28]
  wire  buffer_8_auto_in_bits_last; // @[Buffer.scala 29:28]
  wire  buffer_8_auto_out_ready; // @[Buffer.scala 29:28]
  wire  buffer_8_auto_out_valid; // @[Buffer.scala 29:28]
  wire [31:0] buffer_8_auto_out_bits_data; // @[Buffer.scala 29:28]
  wire  buffer_8_auto_out_bits_last; // @[Buffer.scala 29:28]
  wire  buffer_9_clock; // @[Buffer.scala 29:28]
  wire  buffer_9_reset; // @[Buffer.scala 29:28]
  wire  buffer_9_auto_in_ready; // @[Buffer.scala 29:28]
  wire  buffer_9_auto_in_valid; // @[Buffer.scala 29:28]
  wire [31:0] buffer_9_auto_in_bits_data; // @[Buffer.scala 29:28]
  wire  buffer_9_auto_in_bits_last; // @[Buffer.scala 29:28]
  wire  buffer_9_auto_out_ready; // @[Buffer.scala 29:28]
  wire  buffer_9_auto_out_valid; // @[Buffer.scala 29:28]
  wire [31:0] buffer_9_auto_out_bits_data; // @[Buffer.scala 29:28]
  wire  buffer_9_auto_out_bits_last; // @[Buffer.scala 29:28]
  wire  converter_auto_in_aw_ready; // @[Node.scala 65:31]
  wire  converter_auto_in_aw_valid; // @[Node.scala 65:31]
  wire  converter_auto_in_aw_bits_id; // @[Node.scala 65:31]
  wire [31:0] converter_auto_in_aw_bits_addr; // @[Node.scala 65:31]
  wire [2:0] converter_auto_in_aw_bits_size; // @[Node.scala 65:31]
  wire  converter_auto_in_w_ready; // @[Node.scala 65:31]
  wire  converter_auto_in_w_valid; // @[Node.scala 65:31]
  wire [31:0] converter_auto_in_w_bits_data; // @[Node.scala 65:31]
  wire [3:0] converter_auto_in_w_bits_strb; // @[Node.scala 65:31]
  wire  converter_auto_in_w_bits_last; // @[Node.scala 65:31]
  wire  converter_auto_in_b_ready; // @[Node.scala 65:31]
  wire  converter_auto_in_b_valid; // @[Node.scala 65:31]
  wire [1:0] converter_auto_in_b_bits_resp; // @[Node.scala 65:31]
  wire  converter_auto_in_ar_ready; // @[Node.scala 65:31]
  wire  converter_auto_in_ar_valid; // @[Node.scala 65:31]
  wire  converter_auto_in_ar_bits_id; // @[Node.scala 65:31]
  wire [31:0] converter_auto_in_ar_bits_addr; // @[Node.scala 65:31]
  wire [2:0] converter_auto_in_ar_bits_size; // @[Node.scala 65:31]
  wire  converter_auto_in_r_ready; // @[Node.scala 65:31]
  wire  converter_auto_in_r_valid; // @[Node.scala 65:31]
  wire [31:0] converter_auto_in_r_bits_data; // @[Node.scala 65:31]
  wire [1:0] converter_auto_in_r_bits_resp; // @[Node.scala 65:31]
  wire  converter_auto_in_r_bits_last; // @[Node.scala 65:31]
  wire  converter_auto_out_aw_ready; // @[Node.scala 65:31]
  wire  converter_auto_out_aw_valid; // @[Node.scala 65:31]
  wire  converter_auto_out_aw_bits_id; // @[Node.scala 65:31]
  wire [29:0] converter_auto_out_aw_bits_addr; // @[Node.scala 65:31]
  wire [2:0] converter_auto_out_aw_bits_size; // @[Node.scala 65:31]
  wire  converter_auto_out_w_ready; // @[Node.scala 65:31]
  wire  converter_auto_out_w_valid; // @[Node.scala 65:31]
  wire [31:0] converter_auto_out_w_bits_data; // @[Node.scala 65:31]
  wire [3:0] converter_auto_out_w_bits_strb; // @[Node.scala 65:31]
  wire  converter_auto_out_w_bits_last; // @[Node.scala 65:31]
  wire  converter_auto_out_b_ready; // @[Node.scala 65:31]
  wire  converter_auto_out_b_valid; // @[Node.scala 65:31]
  wire [1:0] converter_auto_out_b_bits_resp; // @[Node.scala 65:31]
  wire  converter_auto_out_ar_ready; // @[Node.scala 65:31]
  wire  converter_auto_out_ar_valid; // @[Node.scala 65:31]
  wire  converter_auto_out_ar_bits_id; // @[Node.scala 65:31]
  wire [29:0] converter_auto_out_ar_bits_addr; // @[Node.scala 65:31]
  wire [2:0] converter_auto_out_ar_bits_size; // @[Node.scala 65:31]
  wire  converter_auto_out_r_ready; // @[Node.scala 65:31]
  wire  converter_auto_out_r_valid; // @[Node.scala 65:31]
  wire [31:0] converter_auto_out_r_bits_data; // @[Node.scala 65:31]
  wire [1:0] converter_auto_out_r_bits_resp; // @[Node.scala 65:31]
  wire  converter_auto_out_r_bits_last; // @[Node.scala 65:31]
  wire  converter_1_auto_in_ready; // @[Nodes.scala 165:31]
  wire  converter_1_auto_in_valid; // @[Nodes.scala 165:31]
  wire [7:0] converter_1_auto_in_bits_data; // @[Nodes.scala 165:31]
  wire  converter_1_auto_in_bits_last; // @[Nodes.scala 165:31]
  wire  converter_1_auto_out_ready; // @[Nodes.scala 165:31]
  wire  converter_1_auto_out_valid; // @[Nodes.scala 165:31]
  wire [7:0] converter_1_auto_out_bits_data; // @[Nodes.scala 165:31]
  wire  converter_1_auto_out_bits_last; // @[Nodes.scala 165:31]
  wire  converter_2_auto_in_ready; // @[Nodes.scala 201:31]
  wire  converter_2_auto_in_valid; // @[Nodes.scala 201:31]
  wire [7:0] converter_2_auto_in_bits_data; // @[Nodes.scala 201:31]
  wire  converter_2_auto_in_bits_last; // @[Nodes.scala 201:31]
  wire  converter_2_auto_out_ready; // @[Nodes.scala 201:31]
  wire  converter_2_auto_out_valid; // @[Nodes.scala 201:31]
  wire [7:0] converter_2_auto_out_bits_data; // @[Nodes.scala 201:31]
  wire  converter_2_auto_out_bits_last; // @[Nodes.scala 201:31]
  AXI4StreamWidthAdapater_4_to_1 widthAdapter ( // @[AXI4StreamWidthAdapter.scala 82:34]
    .clock(widthAdapter_clock),
    .reset(widthAdapter_reset),
    .auto_in_ready(widthAdapter_auto_in_ready),
    .auto_in_valid(widthAdapter_auto_in_valid),
    .auto_in_bits_data(widthAdapter_auto_in_bits_data),
    .auto_in_bits_last(widthAdapter_auto_in_bits_last),
    .auto_out_ready(widthAdapter_auto_out_ready),
    .auto_out_valid(widthAdapter_auto_out_valid),
    .auto_out_bits_data(widthAdapter_auto_out_bits_data),
    .auto_out_bits_last(widthAdapter_auto_out_bits_last)
  );
  AXI4Splitter in_split ( // @[SpectrometerTestWithoutLA.scala 59:29]
    .clock(in_split_clock),
    .reset(in_split_reset),
    .auto_mem_in_aw_ready(in_split_auto_mem_in_aw_ready),
    .auto_mem_in_aw_valid(in_split_auto_mem_in_aw_valid),
    .auto_mem_in_aw_bits_id(in_split_auto_mem_in_aw_bits_id),
    .auto_mem_in_aw_bits_addr(in_split_auto_mem_in_aw_bits_addr),
    .auto_mem_in_w_ready(in_split_auto_mem_in_w_ready),
    .auto_mem_in_w_valid(in_split_auto_mem_in_w_valid),
    .auto_mem_in_w_bits_data(in_split_auto_mem_in_w_bits_data),
    .auto_mem_in_w_bits_strb(in_split_auto_mem_in_w_bits_strb),
    .auto_mem_in_b_ready(in_split_auto_mem_in_b_ready),
    .auto_mem_in_b_valid(in_split_auto_mem_in_b_valid),
    .auto_mem_in_b_bits_id(in_split_auto_mem_in_b_bits_id),
    .auto_mem_in_ar_ready(in_split_auto_mem_in_ar_ready),
    .auto_mem_in_ar_valid(in_split_auto_mem_in_ar_valid),
    .auto_mem_in_ar_bits_id(in_split_auto_mem_in_ar_bits_id),
    .auto_mem_in_ar_bits_addr(in_split_auto_mem_in_ar_bits_addr),
    .auto_mem_in_ar_bits_size(in_split_auto_mem_in_ar_bits_size),
    .auto_mem_in_r_ready(in_split_auto_mem_in_r_ready),
    .auto_mem_in_r_valid(in_split_auto_mem_in_r_valid),
    .auto_mem_in_r_bits_id(in_split_auto_mem_in_r_bits_id),
    .auto_mem_in_r_bits_data(in_split_auto_mem_in_r_bits_data),
    .auto_stream_in_ready(in_split_auto_stream_in_ready),
    .auto_stream_in_valid(in_split_auto_stream_in_valid),
    .auto_stream_in_bits_data(in_split_auto_stream_in_bits_data),
    .auto_stream_in_bits_last(in_split_auto_stream_in_bits_last),
    .auto_stream_out_4_ready(in_split_auto_stream_out_4_ready),
    .auto_stream_out_4_valid(in_split_auto_stream_out_4_valid),
    .auto_stream_out_4_bits_data(in_split_auto_stream_out_4_bits_data),
    .auto_stream_out_4_bits_last(in_split_auto_stream_out_4_bits_last),
    .auto_stream_out_3_ready(in_split_auto_stream_out_3_ready),
    .auto_stream_out_3_valid(in_split_auto_stream_out_3_valid),
    .auto_stream_out_3_bits_data(in_split_auto_stream_out_3_bits_data),
    .auto_stream_out_3_bits_last(in_split_auto_stream_out_3_bits_last),
    .auto_stream_out_2_ready(in_split_auto_stream_out_2_ready),
    .auto_stream_out_2_valid(in_split_auto_stream_out_2_valid),
    .auto_stream_out_2_bits_data(in_split_auto_stream_out_2_bits_data),
    .auto_stream_out_2_bits_last(in_split_auto_stream_out_2_bits_last),
    .auto_stream_out_1_ready(in_split_auto_stream_out_1_ready),
    .auto_stream_out_1_valid(in_split_auto_stream_out_1_valid),
    .auto_stream_out_1_bits_data(in_split_auto_stream_out_1_bits_data),
    .auto_stream_out_1_bits_last(in_split_auto_stream_out_1_bits_last),
    .auto_stream_out_0_ready(in_split_auto_stream_out_0_ready),
    .auto_stream_out_0_valid(in_split_auto_stream_out_0_valid),
    .auto_stream_out_0_bits_data(in_split_auto_stream_out_0_bits_data),
    .auto_stream_out_0_bits_last(in_split_auto_stream_out_0_bits_last)
  );
  StreamBuffer in_queue ( // @[SpectrometerTestWithoutLA.scala 60:29]
    .clock(in_queue_clock),
    .reset(in_queue_reset),
    .auto_out_out_ready(in_queue_auto_out_out_ready),
    .auto_out_out_valid(in_queue_auto_out_out_valid),
    .auto_out_out_bits_data(in_queue_auto_out_out_bits_data),
    .auto_out_out_bits_last(in_queue_auto_out_out_bits_last),
    .auto_in_in_ready(in_queue_auto_in_in_ready),
    .auto_in_in_valid(in_queue_auto_in_in_valid),
    .auto_in_in_bits_data(in_queue_auto_in_in_bits_data),
    .auto_in_in_bits_last(in_queue_auto_in_in_bits_last)
  );
  PLFGDspBlockMem plfg ( // @[SpectrometerTestWithoutLA.scala 62:30]
    .clock(plfg_clock),
    .reset(plfg_reset),
    .auto_mem_in_aw_ready(plfg_auto_mem_in_aw_ready),
    .auto_mem_in_aw_valid(plfg_auto_mem_in_aw_valid),
    .auto_mem_in_aw_bits_id(plfg_auto_mem_in_aw_bits_id),
    .auto_mem_in_aw_bits_addr(plfg_auto_mem_in_aw_bits_addr),
    .auto_mem_in_w_ready(plfg_auto_mem_in_w_ready),
    .auto_mem_in_w_valid(plfg_auto_mem_in_w_valid),
    .auto_mem_in_w_bits_data(plfg_auto_mem_in_w_bits_data),
    .auto_mem_in_w_bits_strb(plfg_auto_mem_in_w_bits_strb),
    .auto_mem_in_w_bits_last(plfg_auto_mem_in_w_bits_last),
    .auto_mem_in_b_ready(plfg_auto_mem_in_b_ready),
    .auto_mem_in_b_valid(plfg_auto_mem_in_b_valid),
    .auto_mem_in_b_bits_resp(plfg_auto_mem_in_b_bits_resp),
    .auto_mem_in_ar_ready(plfg_auto_mem_in_ar_ready),
    .auto_mem_in_ar_valid(plfg_auto_mem_in_ar_valid),
    .auto_mem_in_ar_bits_id(plfg_auto_mem_in_ar_bits_id),
    .auto_mem_in_ar_bits_addr(plfg_auto_mem_in_ar_bits_addr),
    .auto_mem_in_ar_bits_size(plfg_auto_mem_in_ar_bits_size),
    .auto_mem_in_r_ready(plfg_auto_mem_in_r_ready),
    .auto_mem_in_r_valid(plfg_auto_mem_in_r_valid),
    .auto_mem_in_r_bits_data(plfg_auto_mem_in_r_bits_data),
    .auto_mem_in_r_bits_resp(plfg_auto_mem_in_r_bits_resp),
    .auto_mem_in_r_bits_last(plfg_auto_mem_in_r_bits_last),
    .auto_stream_out_ready(plfg_auto_stream_out_ready),
    .auto_stream_out_valid(plfg_auto_stream_out_valid),
    .auto_stream_out_bits_data(plfg_auto_stream_out_bits_data),
    .auto_stream_out_bits_last(plfg_auto_stream_out_bits_last)
  );
  AXI4Splitter_1 plfg_split ( // @[SpectrometerTestWithoutLA.scala 63:30]
    .clock(plfg_split_clock),
    .reset(plfg_split_reset),
    .auto_mem_in_aw_ready(plfg_split_auto_mem_in_aw_ready),
    .auto_mem_in_aw_valid(plfg_split_auto_mem_in_aw_valid),
    .auto_mem_in_aw_bits_id(plfg_split_auto_mem_in_aw_bits_id),
    .auto_mem_in_aw_bits_addr(plfg_split_auto_mem_in_aw_bits_addr),
    .auto_mem_in_w_ready(plfg_split_auto_mem_in_w_ready),
    .auto_mem_in_w_valid(plfg_split_auto_mem_in_w_valid),
    .auto_mem_in_w_bits_data(plfg_split_auto_mem_in_w_bits_data),
    .auto_mem_in_w_bits_strb(plfg_split_auto_mem_in_w_bits_strb),
    .auto_mem_in_b_ready(plfg_split_auto_mem_in_b_ready),
    .auto_mem_in_b_valid(plfg_split_auto_mem_in_b_valid),
    .auto_mem_in_b_bits_id(plfg_split_auto_mem_in_b_bits_id),
    .auto_mem_in_ar_ready(plfg_split_auto_mem_in_ar_ready),
    .auto_mem_in_ar_valid(plfg_split_auto_mem_in_ar_valid),
    .auto_mem_in_ar_bits_id(plfg_split_auto_mem_in_ar_bits_id),
    .auto_mem_in_ar_bits_addr(plfg_split_auto_mem_in_ar_bits_addr),
    .auto_mem_in_ar_bits_size(plfg_split_auto_mem_in_ar_bits_size),
    .auto_mem_in_r_ready(plfg_split_auto_mem_in_r_ready),
    .auto_mem_in_r_valid(plfg_split_auto_mem_in_r_valid),
    .auto_mem_in_r_bits_id(plfg_split_auto_mem_in_r_bits_id),
    .auto_mem_in_r_bits_data(plfg_split_auto_mem_in_r_bits_data),
    .auto_stream_in_ready(plfg_split_auto_stream_in_ready),
    .auto_stream_in_valid(plfg_split_auto_stream_in_valid),
    .auto_stream_in_bits_data(plfg_split_auto_stream_in_bits_data),
    .auto_stream_in_bits_last(plfg_split_auto_stream_in_bits_last),
    .auto_stream_out_1_ready(plfg_split_auto_stream_out_1_ready),
    .auto_stream_out_1_valid(plfg_split_auto_stream_out_1_valid),
    .auto_stream_out_1_bits_data(plfg_split_auto_stream_out_1_bits_data),
    .auto_stream_out_1_bits_last(plfg_split_auto_stream_out_1_bits_last),
    .auto_stream_out_0_ready(plfg_split_auto_stream_out_0_ready),
    .auto_stream_out_0_valid(plfg_split_auto_stream_out_0_valid),
    .auto_stream_out_0_bits_data(plfg_split_auto_stream_out_0_bits_data),
    .auto_stream_out_0_bits_last(plfg_split_auto_stream_out_0_bits_last)
  );
  AXI4StreamMux plfg_mux_0 ( // @[SpectrometerTestWithoutLA.scala 64:30]
    .clock(plfg_mux_0_clock),
    .reset(plfg_mux_0_reset),
    .auto_register_in_aw_ready(plfg_mux_0_auto_register_in_aw_ready),
    .auto_register_in_aw_valid(plfg_mux_0_auto_register_in_aw_valid),
    .auto_register_in_aw_bits_id(plfg_mux_0_auto_register_in_aw_bits_id),
    .auto_register_in_aw_bits_addr(plfg_mux_0_auto_register_in_aw_bits_addr),
    .auto_register_in_w_ready(plfg_mux_0_auto_register_in_w_ready),
    .auto_register_in_w_valid(plfg_mux_0_auto_register_in_w_valid),
    .auto_register_in_w_bits_data(plfg_mux_0_auto_register_in_w_bits_data),
    .auto_register_in_w_bits_strb(plfg_mux_0_auto_register_in_w_bits_strb),
    .auto_register_in_b_ready(plfg_mux_0_auto_register_in_b_ready),
    .auto_register_in_b_valid(plfg_mux_0_auto_register_in_b_valid),
    .auto_register_in_b_bits_id(plfg_mux_0_auto_register_in_b_bits_id),
    .auto_register_in_ar_ready(plfg_mux_0_auto_register_in_ar_ready),
    .auto_register_in_ar_valid(plfg_mux_0_auto_register_in_ar_valid),
    .auto_register_in_ar_bits_id(plfg_mux_0_auto_register_in_ar_bits_id),
    .auto_register_in_ar_bits_addr(plfg_mux_0_auto_register_in_ar_bits_addr),
    .auto_register_in_ar_bits_size(plfg_mux_0_auto_register_in_ar_bits_size),
    .auto_register_in_r_ready(plfg_mux_0_auto_register_in_r_ready),
    .auto_register_in_r_valid(plfg_mux_0_auto_register_in_r_valid),
    .auto_register_in_r_bits_id(plfg_mux_0_auto_register_in_r_bits_id),
    .auto_register_in_r_bits_data(plfg_mux_0_auto_register_in_r_bits_data),
    .auto_stream_in_2_ready(plfg_mux_0_auto_stream_in_2_ready),
    .auto_stream_in_2_valid(plfg_mux_0_auto_stream_in_2_valid),
    .auto_stream_in_2_bits_data(plfg_mux_0_auto_stream_in_2_bits_data),
    .auto_stream_in_2_bits_last(plfg_mux_0_auto_stream_in_2_bits_last),
    .auto_stream_in_1_ready(plfg_mux_0_auto_stream_in_1_ready),
    .auto_stream_in_1_valid(plfg_mux_0_auto_stream_in_1_valid),
    .auto_stream_in_1_bits_data(plfg_mux_0_auto_stream_in_1_bits_data),
    .auto_stream_in_1_bits_last(plfg_mux_0_auto_stream_in_1_bits_last),
    .auto_stream_in_0_ready(plfg_mux_0_auto_stream_in_0_ready),
    .auto_stream_in_0_valid(plfg_mux_0_auto_stream_in_0_valid),
    .auto_stream_in_0_bits_data(plfg_mux_0_auto_stream_in_0_bits_data),
    .auto_stream_in_0_bits_last(plfg_mux_0_auto_stream_in_0_bits_last),
    .auto_stream_out_0_ready(plfg_mux_0_auto_stream_out_0_ready),
    .auto_stream_out_0_valid(plfg_mux_0_auto_stream_out_0_valid),
    .auto_stream_out_0_bits_data(plfg_mux_0_auto_stream_out_0_bits_data),
    .auto_stream_out_0_bits_last(plfg_mux_0_auto_stream_out_0_bits_last)
  );
  AXI4StreamMux_1 plfg_mux_1 ( // @[SpectrometerTestWithoutLA.scala 65:30]
    .clock(plfg_mux_1_clock),
    .reset(plfg_mux_1_reset),
    .auto_register_in_aw_ready(plfg_mux_1_auto_register_in_aw_ready),
    .auto_register_in_aw_valid(plfg_mux_1_auto_register_in_aw_valid),
    .auto_register_in_aw_bits_id(plfg_mux_1_auto_register_in_aw_bits_id),
    .auto_register_in_aw_bits_addr(plfg_mux_1_auto_register_in_aw_bits_addr),
    .auto_register_in_w_ready(plfg_mux_1_auto_register_in_w_ready),
    .auto_register_in_w_valid(plfg_mux_1_auto_register_in_w_valid),
    .auto_register_in_w_bits_data(plfg_mux_1_auto_register_in_w_bits_data),
    .auto_register_in_w_bits_strb(plfg_mux_1_auto_register_in_w_bits_strb),
    .auto_register_in_b_ready(plfg_mux_1_auto_register_in_b_ready),
    .auto_register_in_b_valid(plfg_mux_1_auto_register_in_b_valid),
    .auto_register_in_b_bits_id(plfg_mux_1_auto_register_in_b_bits_id),
    .auto_register_in_ar_ready(plfg_mux_1_auto_register_in_ar_ready),
    .auto_register_in_ar_valid(plfg_mux_1_auto_register_in_ar_valid),
    .auto_register_in_ar_bits_id(plfg_mux_1_auto_register_in_ar_bits_id),
    .auto_register_in_ar_bits_addr(plfg_mux_1_auto_register_in_ar_bits_addr),
    .auto_register_in_ar_bits_size(plfg_mux_1_auto_register_in_ar_bits_size),
    .auto_register_in_r_ready(plfg_mux_1_auto_register_in_r_ready),
    .auto_register_in_r_valid(plfg_mux_1_auto_register_in_r_valid),
    .auto_register_in_r_bits_id(plfg_mux_1_auto_register_in_r_bits_id),
    .auto_register_in_r_bits_data(plfg_mux_1_auto_register_in_r_bits_data),
    .auto_stream_in_ready(plfg_mux_1_auto_stream_in_ready),
    .auto_stream_in_valid(plfg_mux_1_auto_stream_in_valid),
    .auto_stream_in_bits_data(plfg_mux_1_auto_stream_in_bits_data),
    .auto_stream_in_bits_last(plfg_mux_1_auto_stream_in_bits_last),
    .auto_stream_out_1_ready(plfg_mux_1_auto_stream_out_1_ready),
    .auto_stream_out_1_valid(plfg_mux_1_auto_stream_out_1_valid),
    .auto_stream_out_1_bits_data(plfg_mux_1_auto_stream_out_1_bits_data),
    .auto_stream_out_1_bits_last(plfg_mux_1_auto_stream_out_1_bits_last)
  );
  AXI4NCOLazyModuleBlock nco ( // @[SpectrometerTestWithoutLA.scala 71:29]
    .clock(nco_clock),
    .reset(nco_reset),
    .auto_stream_out_ready(nco_auto_stream_out_ready),
    .auto_stream_out_valid(nco_auto_stream_out_valid),
    .auto_stream_out_bits_data(nco_auto_stream_out_bits_data),
    .auto_stream_out_bits_last(nco_auto_stream_out_bits_last),
    .auto_freq_in_ready(nco_auto_freq_in_ready),
    .auto_freq_in_valid(nco_auto_freq_in_valid),
    .auto_freq_in_bits_data(nco_auto_freq_in_bits_data),
    .auto_freq_in_bits_last(nco_auto_freq_in_bits_last)
  );
  AXI4Splitter_2 nco_split ( // @[SpectrometerTestWithoutLA.scala 72:29]
    .clock(nco_split_clock),
    .reset(nco_split_reset),
    .auto_mem_in_aw_ready(nco_split_auto_mem_in_aw_ready),
    .auto_mem_in_aw_valid(nco_split_auto_mem_in_aw_valid),
    .auto_mem_in_aw_bits_id(nco_split_auto_mem_in_aw_bits_id),
    .auto_mem_in_aw_bits_addr(nco_split_auto_mem_in_aw_bits_addr),
    .auto_mem_in_w_ready(nco_split_auto_mem_in_w_ready),
    .auto_mem_in_w_valid(nco_split_auto_mem_in_w_valid),
    .auto_mem_in_w_bits_data(nco_split_auto_mem_in_w_bits_data),
    .auto_mem_in_w_bits_strb(nco_split_auto_mem_in_w_bits_strb),
    .auto_mem_in_b_ready(nco_split_auto_mem_in_b_ready),
    .auto_mem_in_b_valid(nco_split_auto_mem_in_b_valid),
    .auto_mem_in_b_bits_id(nco_split_auto_mem_in_b_bits_id),
    .auto_mem_in_ar_ready(nco_split_auto_mem_in_ar_ready),
    .auto_mem_in_ar_valid(nco_split_auto_mem_in_ar_valid),
    .auto_mem_in_ar_bits_id(nco_split_auto_mem_in_ar_bits_id),
    .auto_mem_in_ar_bits_addr(nco_split_auto_mem_in_ar_bits_addr),
    .auto_mem_in_ar_bits_size(nco_split_auto_mem_in_ar_bits_size),
    .auto_mem_in_r_ready(nco_split_auto_mem_in_r_ready),
    .auto_mem_in_r_valid(nco_split_auto_mem_in_r_valid),
    .auto_mem_in_r_bits_id(nco_split_auto_mem_in_r_bits_id),
    .auto_mem_in_r_bits_data(nco_split_auto_mem_in_r_bits_data),
    .auto_stream_in_ready(nco_split_auto_stream_in_ready),
    .auto_stream_in_valid(nco_split_auto_stream_in_valid),
    .auto_stream_in_bits_data(nco_split_auto_stream_in_bits_data),
    .auto_stream_in_bits_last(nco_split_auto_stream_in_bits_last),
    .auto_stream_out_1_ready(nco_split_auto_stream_out_1_ready),
    .auto_stream_out_1_valid(nco_split_auto_stream_out_1_valid),
    .auto_stream_out_1_bits_data(nco_split_auto_stream_out_1_bits_data),
    .auto_stream_out_1_bits_last(nco_split_auto_stream_out_1_bits_last),
    .auto_stream_out_0_ready(nco_split_auto_stream_out_0_ready),
    .auto_stream_out_0_valid(nco_split_auto_stream_out_0_valid),
    .auto_stream_out_0_bits_data(nco_split_auto_stream_out_0_bits_data),
    .auto_stream_out_0_bits_last(nco_split_auto_stream_out_0_bits_last)
  );
  AXI4StreamMux_2 nco_mux_0 ( // @[SpectrometerTestWithoutLA.scala 73:29]
    .clock(nco_mux_0_clock),
    .reset(nco_mux_0_reset),
    .auto_register_in_aw_ready(nco_mux_0_auto_register_in_aw_ready),
    .auto_register_in_aw_valid(nco_mux_0_auto_register_in_aw_valid),
    .auto_register_in_aw_bits_id(nco_mux_0_auto_register_in_aw_bits_id),
    .auto_register_in_aw_bits_addr(nco_mux_0_auto_register_in_aw_bits_addr),
    .auto_register_in_w_ready(nco_mux_0_auto_register_in_w_ready),
    .auto_register_in_w_valid(nco_mux_0_auto_register_in_w_valid),
    .auto_register_in_w_bits_data(nco_mux_0_auto_register_in_w_bits_data),
    .auto_register_in_w_bits_strb(nco_mux_0_auto_register_in_w_bits_strb),
    .auto_register_in_b_ready(nco_mux_0_auto_register_in_b_ready),
    .auto_register_in_b_valid(nco_mux_0_auto_register_in_b_valid),
    .auto_register_in_b_bits_id(nco_mux_0_auto_register_in_b_bits_id),
    .auto_register_in_ar_ready(nco_mux_0_auto_register_in_ar_ready),
    .auto_register_in_ar_valid(nco_mux_0_auto_register_in_ar_valid),
    .auto_register_in_ar_bits_id(nco_mux_0_auto_register_in_ar_bits_id),
    .auto_register_in_ar_bits_addr(nco_mux_0_auto_register_in_ar_bits_addr),
    .auto_register_in_ar_bits_size(nco_mux_0_auto_register_in_ar_bits_size),
    .auto_register_in_r_ready(nco_mux_0_auto_register_in_r_ready),
    .auto_register_in_r_valid(nco_mux_0_auto_register_in_r_valid),
    .auto_register_in_r_bits_id(nco_mux_0_auto_register_in_r_bits_id),
    .auto_register_in_r_bits_data(nco_mux_0_auto_register_in_r_bits_data),
    .auto_stream_in_2_ready(nco_mux_0_auto_stream_in_2_ready),
    .auto_stream_in_2_valid(nco_mux_0_auto_stream_in_2_valid),
    .auto_stream_in_2_bits_data(nco_mux_0_auto_stream_in_2_bits_data),
    .auto_stream_in_2_bits_last(nco_mux_0_auto_stream_in_2_bits_last),
    .auto_stream_in_1_ready(nco_mux_0_auto_stream_in_1_ready),
    .auto_stream_in_1_valid(nco_mux_0_auto_stream_in_1_valid),
    .auto_stream_in_1_bits_data(nco_mux_0_auto_stream_in_1_bits_data),
    .auto_stream_in_1_bits_last(nco_mux_0_auto_stream_in_1_bits_last),
    .auto_stream_in_0_ready(nco_mux_0_auto_stream_in_0_ready),
    .auto_stream_in_0_valid(nco_mux_0_auto_stream_in_0_valid),
    .auto_stream_in_0_bits_data(nco_mux_0_auto_stream_in_0_bits_data),
    .auto_stream_in_0_bits_last(nco_mux_0_auto_stream_in_0_bits_last),
    .auto_stream_out_0_ready(nco_mux_0_auto_stream_out_0_ready),
    .auto_stream_out_0_valid(nco_mux_0_auto_stream_out_0_valid),
    .auto_stream_out_0_bits_data(nco_mux_0_auto_stream_out_0_bits_data),
    .auto_stream_out_0_bits_last(nco_mux_0_auto_stream_out_0_bits_last)
  );
  AXI4StreamMux_1 nco_mux_1 ( // @[SpectrometerTestWithoutLA.scala 74:29]
    .clock(nco_mux_1_clock),
    .reset(nco_mux_1_reset),
    .auto_register_in_aw_ready(nco_mux_1_auto_register_in_aw_ready),
    .auto_register_in_aw_valid(nco_mux_1_auto_register_in_aw_valid),
    .auto_register_in_aw_bits_id(nco_mux_1_auto_register_in_aw_bits_id),
    .auto_register_in_aw_bits_addr(nco_mux_1_auto_register_in_aw_bits_addr),
    .auto_register_in_w_ready(nco_mux_1_auto_register_in_w_ready),
    .auto_register_in_w_valid(nco_mux_1_auto_register_in_w_valid),
    .auto_register_in_w_bits_data(nco_mux_1_auto_register_in_w_bits_data),
    .auto_register_in_w_bits_strb(nco_mux_1_auto_register_in_w_bits_strb),
    .auto_register_in_b_ready(nco_mux_1_auto_register_in_b_ready),
    .auto_register_in_b_valid(nco_mux_1_auto_register_in_b_valid),
    .auto_register_in_b_bits_id(nco_mux_1_auto_register_in_b_bits_id),
    .auto_register_in_ar_ready(nco_mux_1_auto_register_in_ar_ready),
    .auto_register_in_ar_valid(nco_mux_1_auto_register_in_ar_valid),
    .auto_register_in_ar_bits_id(nco_mux_1_auto_register_in_ar_bits_id),
    .auto_register_in_ar_bits_addr(nco_mux_1_auto_register_in_ar_bits_addr),
    .auto_register_in_ar_bits_size(nco_mux_1_auto_register_in_ar_bits_size),
    .auto_register_in_r_ready(nco_mux_1_auto_register_in_r_ready),
    .auto_register_in_r_valid(nco_mux_1_auto_register_in_r_valid),
    .auto_register_in_r_bits_id(nco_mux_1_auto_register_in_r_bits_id),
    .auto_register_in_r_bits_data(nco_mux_1_auto_register_in_r_bits_data),
    .auto_stream_in_ready(nco_mux_1_auto_stream_in_ready),
    .auto_stream_in_valid(nco_mux_1_auto_stream_in_valid),
    .auto_stream_in_bits_data(nco_mux_1_auto_stream_in_bits_data),
    .auto_stream_in_bits_last(nco_mux_1_auto_stream_in_bits_last),
    .auto_stream_out_1_ready(nco_mux_1_auto_stream_out_1_ready),
    .auto_stream_out_1_valid(nco_mux_1_auto_stream_out_1_valid),
    .auto_stream_out_1_bits_data(nco_mux_1_auto_stream_out_1_bits_data),
    .auto_stream_out_1_bits_last(nco_mux_1_auto_stream_out_1_bits_last)
  );
  AXI4FFTBlock fft ( // @[SpectrometerTestWithoutLA.scala 80:29]
    .clock(fft_clock),
    .reset(fft_reset),
    .auto_mem_in_aw_ready(fft_auto_mem_in_aw_ready),
    .auto_mem_in_aw_valid(fft_auto_mem_in_aw_valid),
    .auto_mem_in_aw_bits_id(fft_auto_mem_in_aw_bits_id),
    .auto_mem_in_aw_bits_addr(fft_auto_mem_in_aw_bits_addr),
    .auto_mem_in_w_ready(fft_auto_mem_in_w_ready),
    .auto_mem_in_w_valid(fft_auto_mem_in_w_valid),
    .auto_mem_in_w_bits_data(fft_auto_mem_in_w_bits_data),
    .auto_mem_in_w_bits_strb(fft_auto_mem_in_w_bits_strb),
    .auto_mem_in_b_ready(fft_auto_mem_in_b_ready),
    .auto_mem_in_b_valid(fft_auto_mem_in_b_valid),
    .auto_mem_in_b_bits_id(fft_auto_mem_in_b_bits_id),
    .auto_mem_in_ar_ready(fft_auto_mem_in_ar_ready),
    .auto_mem_in_ar_valid(fft_auto_mem_in_ar_valid),
    .auto_mem_in_ar_bits_id(fft_auto_mem_in_ar_bits_id),
    .auto_mem_in_ar_bits_addr(fft_auto_mem_in_ar_bits_addr),
    .auto_mem_in_ar_bits_size(fft_auto_mem_in_ar_bits_size),
    .auto_mem_in_r_ready(fft_auto_mem_in_r_ready),
    .auto_mem_in_r_valid(fft_auto_mem_in_r_valid),
    .auto_mem_in_r_bits_id(fft_auto_mem_in_r_bits_id),
    .auto_mem_in_r_bits_data(fft_auto_mem_in_r_bits_data),
    .auto_stream_in_ready(fft_auto_stream_in_ready),
    .auto_stream_in_valid(fft_auto_stream_in_valid),
    .auto_stream_in_bits_data(fft_auto_stream_in_bits_data),
    .auto_stream_in_bits_last(fft_auto_stream_in_bits_last),
    .auto_stream_out_ready(fft_auto_stream_out_ready),
    .auto_stream_out_valid(fft_auto_stream_out_valid),
    .auto_stream_out_bits_data(fft_auto_stream_out_bits_data),
    .auto_stream_out_bits_last(fft_auto_stream_out_bits_last)
  );
  AXI4Splitter_3 fft_split ( // @[SpectrometerTestWithoutLA.scala 81:29]
    .clock(fft_split_clock),
    .reset(fft_split_reset),
    .auto_mem_in_aw_ready(fft_split_auto_mem_in_aw_ready),
    .auto_mem_in_aw_valid(fft_split_auto_mem_in_aw_valid),
    .auto_mem_in_aw_bits_id(fft_split_auto_mem_in_aw_bits_id),
    .auto_mem_in_aw_bits_addr(fft_split_auto_mem_in_aw_bits_addr),
    .auto_mem_in_w_ready(fft_split_auto_mem_in_w_ready),
    .auto_mem_in_w_valid(fft_split_auto_mem_in_w_valid),
    .auto_mem_in_w_bits_data(fft_split_auto_mem_in_w_bits_data),
    .auto_mem_in_w_bits_strb(fft_split_auto_mem_in_w_bits_strb),
    .auto_mem_in_b_ready(fft_split_auto_mem_in_b_ready),
    .auto_mem_in_b_valid(fft_split_auto_mem_in_b_valid),
    .auto_mem_in_b_bits_id(fft_split_auto_mem_in_b_bits_id),
    .auto_mem_in_ar_ready(fft_split_auto_mem_in_ar_ready),
    .auto_mem_in_ar_valid(fft_split_auto_mem_in_ar_valid),
    .auto_mem_in_ar_bits_id(fft_split_auto_mem_in_ar_bits_id),
    .auto_mem_in_ar_bits_addr(fft_split_auto_mem_in_ar_bits_addr),
    .auto_mem_in_ar_bits_size(fft_split_auto_mem_in_ar_bits_size),
    .auto_mem_in_r_ready(fft_split_auto_mem_in_r_ready),
    .auto_mem_in_r_valid(fft_split_auto_mem_in_r_valid),
    .auto_mem_in_r_bits_id(fft_split_auto_mem_in_r_bits_id),
    .auto_mem_in_r_bits_data(fft_split_auto_mem_in_r_bits_data),
    .auto_stream_in_ready(fft_split_auto_stream_in_ready),
    .auto_stream_in_valid(fft_split_auto_stream_in_valid),
    .auto_stream_in_bits_data(fft_split_auto_stream_in_bits_data),
    .auto_stream_in_bits_last(fft_split_auto_stream_in_bits_last),
    .auto_stream_out_1_ready(fft_split_auto_stream_out_1_ready),
    .auto_stream_out_1_valid(fft_split_auto_stream_out_1_valid),
    .auto_stream_out_1_bits_data(fft_split_auto_stream_out_1_bits_data),
    .auto_stream_out_1_bits_last(fft_split_auto_stream_out_1_bits_last),
    .auto_stream_out_0_ready(fft_split_auto_stream_out_0_ready),
    .auto_stream_out_0_valid(fft_split_auto_stream_out_0_valid),
    .auto_stream_out_0_bits_data(fft_split_auto_stream_out_0_bits_data),
    .auto_stream_out_0_bits_last(fft_split_auto_stream_out_0_bits_last)
  );
  AXI4StreamMux_4 fft_mux_0 ( // @[SpectrometerTestWithoutLA.scala 82:29]
    .clock(fft_mux_0_clock),
    .reset(fft_mux_0_reset),
    .auto_register_in_aw_ready(fft_mux_0_auto_register_in_aw_ready),
    .auto_register_in_aw_valid(fft_mux_0_auto_register_in_aw_valid),
    .auto_register_in_aw_bits_id(fft_mux_0_auto_register_in_aw_bits_id),
    .auto_register_in_aw_bits_addr(fft_mux_0_auto_register_in_aw_bits_addr),
    .auto_register_in_w_ready(fft_mux_0_auto_register_in_w_ready),
    .auto_register_in_w_valid(fft_mux_0_auto_register_in_w_valid),
    .auto_register_in_w_bits_data(fft_mux_0_auto_register_in_w_bits_data),
    .auto_register_in_w_bits_strb(fft_mux_0_auto_register_in_w_bits_strb),
    .auto_register_in_b_ready(fft_mux_0_auto_register_in_b_ready),
    .auto_register_in_b_valid(fft_mux_0_auto_register_in_b_valid),
    .auto_register_in_b_bits_id(fft_mux_0_auto_register_in_b_bits_id),
    .auto_register_in_ar_ready(fft_mux_0_auto_register_in_ar_ready),
    .auto_register_in_ar_valid(fft_mux_0_auto_register_in_ar_valid),
    .auto_register_in_ar_bits_id(fft_mux_0_auto_register_in_ar_bits_id),
    .auto_register_in_ar_bits_addr(fft_mux_0_auto_register_in_ar_bits_addr),
    .auto_register_in_ar_bits_size(fft_mux_0_auto_register_in_ar_bits_size),
    .auto_register_in_r_ready(fft_mux_0_auto_register_in_r_ready),
    .auto_register_in_r_valid(fft_mux_0_auto_register_in_r_valid),
    .auto_register_in_r_bits_id(fft_mux_0_auto_register_in_r_bits_id),
    .auto_register_in_r_bits_data(fft_mux_0_auto_register_in_r_bits_data),
    .auto_stream_in_2_ready(fft_mux_0_auto_stream_in_2_ready),
    .auto_stream_in_2_valid(fft_mux_0_auto_stream_in_2_valid),
    .auto_stream_in_2_bits_data(fft_mux_0_auto_stream_in_2_bits_data),
    .auto_stream_in_2_bits_last(fft_mux_0_auto_stream_in_2_bits_last),
    .auto_stream_in_1_ready(fft_mux_0_auto_stream_in_1_ready),
    .auto_stream_in_1_valid(fft_mux_0_auto_stream_in_1_valid),
    .auto_stream_in_1_bits_data(fft_mux_0_auto_stream_in_1_bits_data),
    .auto_stream_in_1_bits_last(fft_mux_0_auto_stream_in_1_bits_last),
    .auto_stream_in_0_ready(fft_mux_0_auto_stream_in_0_ready),
    .auto_stream_in_0_valid(fft_mux_0_auto_stream_in_0_valid),
    .auto_stream_in_0_bits_data(fft_mux_0_auto_stream_in_0_bits_data),
    .auto_stream_in_0_bits_last(fft_mux_0_auto_stream_in_0_bits_last),
    .auto_stream_out_0_ready(fft_mux_0_auto_stream_out_0_ready),
    .auto_stream_out_0_valid(fft_mux_0_auto_stream_out_0_valid),
    .auto_stream_out_0_bits_data(fft_mux_0_auto_stream_out_0_bits_data),
    .auto_stream_out_0_bits_last(fft_mux_0_auto_stream_out_0_bits_last)
  );
  AXI4StreamMux_5 fft_mux_1 ( // @[SpectrometerTestWithoutLA.scala 83:29]
    .clock(fft_mux_1_clock),
    .reset(fft_mux_1_reset),
    .auto_register_in_aw_ready(fft_mux_1_auto_register_in_aw_ready),
    .auto_register_in_aw_valid(fft_mux_1_auto_register_in_aw_valid),
    .auto_register_in_aw_bits_id(fft_mux_1_auto_register_in_aw_bits_id),
    .auto_register_in_aw_bits_addr(fft_mux_1_auto_register_in_aw_bits_addr),
    .auto_register_in_w_ready(fft_mux_1_auto_register_in_w_ready),
    .auto_register_in_w_valid(fft_mux_1_auto_register_in_w_valid),
    .auto_register_in_w_bits_data(fft_mux_1_auto_register_in_w_bits_data),
    .auto_register_in_w_bits_strb(fft_mux_1_auto_register_in_w_bits_strb),
    .auto_register_in_b_ready(fft_mux_1_auto_register_in_b_ready),
    .auto_register_in_b_valid(fft_mux_1_auto_register_in_b_valid),
    .auto_register_in_b_bits_id(fft_mux_1_auto_register_in_b_bits_id),
    .auto_register_in_ar_ready(fft_mux_1_auto_register_in_ar_ready),
    .auto_register_in_ar_valid(fft_mux_1_auto_register_in_ar_valid),
    .auto_register_in_ar_bits_id(fft_mux_1_auto_register_in_ar_bits_id),
    .auto_register_in_ar_bits_addr(fft_mux_1_auto_register_in_ar_bits_addr),
    .auto_register_in_ar_bits_size(fft_mux_1_auto_register_in_ar_bits_size),
    .auto_register_in_r_ready(fft_mux_1_auto_register_in_r_ready),
    .auto_register_in_r_valid(fft_mux_1_auto_register_in_r_valid),
    .auto_register_in_r_bits_id(fft_mux_1_auto_register_in_r_bits_id),
    .auto_register_in_r_bits_data(fft_mux_1_auto_register_in_r_bits_data),
    .auto_stream_in_ready(fft_mux_1_auto_stream_in_ready),
    .auto_stream_in_valid(fft_mux_1_auto_stream_in_valid),
    .auto_stream_in_bits_data(fft_mux_1_auto_stream_in_bits_data),
    .auto_stream_in_bits_last(fft_mux_1_auto_stream_in_bits_last),
    .auto_stream_out_1_ready(fft_mux_1_auto_stream_out_1_ready),
    .auto_stream_out_1_valid(fft_mux_1_auto_stream_out_1_valid),
    .auto_stream_out_1_bits_data(fft_mux_1_auto_stream_out_1_bits_data),
    .auto_stream_out_1_bits_last(fft_mux_1_auto_stream_out_1_bits_last)
  );
  AXI4LogMagMuxBlock mag ( // @[SpectrometerTestWithoutLA.scala 89:29]
    .clock(mag_clock),
    .reset(mag_reset),
    .auto_mem_in_aw_ready(mag_auto_mem_in_aw_ready),
    .auto_mem_in_aw_valid(mag_auto_mem_in_aw_valid),
    .auto_mem_in_aw_bits_id(mag_auto_mem_in_aw_bits_id),
    .auto_mem_in_aw_bits_addr(mag_auto_mem_in_aw_bits_addr),
    .auto_mem_in_w_ready(mag_auto_mem_in_w_ready),
    .auto_mem_in_w_valid(mag_auto_mem_in_w_valid),
    .auto_mem_in_w_bits_data(mag_auto_mem_in_w_bits_data),
    .auto_mem_in_w_bits_strb(mag_auto_mem_in_w_bits_strb),
    .auto_mem_in_b_ready(mag_auto_mem_in_b_ready),
    .auto_mem_in_b_valid(mag_auto_mem_in_b_valid),
    .auto_mem_in_b_bits_id(mag_auto_mem_in_b_bits_id),
    .auto_mem_in_ar_ready(mag_auto_mem_in_ar_ready),
    .auto_mem_in_ar_valid(mag_auto_mem_in_ar_valid),
    .auto_mem_in_ar_bits_id(mag_auto_mem_in_ar_bits_id),
    .auto_mem_in_ar_bits_addr(mag_auto_mem_in_ar_bits_addr),
    .auto_mem_in_ar_bits_size(mag_auto_mem_in_ar_bits_size),
    .auto_mem_in_r_ready(mag_auto_mem_in_r_ready),
    .auto_mem_in_r_valid(mag_auto_mem_in_r_valid),
    .auto_mem_in_r_bits_id(mag_auto_mem_in_r_bits_id),
    .auto_mem_in_r_bits_data(mag_auto_mem_in_r_bits_data),
    .auto_stream_in_ready(mag_auto_stream_in_ready),
    .auto_stream_in_valid(mag_auto_stream_in_valid),
    .auto_stream_in_bits_data(mag_auto_stream_in_bits_data),
    .auto_stream_in_bits_last(mag_auto_stream_in_bits_last),
    .auto_stream_out_ready(mag_auto_stream_out_ready),
    .auto_stream_out_valid(mag_auto_stream_out_valid),
    .auto_stream_out_bits_data(mag_auto_stream_out_bits_data),
    .auto_stream_out_bits_last(mag_auto_stream_out_bits_last)
  );
  AXI4Splitter_4 mag_split ( // @[SpectrometerTestWithoutLA.scala 90:29]
    .clock(mag_split_clock),
    .reset(mag_split_reset),
    .auto_mem_in_aw_ready(mag_split_auto_mem_in_aw_ready),
    .auto_mem_in_aw_valid(mag_split_auto_mem_in_aw_valid),
    .auto_mem_in_aw_bits_id(mag_split_auto_mem_in_aw_bits_id),
    .auto_mem_in_aw_bits_addr(mag_split_auto_mem_in_aw_bits_addr),
    .auto_mem_in_w_ready(mag_split_auto_mem_in_w_ready),
    .auto_mem_in_w_valid(mag_split_auto_mem_in_w_valid),
    .auto_mem_in_w_bits_data(mag_split_auto_mem_in_w_bits_data),
    .auto_mem_in_w_bits_strb(mag_split_auto_mem_in_w_bits_strb),
    .auto_mem_in_b_ready(mag_split_auto_mem_in_b_ready),
    .auto_mem_in_b_valid(mag_split_auto_mem_in_b_valid),
    .auto_mem_in_b_bits_id(mag_split_auto_mem_in_b_bits_id),
    .auto_mem_in_ar_ready(mag_split_auto_mem_in_ar_ready),
    .auto_mem_in_ar_valid(mag_split_auto_mem_in_ar_valid),
    .auto_mem_in_ar_bits_id(mag_split_auto_mem_in_ar_bits_id),
    .auto_mem_in_ar_bits_addr(mag_split_auto_mem_in_ar_bits_addr),
    .auto_mem_in_ar_bits_size(mag_split_auto_mem_in_ar_bits_size),
    .auto_mem_in_r_ready(mag_split_auto_mem_in_r_ready),
    .auto_mem_in_r_valid(mag_split_auto_mem_in_r_valid),
    .auto_mem_in_r_bits_id(mag_split_auto_mem_in_r_bits_id),
    .auto_mem_in_r_bits_data(mag_split_auto_mem_in_r_bits_data),
    .auto_stream_in_ready(mag_split_auto_stream_in_ready),
    .auto_stream_in_valid(mag_split_auto_stream_in_valid),
    .auto_stream_in_bits_data(mag_split_auto_stream_in_bits_data),
    .auto_stream_in_bits_last(mag_split_auto_stream_in_bits_last),
    .auto_stream_out_1_ready(mag_split_auto_stream_out_1_ready),
    .auto_stream_out_1_valid(mag_split_auto_stream_out_1_valid),
    .auto_stream_out_1_bits_data(mag_split_auto_stream_out_1_bits_data),
    .auto_stream_out_1_bits_last(mag_split_auto_stream_out_1_bits_last),
    .auto_stream_out_0_ready(mag_split_auto_stream_out_0_ready),
    .auto_stream_out_0_valid(mag_split_auto_stream_out_0_valid),
    .auto_stream_out_0_bits_data(mag_split_auto_stream_out_0_bits_data),
    .auto_stream_out_0_bits_last(mag_split_auto_stream_out_0_bits_last)
  );
  AXI4StreamMux_6 mag_mux_0 ( // @[SpectrometerTestWithoutLA.scala 91:29]
    .clock(mag_mux_0_clock),
    .reset(mag_mux_0_reset),
    .auto_register_in_aw_ready(mag_mux_0_auto_register_in_aw_ready),
    .auto_register_in_aw_valid(mag_mux_0_auto_register_in_aw_valid),
    .auto_register_in_aw_bits_id(mag_mux_0_auto_register_in_aw_bits_id),
    .auto_register_in_aw_bits_addr(mag_mux_0_auto_register_in_aw_bits_addr),
    .auto_register_in_w_ready(mag_mux_0_auto_register_in_w_ready),
    .auto_register_in_w_valid(mag_mux_0_auto_register_in_w_valid),
    .auto_register_in_w_bits_data(mag_mux_0_auto_register_in_w_bits_data),
    .auto_register_in_w_bits_strb(mag_mux_0_auto_register_in_w_bits_strb),
    .auto_register_in_b_ready(mag_mux_0_auto_register_in_b_ready),
    .auto_register_in_b_valid(mag_mux_0_auto_register_in_b_valid),
    .auto_register_in_b_bits_id(mag_mux_0_auto_register_in_b_bits_id),
    .auto_register_in_ar_ready(mag_mux_0_auto_register_in_ar_ready),
    .auto_register_in_ar_valid(mag_mux_0_auto_register_in_ar_valid),
    .auto_register_in_ar_bits_id(mag_mux_0_auto_register_in_ar_bits_id),
    .auto_register_in_ar_bits_addr(mag_mux_0_auto_register_in_ar_bits_addr),
    .auto_register_in_ar_bits_size(mag_mux_0_auto_register_in_ar_bits_size),
    .auto_register_in_r_ready(mag_mux_0_auto_register_in_r_ready),
    .auto_register_in_r_valid(mag_mux_0_auto_register_in_r_valid),
    .auto_register_in_r_bits_id(mag_mux_0_auto_register_in_r_bits_id),
    .auto_register_in_r_bits_data(mag_mux_0_auto_register_in_r_bits_data),
    .auto_stream_in_2_ready(mag_mux_0_auto_stream_in_2_ready),
    .auto_stream_in_2_valid(mag_mux_0_auto_stream_in_2_valid),
    .auto_stream_in_2_bits_data(mag_mux_0_auto_stream_in_2_bits_data),
    .auto_stream_in_2_bits_last(mag_mux_0_auto_stream_in_2_bits_last),
    .auto_stream_in_1_ready(mag_mux_0_auto_stream_in_1_ready),
    .auto_stream_in_1_valid(mag_mux_0_auto_stream_in_1_valid),
    .auto_stream_in_1_bits_data(mag_mux_0_auto_stream_in_1_bits_data),
    .auto_stream_in_1_bits_last(mag_mux_0_auto_stream_in_1_bits_last),
    .auto_stream_in_0_ready(mag_mux_0_auto_stream_in_0_ready),
    .auto_stream_in_0_valid(mag_mux_0_auto_stream_in_0_valid),
    .auto_stream_in_0_bits_data(mag_mux_0_auto_stream_in_0_bits_data),
    .auto_stream_in_0_bits_last(mag_mux_0_auto_stream_in_0_bits_last),
    .auto_stream_out_0_ready(mag_mux_0_auto_stream_out_0_ready),
    .auto_stream_out_0_valid(mag_mux_0_auto_stream_out_0_valid),
    .auto_stream_out_0_bits_data(mag_mux_0_auto_stream_out_0_bits_data),
    .auto_stream_out_0_bits_last(mag_mux_0_auto_stream_out_0_bits_last)
  );
  AXI4StreamMux_7 mag_mux_1 ( // @[SpectrometerTestWithoutLA.scala 92:29]
    .clock(mag_mux_1_clock),
    .reset(mag_mux_1_reset),
    .auto_register_in_aw_ready(mag_mux_1_auto_register_in_aw_ready),
    .auto_register_in_aw_valid(mag_mux_1_auto_register_in_aw_valid),
    .auto_register_in_aw_bits_id(mag_mux_1_auto_register_in_aw_bits_id),
    .auto_register_in_aw_bits_addr(mag_mux_1_auto_register_in_aw_bits_addr),
    .auto_register_in_w_ready(mag_mux_1_auto_register_in_w_ready),
    .auto_register_in_w_valid(mag_mux_1_auto_register_in_w_valid),
    .auto_register_in_w_bits_data(mag_mux_1_auto_register_in_w_bits_data),
    .auto_register_in_w_bits_strb(mag_mux_1_auto_register_in_w_bits_strb),
    .auto_register_in_b_ready(mag_mux_1_auto_register_in_b_ready),
    .auto_register_in_b_valid(mag_mux_1_auto_register_in_b_valid),
    .auto_register_in_b_bits_id(mag_mux_1_auto_register_in_b_bits_id),
    .auto_register_in_ar_ready(mag_mux_1_auto_register_in_ar_ready),
    .auto_register_in_ar_valid(mag_mux_1_auto_register_in_ar_valid),
    .auto_register_in_ar_bits_id(mag_mux_1_auto_register_in_ar_bits_id),
    .auto_register_in_ar_bits_addr(mag_mux_1_auto_register_in_ar_bits_addr),
    .auto_register_in_ar_bits_size(mag_mux_1_auto_register_in_ar_bits_size),
    .auto_register_in_r_ready(mag_mux_1_auto_register_in_r_ready),
    .auto_register_in_r_valid(mag_mux_1_auto_register_in_r_valid),
    .auto_register_in_r_bits_id(mag_mux_1_auto_register_in_r_bits_id),
    .auto_register_in_r_bits_data(mag_mux_1_auto_register_in_r_bits_data),
    .auto_stream_in_ready(mag_mux_1_auto_stream_in_ready),
    .auto_stream_in_valid(mag_mux_1_auto_stream_in_valid),
    .auto_stream_in_bits_data(mag_mux_1_auto_stream_in_bits_data),
    .auto_stream_in_bits_last(mag_mux_1_auto_stream_in_bits_last),
    .auto_stream_out_1_ready(mag_mux_1_auto_stream_out_1_ready),
    .auto_stream_out_1_valid(mag_mux_1_auto_stream_out_1_valid),
    .auto_stream_out_1_bits_data(mag_mux_1_auto_stream_out_1_bits_data),
    .auto_stream_out_1_bits_last(mag_mux_1_auto_stream_out_1_bits_last)
  );
  AccumulatorChain acc ( // @[SpectrometerTestWithoutLA.scala 98:29]
    .clock(acc_clock),
    .reset(acc_reset),
    .auto_bus_in_aw_ready(acc_auto_bus_in_aw_ready),
    .auto_bus_in_aw_valid(acc_auto_bus_in_aw_valid),
    .auto_bus_in_aw_bits_id(acc_auto_bus_in_aw_bits_id),
    .auto_bus_in_aw_bits_addr(acc_auto_bus_in_aw_bits_addr),
    .auto_bus_in_aw_bits_size(acc_auto_bus_in_aw_bits_size),
    .auto_bus_in_w_ready(acc_auto_bus_in_w_ready),
    .auto_bus_in_w_valid(acc_auto_bus_in_w_valid),
    .auto_bus_in_w_bits_data(acc_auto_bus_in_w_bits_data),
    .auto_bus_in_w_bits_strb(acc_auto_bus_in_w_bits_strb),
    .auto_bus_in_w_bits_last(acc_auto_bus_in_w_bits_last),
    .auto_bus_in_b_ready(acc_auto_bus_in_b_ready),
    .auto_bus_in_b_valid(acc_auto_bus_in_b_valid),
    .auto_bus_in_b_bits_resp(acc_auto_bus_in_b_bits_resp),
    .auto_bus_in_ar_ready(acc_auto_bus_in_ar_ready),
    .auto_bus_in_ar_valid(acc_auto_bus_in_ar_valid),
    .auto_bus_in_ar_bits_id(acc_auto_bus_in_ar_bits_id),
    .auto_bus_in_ar_bits_addr(acc_auto_bus_in_ar_bits_addr),
    .auto_bus_in_ar_bits_size(acc_auto_bus_in_ar_bits_size),
    .auto_bus_in_r_ready(acc_auto_bus_in_r_ready),
    .auto_bus_in_r_valid(acc_auto_bus_in_r_valid),
    .auto_bus_in_r_bits_data(acc_auto_bus_in_r_bits_data),
    .auto_bus_in_r_bits_resp(acc_auto_bus_in_r_bits_resp),
    .auto_bus_in_r_bits_last(acc_auto_bus_in_r_bits_last),
    .auto_dspQueue_stream_out_ready(acc_auto_dspQueue_stream_out_ready),
    .auto_dspQueue_stream_out_valid(acc_auto_dspQueue_stream_out_valid),
    .auto_dspQueue_stream_out_bits_data(acc_auto_dspQueue_stream_out_bits_data),
    .auto_dspQueue_stream_out_bits_last(acc_auto_dspQueue_stream_out_bits_last),
    .auto_accumulator_slave_in_ready(acc_auto_accumulator_slave_in_ready),
    .auto_accumulator_slave_in_valid(acc_auto_accumulator_slave_in_valid),
    .auto_accumulator_slave_in_bits_data(acc_auto_accumulator_slave_in_bits_data),
    .auto_accumulator_slave_in_bits_last(acc_auto_accumulator_slave_in_bits_last)
  );
  AXI4StreamWidthAdapater_2_to_1 widthAdapter_1 ( // @[AXI4StreamWidthAdapter.scala 82:34]
    .clock(widthAdapter_1_clock),
    .reset(widthAdapter_1_reset),
    .auto_in_ready(widthAdapter_1_auto_in_ready),
    .auto_in_valid(widthAdapter_1_auto_in_valid),
    .auto_in_bits_data(widthAdapter_1_auto_in_bits_data),
    .auto_in_bits_last(widthAdapter_1_auto_in_bits_last),
    .auto_out_ready(widthAdapter_1_auto_out_ready),
    .auto_out_valid(widthAdapter_1_auto_out_valid),
    .auto_out_bits_data(widthAdapter_1_auto_out_bits_data),
    .auto_out_bits_last(widthAdapter_1_auto_out_bits_last)
  );
  StreamBuffer_1 acc_queue ( // @[SpectrometerTestWithoutLA.scala 100:29]
    .clock(acc_queue_clock),
    .reset(acc_queue_reset),
    .auto_out_out_ready(acc_queue_auto_out_out_ready),
    .auto_out_out_valid(acc_queue_auto_out_out_valid),
    .auto_out_out_bits_data(acc_queue_auto_out_out_bits_data),
    .auto_out_out_bits_last(acc_queue_auto_out_out_bits_last),
    .auto_in_in_ready(acc_queue_auto_in_in_ready),
    .auto_in_in_valid(acc_queue_auto_in_in_valid),
    .auto_in_in_bits_data(acc_queue_auto_in_in_bits_data),
    .auto_in_in_bits_last(acc_queue_auto_in_in_bits_last)
  );
  AXI4StreamMux_8 out_mux ( // @[SpectrometerTestWithoutLA.scala 102:29]
    .clock(out_mux_clock),
    .reset(out_mux_reset),
    .auto_register_in_aw_ready(out_mux_auto_register_in_aw_ready),
    .auto_register_in_aw_valid(out_mux_auto_register_in_aw_valid),
    .auto_register_in_aw_bits_id(out_mux_auto_register_in_aw_bits_id),
    .auto_register_in_aw_bits_addr(out_mux_auto_register_in_aw_bits_addr),
    .auto_register_in_w_ready(out_mux_auto_register_in_w_ready),
    .auto_register_in_w_valid(out_mux_auto_register_in_w_valid),
    .auto_register_in_w_bits_data(out_mux_auto_register_in_w_bits_data),
    .auto_register_in_w_bits_strb(out_mux_auto_register_in_w_bits_strb),
    .auto_register_in_b_ready(out_mux_auto_register_in_b_ready),
    .auto_register_in_b_valid(out_mux_auto_register_in_b_valid),
    .auto_register_in_b_bits_id(out_mux_auto_register_in_b_bits_id),
    .auto_register_in_ar_ready(out_mux_auto_register_in_ar_ready),
    .auto_register_in_ar_valid(out_mux_auto_register_in_ar_valid),
    .auto_register_in_ar_bits_id(out_mux_auto_register_in_ar_bits_id),
    .auto_register_in_ar_bits_addr(out_mux_auto_register_in_ar_bits_addr),
    .auto_register_in_ar_bits_size(out_mux_auto_register_in_ar_bits_size),
    .auto_register_in_r_ready(out_mux_auto_register_in_r_ready),
    .auto_register_in_r_valid(out_mux_auto_register_in_r_valid),
    .auto_register_in_r_bits_id(out_mux_auto_register_in_r_bits_id),
    .auto_register_in_r_bits_data(out_mux_auto_register_in_r_bits_data),
    .auto_stream_in_6_ready(out_mux_auto_stream_in_6_ready),
    .auto_stream_in_6_valid(out_mux_auto_stream_in_6_valid),
    .auto_stream_in_6_bits_data(out_mux_auto_stream_in_6_bits_data),
    .auto_stream_in_6_bits_last(out_mux_auto_stream_in_6_bits_last),
    .auto_stream_in_5_ready(out_mux_auto_stream_in_5_ready),
    .auto_stream_in_5_valid(out_mux_auto_stream_in_5_valid),
    .auto_stream_in_5_bits_data(out_mux_auto_stream_in_5_bits_data),
    .auto_stream_in_5_bits_last(out_mux_auto_stream_in_5_bits_last),
    .auto_stream_in_4_ready(out_mux_auto_stream_in_4_ready),
    .auto_stream_in_4_valid(out_mux_auto_stream_in_4_valid),
    .auto_stream_in_4_bits_data(out_mux_auto_stream_in_4_bits_data),
    .auto_stream_in_4_bits_last(out_mux_auto_stream_in_4_bits_last),
    .auto_stream_in_3_ready(out_mux_auto_stream_in_3_ready),
    .auto_stream_in_3_valid(out_mux_auto_stream_in_3_valid),
    .auto_stream_in_3_bits_data(out_mux_auto_stream_in_3_bits_data),
    .auto_stream_in_3_bits_last(out_mux_auto_stream_in_3_bits_last),
    .auto_stream_in_2_ready(out_mux_auto_stream_in_2_ready),
    .auto_stream_in_2_valid(out_mux_auto_stream_in_2_valid),
    .auto_stream_in_2_bits_data(out_mux_auto_stream_in_2_bits_data),
    .auto_stream_in_2_bits_last(out_mux_auto_stream_in_2_bits_last),
    .auto_stream_in_1_ready(out_mux_auto_stream_in_1_ready),
    .auto_stream_in_1_valid(out_mux_auto_stream_in_1_valid),
    .auto_stream_in_1_bits_data(out_mux_auto_stream_in_1_bits_data),
    .auto_stream_in_1_bits_last(out_mux_auto_stream_in_1_bits_last),
    .auto_stream_in_0_ready(out_mux_auto_stream_in_0_ready),
    .auto_stream_in_0_valid(out_mux_auto_stream_in_0_valid),
    .auto_stream_in_0_bits_data(out_mux_auto_stream_in_0_bits_data),
    .auto_stream_in_0_bits_last(out_mux_auto_stream_in_0_bits_last),
    .auto_stream_out_1_ready(out_mux_auto_stream_out_1_ready),
    .auto_stream_out_1_valid(out_mux_auto_stream_out_1_valid),
    .auto_stream_out_1_bits_data(out_mux_auto_stream_out_1_bits_data),
    .auto_stream_out_1_bits_last(out_mux_auto_stream_out_1_bits_last),
    .auto_stream_out_0_ready(out_mux_auto_stream_out_0_ready),
    .auto_stream_out_0_valid(out_mux_auto_stream_out_0_valid),
    .auto_stream_out_0_bits_data(out_mux_auto_stream_out_0_bits_data),
    .auto_stream_out_0_bits_last(out_mux_auto_stream_out_0_bits_last)
  );
  AXI4Splitter_5 out_split ( // @[SpectrometerTestWithoutLA.scala 103:29]
    .clock(out_split_clock),
    .reset(out_split_reset),
    .auto_mem_in_aw_ready(out_split_auto_mem_in_aw_ready),
    .auto_mem_in_aw_valid(out_split_auto_mem_in_aw_valid),
    .auto_mem_in_aw_bits_id(out_split_auto_mem_in_aw_bits_id),
    .auto_mem_in_aw_bits_addr(out_split_auto_mem_in_aw_bits_addr),
    .auto_mem_in_w_ready(out_split_auto_mem_in_w_ready),
    .auto_mem_in_w_valid(out_split_auto_mem_in_w_valid),
    .auto_mem_in_w_bits_data(out_split_auto_mem_in_w_bits_data),
    .auto_mem_in_w_bits_strb(out_split_auto_mem_in_w_bits_strb),
    .auto_mem_in_b_ready(out_split_auto_mem_in_b_ready),
    .auto_mem_in_b_valid(out_split_auto_mem_in_b_valid),
    .auto_mem_in_b_bits_id(out_split_auto_mem_in_b_bits_id),
    .auto_mem_in_ar_ready(out_split_auto_mem_in_ar_ready),
    .auto_mem_in_ar_valid(out_split_auto_mem_in_ar_valid),
    .auto_mem_in_ar_bits_id(out_split_auto_mem_in_ar_bits_id),
    .auto_mem_in_ar_bits_addr(out_split_auto_mem_in_ar_bits_addr),
    .auto_mem_in_ar_bits_size(out_split_auto_mem_in_ar_bits_size),
    .auto_mem_in_r_ready(out_split_auto_mem_in_r_ready),
    .auto_mem_in_r_valid(out_split_auto_mem_in_r_valid),
    .auto_mem_in_r_bits_id(out_split_auto_mem_in_r_bits_id),
    .auto_mem_in_r_bits_data(out_split_auto_mem_in_r_bits_data),
    .auto_stream_in_ready(out_split_auto_stream_in_ready),
    .auto_stream_in_valid(out_split_auto_stream_in_valid),
    .auto_stream_in_bits_data(out_split_auto_stream_in_bits_data),
    .auto_stream_in_bits_last(out_split_auto_stream_in_bits_last),
    .auto_stream_out_ready(out_split_auto_stream_out_ready),
    .auto_stream_out_valid(out_split_auto_stream_out_valid),
    .auto_stream_out_bits_data(out_split_auto_stream_out_bits_data),
    .auto_stream_out_bits_last(out_split_auto_stream_out_bits_last)
  );
  StreamBuffer_2 out_queue ( // @[SpectrometerTestWithoutLA.scala 104:29]
    .clock(out_queue_clock),
    .reset(out_queue_reset),
    .auto_out_out_ready(out_queue_auto_out_out_ready),
    .auto_out_out_valid(out_queue_auto_out_out_valid),
    .auto_out_out_bits_data(out_queue_auto_out_out_bits_data),
    .auto_out_out_bits_last(out_queue_auto_out_out_bits_last),
    .auto_in_in_ready(out_queue_auto_in_in_ready),
    .auto_in_in_valid(out_queue_auto_in_in_valid),
    .auto_in_in_bits_data(out_queue_auto_in_in_bits_data),
    .auto_in_in_bits_last(out_queue_auto_in_in_bits_last)
  );
  AXI4StreamWidthAdapater_1_to_4 widthAdapter_2 ( // @[AXI4StreamWidthAdapter.scala 82:34]
    .clock(widthAdapter_2_clock),
    .reset(widthAdapter_2_reset),
    .auto_in_ready(widthAdapter_2_auto_in_ready),
    .auto_in_valid(widthAdapter_2_auto_in_valid),
    .auto_in_bits_data(widthAdapter_2_auto_in_bits_data),
    .auto_in_bits_last(widthAdapter_2_auto_in_bits_last),
    .auto_out_ready(widthAdapter_2_auto_out_ready),
    .auto_out_valid(widthAdapter_2_auto_out_valid),
    .auto_out_bits_data(widthAdapter_2_auto_out_bits_data),
    .auto_out_bits_last(widthAdapter_2_auto_out_bits_last)
  );
  StreamBuffer_3 uTx_queue ( // @[SpectrometerTestWithoutLA.scala 108:29]
    .clock(uTx_queue_clock),
    .reset(uTx_queue_reset),
    .auto_out_out_ready(uTx_queue_auto_out_out_ready),
    .auto_out_out_valid(uTx_queue_auto_out_out_valid),
    .auto_out_out_bits_data(uTx_queue_auto_out_out_bits_data),
    .auto_out_out_bits_last(uTx_queue_auto_out_out_bits_last),
    .auto_in_in_ready(uTx_queue_auto_in_in_ready),
    .auto_in_in_valid(uTx_queue_auto_in_in_valid),
    .auto_in_in_bits_data(uTx_queue_auto_in_in_bits_data),
    .auto_in_in_bits_last(uTx_queue_auto_in_in_bits_last)
  );
  AXI4StreamWidthAdapater_1_to_4 widthAdapter_3 ( // @[AXI4StreamWidthAdapter.scala 82:34]
    .clock(widthAdapter_3_clock),
    .reset(widthAdapter_3_reset),
    .auto_in_ready(widthAdapter_3_auto_in_ready),
    .auto_in_valid(widthAdapter_3_auto_in_valid),
    .auto_in_bits_data(widthAdapter_3_auto_in_bits_data),
    .auto_in_bits_last(widthAdapter_3_auto_in_bits_last),
    .auto_out_ready(widthAdapter_3_auto_out_ready),
    .auto_out_valid(widthAdapter_3_auto_out_valid),
    .auto_out_bits_data(widthAdapter_3_auto_out_bits_data),
    .auto_out_bits_last(widthAdapter_3_auto_out_bits_last)
  );
  AXI4StreamWidthAdapater_4_to_1 widthAdapter_4 ( // @[AXI4StreamWidthAdapter.scala 82:34]
    .clock(widthAdapter_4_clock),
    .reset(widthAdapter_4_reset),
    .auto_in_ready(widthAdapter_4_auto_in_ready),
    .auto_in_valid(widthAdapter_4_auto_in_valid),
    .auto_in_bits_data(widthAdapter_4_auto_in_bits_data),
    .auto_in_bits_last(widthAdapter_4_auto_in_bits_last),
    .auto_out_ready(widthAdapter_4_auto_out_ready),
    .auto_out_valid(widthAdapter_4_auto_out_valid),
    .auto_out_bits_data(widthAdapter_4_auto_out_bits_data),
    .auto_out_bits_last(widthAdapter_4_auto_out_bits_last)
  );
  AXI4Splitter uRx_split ( // @[SpectrometerTestWithoutLA.scala 111:29]
    .clock(uRx_split_clock),
    .reset(uRx_split_reset),
    .auto_mem_in_aw_ready(uRx_split_auto_mem_in_aw_ready),
    .auto_mem_in_aw_valid(uRx_split_auto_mem_in_aw_valid),
    .auto_mem_in_aw_bits_id(uRx_split_auto_mem_in_aw_bits_id),
    .auto_mem_in_aw_bits_addr(uRx_split_auto_mem_in_aw_bits_addr),
    .auto_mem_in_w_ready(uRx_split_auto_mem_in_w_ready),
    .auto_mem_in_w_valid(uRx_split_auto_mem_in_w_valid),
    .auto_mem_in_w_bits_data(uRx_split_auto_mem_in_w_bits_data),
    .auto_mem_in_w_bits_strb(uRx_split_auto_mem_in_w_bits_strb),
    .auto_mem_in_b_ready(uRx_split_auto_mem_in_b_ready),
    .auto_mem_in_b_valid(uRx_split_auto_mem_in_b_valid),
    .auto_mem_in_b_bits_id(uRx_split_auto_mem_in_b_bits_id),
    .auto_mem_in_ar_ready(uRx_split_auto_mem_in_ar_ready),
    .auto_mem_in_ar_valid(uRx_split_auto_mem_in_ar_valid),
    .auto_mem_in_ar_bits_id(uRx_split_auto_mem_in_ar_bits_id),
    .auto_mem_in_ar_bits_addr(uRx_split_auto_mem_in_ar_bits_addr),
    .auto_mem_in_ar_bits_size(uRx_split_auto_mem_in_ar_bits_size),
    .auto_mem_in_r_ready(uRx_split_auto_mem_in_r_ready),
    .auto_mem_in_r_valid(uRx_split_auto_mem_in_r_valid),
    .auto_mem_in_r_bits_id(uRx_split_auto_mem_in_r_bits_id),
    .auto_mem_in_r_bits_data(uRx_split_auto_mem_in_r_bits_data),
    .auto_stream_in_ready(uRx_split_auto_stream_in_ready),
    .auto_stream_in_valid(uRx_split_auto_stream_in_valid),
    .auto_stream_in_bits_data(uRx_split_auto_stream_in_bits_data),
    .auto_stream_in_bits_last(uRx_split_auto_stream_in_bits_last),
    .auto_stream_out_4_ready(uRx_split_auto_stream_out_4_ready),
    .auto_stream_out_4_valid(uRx_split_auto_stream_out_4_valid),
    .auto_stream_out_4_bits_data(uRx_split_auto_stream_out_4_bits_data),
    .auto_stream_out_4_bits_last(uRx_split_auto_stream_out_4_bits_last),
    .auto_stream_out_3_ready(uRx_split_auto_stream_out_3_ready),
    .auto_stream_out_3_valid(uRx_split_auto_stream_out_3_valid),
    .auto_stream_out_3_bits_data(uRx_split_auto_stream_out_3_bits_data),
    .auto_stream_out_3_bits_last(uRx_split_auto_stream_out_3_bits_last),
    .auto_stream_out_2_ready(uRx_split_auto_stream_out_2_ready),
    .auto_stream_out_2_valid(uRx_split_auto_stream_out_2_valid),
    .auto_stream_out_2_bits_data(uRx_split_auto_stream_out_2_bits_data),
    .auto_stream_out_2_bits_last(uRx_split_auto_stream_out_2_bits_last),
    .auto_stream_out_1_ready(uRx_split_auto_stream_out_1_ready),
    .auto_stream_out_1_valid(uRx_split_auto_stream_out_1_valid),
    .auto_stream_out_1_bits_data(uRx_split_auto_stream_out_1_bits_data),
    .auto_stream_out_1_bits_last(uRx_split_auto_stream_out_1_bits_last),
    .auto_stream_out_0_ready(uRx_split_auto_stream_out_0_ready),
    .auto_stream_out_0_valid(uRx_split_auto_stream_out_0_valid),
    .auto_stream_out_0_bits_data(uRx_split_auto_stream_out_0_bits_data),
    .auto_stream_out_0_bits_last(uRx_split_auto_stream_out_0_bits_last)
  );
  AXI4UARTBlock uart ( // @[SpectrometerTestWithoutLA.scala 112:29]
    .clock(uart_clock),
    .reset(uart_reset),
    .auto_mem_in_aw_ready(uart_auto_mem_in_aw_ready),
    .auto_mem_in_aw_valid(uart_auto_mem_in_aw_valid),
    .auto_mem_in_aw_bits_id(uart_auto_mem_in_aw_bits_id),
    .auto_mem_in_aw_bits_addr(uart_auto_mem_in_aw_bits_addr),
    .auto_mem_in_w_ready(uart_auto_mem_in_w_ready),
    .auto_mem_in_w_valid(uart_auto_mem_in_w_valid),
    .auto_mem_in_w_bits_data(uart_auto_mem_in_w_bits_data),
    .auto_mem_in_w_bits_strb(uart_auto_mem_in_w_bits_strb),
    .auto_mem_in_b_ready(uart_auto_mem_in_b_ready),
    .auto_mem_in_b_valid(uart_auto_mem_in_b_valid),
    .auto_mem_in_b_bits_id(uart_auto_mem_in_b_bits_id),
    .auto_mem_in_ar_ready(uart_auto_mem_in_ar_ready),
    .auto_mem_in_ar_valid(uart_auto_mem_in_ar_valid),
    .auto_mem_in_ar_bits_id(uart_auto_mem_in_ar_bits_id),
    .auto_mem_in_ar_bits_addr(uart_auto_mem_in_ar_bits_addr),
    .auto_mem_in_ar_bits_size(uart_auto_mem_in_ar_bits_size),
    .auto_mem_in_r_ready(uart_auto_mem_in_r_ready),
    .auto_mem_in_r_valid(uart_auto_mem_in_r_valid),
    .auto_mem_in_r_bits_id(uart_auto_mem_in_r_bits_id),
    .auto_mem_in_r_bits_data(uart_auto_mem_in_r_bits_data),
    .auto_in_in_ready(uart_auto_in_in_ready),
    .auto_in_in_valid(uart_auto_in_in_valid),
    .auto_in_in_bits_data(uart_auto_in_in_bits_data),
    .auto_out_out_ready(uart_auto_out_out_ready),
    .auto_out_out_valid(uart_auto_out_out_valid),
    .auto_out_out_bits_data(uart_auto_out_out_bits_data),
    .int_0(uart_int_0),
    .io_txd(uart_io_txd),
    .io_rxd(uart_io_rxd)
  );
  AXI4Xbar_2 bus ( // @[SpectrometerTestWithoutLA.scala 126:23]
    .clock(bus_clock),
    .reset(bus_reset),
    .auto_in_aw_ready(bus_auto_in_aw_ready),
    .auto_in_aw_valid(bus_auto_in_aw_valid),
    .auto_in_aw_bits_id(bus_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(bus_auto_in_aw_bits_addr),
    .auto_in_aw_bits_size(bus_auto_in_aw_bits_size),
    .auto_in_w_ready(bus_auto_in_w_ready),
    .auto_in_w_valid(bus_auto_in_w_valid),
    .auto_in_w_bits_data(bus_auto_in_w_bits_data),
    .auto_in_w_bits_strb(bus_auto_in_w_bits_strb),
    .auto_in_w_bits_last(bus_auto_in_w_bits_last),
    .auto_in_b_ready(bus_auto_in_b_ready),
    .auto_in_b_valid(bus_auto_in_b_valid),
    .auto_in_b_bits_resp(bus_auto_in_b_bits_resp),
    .auto_in_ar_ready(bus_auto_in_ar_ready),
    .auto_in_ar_valid(bus_auto_in_ar_valid),
    .auto_in_ar_bits_id(bus_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(bus_auto_in_ar_bits_addr),
    .auto_in_ar_bits_size(bus_auto_in_ar_bits_size),
    .auto_in_r_ready(bus_auto_in_r_ready),
    .auto_in_r_valid(bus_auto_in_r_valid),
    .auto_in_r_bits_data(bus_auto_in_r_bits_data),
    .auto_in_r_bits_resp(bus_auto_in_r_bits_resp),
    .auto_in_r_bits_last(bus_auto_in_r_bits_last),
    .auto_out_21_aw_ready(bus_auto_out_21_aw_ready),
    .auto_out_21_aw_valid(bus_auto_out_21_aw_valid),
    .auto_out_21_aw_bits_id(bus_auto_out_21_aw_bits_id),
    .auto_out_21_aw_bits_addr(bus_auto_out_21_aw_bits_addr),
    .auto_out_21_aw_bits_size(bus_auto_out_21_aw_bits_size),
    .auto_out_21_w_ready(bus_auto_out_21_w_ready),
    .auto_out_21_w_valid(bus_auto_out_21_w_valid),
    .auto_out_21_w_bits_data(bus_auto_out_21_w_bits_data),
    .auto_out_21_w_bits_strb(bus_auto_out_21_w_bits_strb),
    .auto_out_21_w_bits_last(bus_auto_out_21_w_bits_last),
    .auto_out_21_b_ready(bus_auto_out_21_b_ready),
    .auto_out_21_b_valid(bus_auto_out_21_b_valid),
    .auto_out_21_b_bits_resp(bus_auto_out_21_b_bits_resp),
    .auto_out_21_ar_ready(bus_auto_out_21_ar_ready),
    .auto_out_21_ar_valid(bus_auto_out_21_ar_valid),
    .auto_out_21_ar_bits_id(bus_auto_out_21_ar_bits_id),
    .auto_out_21_ar_bits_addr(bus_auto_out_21_ar_bits_addr),
    .auto_out_21_ar_bits_size(bus_auto_out_21_ar_bits_size),
    .auto_out_21_r_ready(bus_auto_out_21_r_ready),
    .auto_out_21_r_valid(bus_auto_out_21_r_valid),
    .auto_out_21_r_bits_data(bus_auto_out_21_r_bits_data),
    .auto_out_21_r_bits_resp(bus_auto_out_21_r_bits_resp),
    .auto_out_21_r_bits_last(bus_auto_out_21_r_bits_last),
    .auto_out_20_aw_ready(bus_auto_out_20_aw_ready),
    .auto_out_20_aw_valid(bus_auto_out_20_aw_valid),
    .auto_out_20_aw_bits_id(bus_auto_out_20_aw_bits_id),
    .auto_out_20_aw_bits_addr(bus_auto_out_20_aw_bits_addr),
    .auto_out_20_aw_bits_size(bus_auto_out_20_aw_bits_size),
    .auto_out_20_w_ready(bus_auto_out_20_w_ready),
    .auto_out_20_w_valid(bus_auto_out_20_w_valid),
    .auto_out_20_w_bits_data(bus_auto_out_20_w_bits_data),
    .auto_out_20_w_bits_strb(bus_auto_out_20_w_bits_strb),
    .auto_out_20_w_bits_last(bus_auto_out_20_w_bits_last),
    .auto_out_20_b_ready(bus_auto_out_20_b_ready),
    .auto_out_20_b_valid(bus_auto_out_20_b_valid),
    .auto_out_20_b_bits_id(bus_auto_out_20_b_bits_id),
    .auto_out_20_b_bits_resp(bus_auto_out_20_b_bits_resp),
    .auto_out_20_ar_ready(bus_auto_out_20_ar_ready),
    .auto_out_20_ar_valid(bus_auto_out_20_ar_valid),
    .auto_out_20_ar_bits_id(bus_auto_out_20_ar_bits_id),
    .auto_out_20_ar_bits_addr(bus_auto_out_20_ar_bits_addr),
    .auto_out_20_ar_bits_size(bus_auto_out_20_ar_bits_size),
    .auto_out_20_r_ready(bus_auto_out_20_r_ready),
    .auto_out_20_r_valid(bus_auto_out_20_r_valid),
    .auto_out_20_r_bits_id(bus_auto_out_20_r_bits_id),
    .auto_out_20_r_bits_data(bus_auto_out_20_r_bits_data),
    .auto_out_20_r_bits_resp(bus_auto_out_20_r_bits_resp),
    .auto_out_20_r_bits_last(bus_auto_out_20_r_bits_last),
    .auto_out_19_aw_ready(bus_auto_out_19_aw_ready),
    .auto_out_19_aw_valid(bus_auto_out_19_aw_valid),
    .auto_out_19_aw_bits_id(bus_auto_out_19_aw_bits_id),
    .auto_out_19_aw_bits_addr(bus_auto_out_19_aw_bits_addr),
    .auto_out_19_aw_bits_size(bus_auto_out_19_aw_bits_size),
    .auto_out_19_w_ready(bus_auto_out_19_w_ready),
    .auto_out_19_w_valid(bus_auto_out_19_w_valid),
    .auto_out_19_w_bits_data(bus_auto_out_19_w_bits_data),
    .auto_out_19_w_bits_strb(bus_auto_out_19_w_bits_strb),
    .auto_out_19_w_bits_last(bus_auto_out_19_w_bits_last),
    .auto_out_19_b_ready(bus_auto_out_19_b_ready),
    .auto_out_19_b_valid(bus_auto_out_19_b_valid),
    .auto_out_19_b_bits_id(bus_auto_out_19_b_bits_id),
    .auto_out_19_b_bits_resp(bus_auto_out_19_b_bits_resp),
    .auto_out_19_ar_ready(bus_auto_out_19_ar_ready),
    .auto_out_19_ar_valid(bus_auto_out_19_ar_valid),
    .auto_out_19_ar_bits_id(bus_auto_out_19_ar_bits_id),
    .auto_out_19_ar_bits_addr(bus_auto_out_19_ar_bits_addr),
    .auto_out_19_ar_bits_size(bus_auto_out_19_ar_bits_size),
    .auto_out_19_r_ready(bus_auto_out_19_r_ready),
    .auto_out_19_r_valid(bus_auto_out_19_r_valid),
    .auto_out_19_r_bits_id(bus_auto_out_19_r_bits_id),
    .auto_out_19_r_bits_data(bus_auto_out_19_r_bits_data),
    .auto_out_19_r_bits_resp(bus_auto_out_19_r_bits_resp),
    .auto_out_19_r_bits_last(bus_auto_out_19_r_bits_last),
    .auto_out_18_aw_ready(bus_auto_out_18_aw_ready),
    .auto_out_18_aw_valid(bus_auto_out_18_aw_valid),
    .auto_out_18_aw_bits_id(bus_auto_out_18_aw_bits_id),
    .auto_out_18_aw_bits_addr(bus_auto_out_18_aw_bits_addr),
    .auto_out_18_aw_bits_size(bus_auto_out_18_aw_bits_size),
    .auto_out_18_w_ready(bus_auto_out_18_w_ready),
    .auto_out_18_w_valid(bus_auto_out_18_w_valid),
    .auto_out_18_w_bits_data(bus_auto_out_18_w_bits_data),
    .auto_out_18_w_bits_strb(bus_auto_out_18_w_bits_strb),
    .auto_out_18_w_bits_last(bus_auto_out_18_w_bits_last),
    .auto_out_18_b_ready(bus_auto_out_18_b_ready),
    .auto_out_18_b_valid(bus_auto_out_18_b_valid),
    .auto_out_18_b_bits_id(bus_auto_out_18_b_bits_id),
    .auto_out_18_b_bits_resp(bus_auto_out_18_b_bits_resp),
    .auto_out_18_ar_ready(bus_auto_out_18_ar_ready),
    .auto_out_18_ar_valid(bus_auto_out_18_ar_valid),
    .auto_out_18_ar_bits_id(bus_auto_out_18_ar_bits_id),
    .auto_out_18_ar_bits_addr(bus_auto_out_18_ar_bits_addr),
    .auto_out_18_ar_bits_size(bus_auto_out_18_ar_bits_size),
    .auto_out_18_r_ready(bus_auto_out_18_r_ready),
    .auto_out_18_r_valid(bus_auto_out_18_r_valid),
    .auto_out_18_r_bits_id(bus_auto_out_18_r_bits_id),
    .auto_out_18_r_bits_data(bus_auto_out_18_r_bits_data),
    .auto_out_18_r_bits_resp(bus_auto_out_18_r_bits_resp),
    .auto_out_18_r_bits_last(bus_auto_out_18_r_bits_last),
    .auto_out_17_aw_ready(bus_auto_out_17_aw_ready),
    .auto_out_17_aw_valid(bus_auto_out_17_aw_valid),
    .auto_out_17_aw_bits_id(bus_auto_out_17_aw_bits_id),
    .auto_out_17_aw_bits_addr(bus_auto_out_17_aw_bits_addr),
    .auto_out_17_aw_bits_size(bus_auto_out_17_aw_bits_size),
    .auto_out_17_w_ready(bus_auto_out_17_w_ready),
    .auto_out_17_w_valid(bus_auto_out_17_w_valid),
    .auto_out_17_w_bits_data(bus_auto_out_17_w_bits_data),
    .auto_out_17_w_bits_strb(bus_auto_out_17_w_bits_strb),
    .auto_out_17_w_bits_last(bus_auto_out_17_w_bits_last),
    .auto_out_17_b_ready(bus_auto_out_17_b_ready),
    .auto_out_17_b_valid(bus_auto_out_17_b_valid),
    .auto_out_17_b_bits_id(bus_auto_out_17_b_bits_id),
    .auto_out_17_b_bits_resp(bus_auto_out_17_b_bits_resp),
    .auto_out_17_ar_ready(bus_auto_out_17_ar_ready),
    .auto_out_17_ar_valid(bus_auto_out_17_ar_valid),
    .auto_out_17_ar_bits_id(bus_auto_out_17_ar_bits_id),
    .auto_out_17_ar_bits_addr(bus_auto_out_17_ar_bits_addr),
    .auto_out_17_ar_bits_size(bus_auto_out_17_ar_bits_size),
    .auto_out_17_r_ready(bus_auto_out_17_r_ready),
    .auto_out_17_r_valid(bus_auto_out_17_r_valid),
    .auto_out_17_r_bits_id(bus_auto_out_17_r_bits_id),
    .auto_out_17_r_bits_data(bus_auto_out_17_r_bits_data),
    .auto_out_17_r_bits_resp(bus_auto_out_17_r_bits_resp),
    .auto_out_17_r_bits_last(bus_auto_out_17_r_bits_last),
    .auto_out_16_aw_ready(bus_auto_out_16_aw_ready),
    .auto_out_16_aw_valid(bus_auto_out_16_aw_valid),
    .auto_out_16_aw_bits_id(bus_auto_out_16_aw_bits_id),
    .auto_out_16_aw_bits_addr(bus_auto_out_16_aw_bits_addr),
    .auto_out_16_aw_bits_size(bus_auto_out_16_aw_bits_size),
    .auto_out_16_w_ready(bus_auto_out_16_w_ready),
    .auto_out_16_w_valid(bus_auto_out_16_w_valid),
    .auto_out_16_w_bits_data(bus_auto_out_16_w_bits_data),
    .auto_out_16_w_bits_strb(bus_auto_out_16_w_bits_strb),
    .auto_out_16_w_bits_last(bus_auto_out_16_w_bits_last),
    .auto_out_16_b_ready(bus_auto_out_16_b_ready),
    .auto_out_16_b_valid(bus_auto_out_16_b_valid),
    .auto_out_16_b_bits_id(bus_auto_out_16_b_bits_id),
    .auto_out_16_b_bits_resp(bus_auto_out_16_b_bits_resp),
    .auto_out_16_ar_ready(bus_auto_out_16_ar_ready),
    .auto_out_16_ar_valid(bus_auto_out_16_ar_valid),
    .auto_out_16_ar_bits_id(bus_auto_out_16_ar_bits_id),
    .auto_out_16_ar_bits_addr(bus_auto_out_16_ar_bits_addr),
    .auto_out_16_ar_bits_size(bus_auto_out_16_ar_bits_size),
    .auto_out_16_r_ready(bus_auto_out_16_r_ready),
    .auto_out_16_r_valid(bus_auto_out_16_r_valid),
    .auto_out_16_r_bits_id(bus_auto_out_16_r_bits_id),
    .auto_out_16_r_bits_data(bus_auto_out_16_r_bits_data),
    .auto_out_16_r_bits_resp(bus_auto_out_16_r_bits_resp),
    .auto_out_16_r_bits_last(bus_auto_out_16_r_bits_last),
    .auto_out_15_aw_ready(bus_auto_out_15_aw_ready),
    .auto_out_15_aw_valid(bus_auto_out_15_aw_valid),
    .auto_out_15_aw_bits_id(bus_auto_out_15_aw_bits_id),
    .auto_out_15_aw_bits_addr(bus_auto_out_15_aw_bits_addr),
    .auto_out_15_aw_bits_size(bus_auto_out_15_aw_bits_size),
    .auto_out_15_w_ready(bus_auto_out_15_w_ready),
    .auto_out_15_w_valid(bus_auto_out_15_w_valid),
    .auto_out_15_w_bits_data(bus_auto_out_15_w_bits_data),
    .auto_out_15_w_bits_strb(bus_auto_out_15_w_bits_strb),
    .auto_out_15_w_bits_last(bus_auto_out_15_w_bits_last),
    .auto_out_15_b_ready(bus_auto_out_15_b_ready),
    .auto_out_15_b_valid(bus_auto_out_15_b_valid),
    .auto_out_15_b_bits_id(bus_auto_out_15_b_bits_id),
    .auto_out_15_b_bits_resp(bus_auto_out_15_b_bits_resp),
    .auto_out_15_ar_ready(bus_auto_out_15_ar_ready),
    .auto_out_15_ar_valid(bus_auto_out_15_ar_valid),
    .auto_out_15_ar_bits_id(bus_auto_out_15_ar_bits_id),
    .auto_out_15_ar_bits_addr(bus_auto_out_15_ar_bits_addr),
    .auto_out_15_ar_bits_size(bus_auto_out_15_ar_bits_size),
    .auto_out_15_r_ready(bus_auto_out_15_r_ready),
    .auto_out_15_r_valid(bus_auto_out_15_r_valid),
    .auto_out_15_r_bits_id(bus_auto_out_15_r_bits_id),
    .auto_out_15_r_bits_data(bus_auto_out_15_r_bits_data),
    .auto_out_15_r_bits_resp(bus_auto_out_15_r_bits_resp),
    .auto_out_15_r_bits_last(bus_auto_out_15_r_bits_last),
    .auto_out_14_aw_ready(bus_auto_out_14_aw_ready),
    .auto_out_14_aw_valid(bus_auto_out_14_aw_valid),
    .auto_out_14_aw_bits_id(bus_auto_out_14_aw_bits_id),
    .auto_out_14_aw_bits_addr(bus_auto_out_14_aw_bits_addr),
    .auto_out_14_aw_bits_size(bus_auto_out_14_aw_bits_size),
    .auto_out_14_w_ready(bus_auto_out_14_w_ready),
    .auto_out_14_w_valid(bus_auto_out_14_w_valid),
    .auto_out_14_w_bits_data(bus_auto_out_14_w_bits_data),
    .auto_out_14_w_bits_strb(bus_auto_out_14_w_bits_strb),
    .auto_out_14_w_bits_last(bus_auto_out_14_w_bits_last),
    .auto_out_14_b_ready(bus_auto_out_14_b_ready),
    .auto_out_14_b_valid(bus_auto_out_14_b_valid),
    .auto_out_14_b_bits_id(bus_auto_out_14_b_bits_id),
    .auto_out_14_b_bits_resp(bus_auto_out_14_b_bits_resp),
    .auto_out_14_ar_ready(bus_auto_out_14_ar_ready),
    .auto_out_14_ar_valid(bus_auto_out_14_ar_valid),
    .auto_out_14_ar_bits_id(bus_auto_out_14_ar_bits_id),
    .auto_out_14_ar_bits_addr(bus_auto_out_14_ar_bits_addr),
    .auto_out_14_ar_bits_size(bus_auto_out_14_ar_bits_size),
    .auto_out_14_r_ready(bus_auto_out_14_r_ready),
    .auto_out_14_r_valid(bus_auto_out_14_r_valid),
    .auto_out_14_r_bits_id(bus_auto_out_14_r_bits_id),
    .auto_out_14_r_bits_data(bus_auto_out_14_r_bits_data),
    .auto_out_14_r_bits_resp(bus_auto_out_14_r_bits_resp),
    .auto_out_14_r_bits_last(bus_auto_out_14_r_bits_last),
    .auto_out_13_aw_ready(bus_auto_out_13_aw_ready),
    .auto_out_13_aw_valid(bus_auto_out_13_aw_valid),
    .auto_out_13_aw_bits_id(bus_auto_out_13_aw_bits_id),
    .auto_out_13_aw_bits_addr(bus_auto_out_13_aw_bits_addr),
    .auto_out_13_aw_bits_size(bus_auto_out_13_aw_bits_size),
    .auto_out_13_w_ready(bus_auto_out_13_w_ready),
    .auto_out_13_w_valid(bus_auto_out_13_w_valid),
    .auto_out_13_w_bits_data(bus_auto_out_13_w_bits_data),
    .auto_out_13_w_bits_strb(bus_auto_out_13_w_bits_strb),
    .auto_out_13_w_bits_last(bus_auto_out_13_w_bits_last),
    .auto_out_13_b_ready(bus_auto_out_13_b_ready),
    .auto_out_13_b_valid(bus_auto_out_13_b_valid),
    .auto_out_13_b_bits_id(bus_auto_out_13_b_bits_id),
    .auto_out_13_b_bits_resp(bus_auto_out_13_b_bits_resp),
    .auto_out_13_ar_ready(bus_auto_out_13_ar_ready),
    .auto_out_13_ar_valid(bus_auto_out_13_ar_valid),
    .auto_out_13_ar_bits_id(bus_auto_out_13_ar_bits_id),
    .auto_out_13_ar_bits_addr(bus_auto_out_13_ar_bits_addr),
    .auto_out_13_ar_bits_size(bus_auto_out_13_ar_bits_size),
    .auto_out_13_r_ready(bus_auto_out_13_r_ready),
    .auto_out_13_r_valid(bus_auto_out_13_r_valid),
    .auto_out_13_r_bits_id(bus_auto_out_13_r_bits_id),
    .auto_out_13_r_bits_data(bus_auto_out_13_r_bits_data),
    .auto_out_13_r_bits_resp(bus_auto_out_13_r_bits_resp),
    .auto_out_13_r_bits_last(bus_auto_out_13_r_bits_last),
    .auto_out_12_aw_ready(bus_auto_out_12_aw_ready),
    .auto_out_12_aw_valid(bus_auto_out_12_aw_valid),
    .auto_out_12_aw_bits_id(bus_auto_out_12_aw_bits_id),
    .auto_out_12_aw_bits_addr(bus_auto_out_12_aw_bits_addr),
    .auto_out_12_aw_bits_size(bus_auto_out_12_aw_bits_size),
    .auto_out_12_w_ready(bus_auto_out_12_w_ready),
    .auto_out_12_w_valid(bus_auto_out_12_w_valid),
    .auto_out_12_w_bits_data(bus_auto_out_12_w_bits_data),
    .auto_out_12_w_bits_strb(bus_auto_out_12_w_bits_strb),
    .auto_out_12_w_bits_last(bus_auto_out_12_w_bits_last),
    .auto_out_12_b_ready(bus_auto_out_12_b_ready),
    .auto_out_12_b_valid(bus_auto_out_12_b_valid),
    .auto_out_12_b_bits_id(bus_auto_out_12_b_bits_id),
    .auto_out_12_b_bits_resp(bus_auto_out_12_b_bits_resp),
    .auto_out_12_ar_ready(bus_auto_out_12_ar_ready),
    .auto_out_12_ar_valid(bus_auto_out_12_ar_valid),
    .auto_out_12_ar_bits_id(bus_auto_out_12_ar_bits_id),
    .auto_out_12_ar_bits_addr(bus_auto_out_12_ar_bits_addr),
    .auto_out_12_ar_bits_size(bus_auto_out_12_ar_bits_size),
    .auto_out_12_r_ready(bus_auto_out_12_r_ready),
    .auto_out_12_r_valid(bus_auto_out_12_r_valid),
    .auto_out_12_r_bits_id(bus_auto_out_12_r_bits_id),
    .auto_out_12_r_bits_data(bus_auto_out_12_r_bits_data),
    .auto_out_12_r_bits_resp(bus_auto_out_12_r_bits_resp),
    .auto_out_12_r_bits_last(bus_auto_out_12_r_bits_last),
    .auto_out_11_aw_ready(bus_auto_out_11_aw_ready),
    .auto_out_11_aw_valid(bus_auto_out_11_aw_valid),
    .auto_out_11_aw_bits_id(bus_auto_out_11_aw_bits_id),
    .auto_out_11_aw_bits_addr(bus_auto_out_11_aw_bits_addr),
    .auto_out_11_aw_bits_size(bus_auto_out_11_aw_bits_size),
    .auto_out_11_w_ready(bus_auto_out_11_w_ready),
    .auto_out_11_w_valid(bus_auto_out_11_w_valid),
    .auto_out_11_w_bits_data(bus_auto_out_11_w_bits_data),
    .auto_out_11_w_bits_strb(bus_auto_out_11_w_bits_strb),
    .auto_out_11_w_bits_last(bus_auto_out_11_w_bits_last),
    .auto_out_11_b_ready(bus_auto_out_11_b_ready),
    .auto_out_11_b_valid(bus_auto_out_11_b_valid),
    .auto_out_11_b_bits_id(bus_auto_out_11_b_bits_id),
    .auto_out_11_b_bits_resp(bus_auto_out_11_b_bits_resp),
    .auto_out_11_ar_ready(bus_auto_out_11_ar_ready),
    .auto_out_11_ar_valid(bus_auto_out_11_ar_valid),
    .auto_out_11_ar_bits_id(bus_auto_out_11_ar_bits_id),
    .auto_out_11_ar_bits_addr(bus_auto_out_11_ar_bits_addr),
    .auto_out_11_ar_bits_size(bus_auto_out_11_ar_bits_size),
    .auto_out_11_r_ready(bus_auto_out_11_r_ready),
    .auto_out_11_r_valid(bus_auto_out_11_r_valid),
    .auto_out_11_r_bits_id(bus_auto_out_11_r_bits_id),
    .auto_out_11_r_bits_data(bus_auto_out_11_r_bits_data),
    .auto_out_11_r_bits_resp(bus_auto_out_11_r_bits_resp),
    .auto_out_11_r_bits_last(bus_auto_out_11_r_bits_last),
    .auto_out_10_aw_ready(bus_auto_out_10_aw_ready),
    .auto_out_10_aw_valid(bus_auto_out_10_aw_valid),
    .auto_out_10_aw_bits_id(bus_auto_out_10_aw_bits_id),
    .auto_out_10_aw_bits_addr(bus_auto_out_10_aw_bits_addr),
    .auto_out_10_aw_bits_size(bus_auto_out_10_aw_bits_size),
    .auto_out_10_w_ready(bus_auto_out_10_w_ready),
    .auto_out_10_w_valid(bus_auto_out_10_w_valid),
    .auto_out_10_w_bits_data(bus_auto_out_10_w_bits_data),
    .auto_out_10_w_bits_strb(bus_auto_out_10_w_bits_strb),
    .auto_out_10_w_bits_last(bus_auto_out_10_w_bits_last),
    .auto_out_10_b_ready(bus_auto_out_10_b_ready),
    .auto_out_10_b_valid(bus_auto_out_10_b_valid),
    .auto_out_10_b_bits_id(bus_auto_out_10_b_bits_id),
    .auto_out_10_b_bits_resp(bus_auto_out_10_b_bits_resp),
    .auto_out_10_ar_ready(bus_auto_out_10_ar_ready),
    .auto_out_10_ar_valid(bus_auto_out_10_ar_valid),
    .auto_out_10_ar_bits_id(bus_auto_out_10_ar_bits_id),
    .auto_out_10_ar_bits_addr(bus_auto_out_10_ar_bits_addr),
    .auto_out_10_ar_bits_size(bus_auto_out_10_ar_bits_size),
    .auto_out_10_r_ready(bus_auto_out_10_r_ready),
    .auto_out_10_r_valid(bus_auto_out_10_r_valid),
    .auto_out_10_r_bits_id(bus_auto_out_10_r_bits_id),
    .auto_out_10_r_bits_data(bus_auto_out_10_r_bits_data),
    .auto_out_10_r_bits_resp(bus_auto_out_10_r_bits_resp),
    .auto_out_10_r_bits_last(bus_auto_out_10_r_bits_last),
    .auto_out_9_aw_ready(bus_auto_out_9_aw_ready),
    .auto_out_9_aw_valid(bus_auto_out_9_aw_valid),
    .auto_out_9_aw_bits_id(bus_auto_out_9_aw_bits_id),
    .auto_out_9_aw_bits_addr(bus_auto_out_9_aw_bits_addr),
    .auto_out_9_aw_bits_size(bus_auto_out_9_aw_bits_size),
    .auto_out_9_w_ready(bus_auto_out_9_w_ready),
    .auto_out_9_w_valid(bus_auto_out_9_w_valid),
    .auto_out_9_w_bits_data(bus_auto_out_9_w_bits_data),
    .auto_out_9_w_bits_strb(bus_auto_out_9_w_bits_strb),
    .auto_out_9_w_bits_last(bus_auto_out_9_w_bits_last),
    .auto_out_9_b_ready(bus_auto_out_9_b_ready),
    .auto_out_9_b_valid(bus_auto_out_9_b_valid),
    .auto_out_9_b_bits_id(bus_auto_out_9_b_bits_id),
    .auto_out_9_b_bits_resp(bus_auto_out_9_b_bits_resp),
    .auto_out_9_ar_ready(bus_auto_out_9_ar_ready),
    .auto_out_9_ar_valid(bus_auto_out_9_ar_valid),
    .auto_out_9_ar_bits_id(bus_auto_out_9_ar_bits_id),
    .auto_out_9_ar_bits_addr(bus_auto_out_9_ar_bits_addr),
    .auto_out_9_ar_bits_size(bus_auto_out_9_ar_bits_size),
    .auto_out_9_r_ready(bus_auto_out_9_r_ready),
    .auto_out_9_r_valid(bus_auto_out_9_r_valid),
    .auto_out_9_r_bits_id(bus_auto_out_9_r_bits_id),
    .auto_out_9_r_bits_data(bus_auto_out_9_r_bits_data),
    .auto_out_9_r_bits_resp(bus_auto_out_9_r_bits_resp),
    .auto_out_9_r_bits_last(bus_auto_out_9_r_bits_last),
    .auto_out_8_aw_ready(bus_auto_out_8_aw_ready),
    .auto_out_8_aw_valid(bus_auto_out_8_aw_valid),
    .auto_out_8_aw_bits_id(bus_auto_out_8_aw_bits_id),
    .auto_out_8_aw_bits_addr(bus_auto_out_8_aw_bits_addr),
    .auto_out_8_aw_bits_size(bus_auto_out_8_aw_bits_size),
    .auto_out_8_w_ready(bus_auto_out_8_w_ready),
    .auto_out_8_w_valid(bus_auto_out_8_w_valid),
    .auto_out_8_w_bits_data(bus_auto_out_8_w_bits_data),
    .auto_out_8_w_bits_strb(bus_auto_out_8_w_bits_strb),
    .auto_out_8_w_bits_last(bus_auto_out_8_w_bits_last),
    .auto_out_8_b_ready(bus_auto_out_8_b_ready),
    .auto_out_8_b_valid(bus_auto_out_8_b_valid),
    .auto_out_8_b_bits_id(bus_auto_out_8_b_bits_id),
    .auto_out_8_b_bits_resp(bus_auto_out_8_b_bits_resp),
    .auto_out_8_ar_ready(bus_auto_out_8_ar_ready),
    .auto_out_8_ar_valid(bus_auto_out_8_ar_valid),
    .auto_out_8_ar_bits_id(bus_auto_out_8_ar_bits_id),
    .auto_out_8_ar_bits_addr(bus_auto_out_8_ar_bits_addr),
    .auto_out_8_ar_bits_size(bus_auto_out_8_ar_bits_size),
    .auto_out_8_r_ready(bus_auto_out_8_r_ready),
    .auto_out_8_r_valid(bus_auto_out_8_r_valid),
    .auto_out_8_r_bits_id(bus_auto_out_8_r_bits_id),
    .auto_out_8_r_bits_data(bus_auto_out_8_r_bits_data),
    .auto_out_8_r_bits_resp(bus_auto_out_8_r_bits_resp),
    .auto_out_8_r_bits_last(bus_auto_out_8_r_bits_last),
    .auto_out_7_aw_ready(bus_auto_out_7_aw_ready),
    .auto_out_7_aw_valid(bus_auto_out_7_aw_valid),
    .auto_out_7_aw_bits_id(bus_auto_out_7_aw_bits_id),
    .auto_out_7_aw_bits_addr(bus_auto_out_7_aw_bits_addr),
    .auto_out_7_aw_bits_size(bus_auto_out_7_aw_bits_size),
    .auto_out_7_w_ready(bus_auto_out_7_w_ready),
    .auto_out_7_w_valid(bus_auto_out_7_w_valid),
    .auto_out_7_w_bits_data(bus_auto_out_7_w_bits_data),
    .auto_out_7_w_bits_strb(bus_auto_out_7_w_bits_strb),
    .auto_out_7_w_bits_last(bus_auto_out_7_w_bits_last),
    .auto_out_7_b_ready(bus_auto_out_7_b_ready),
    .auto_out_7_b_valid(bus_auto_out_7_b_valid),
    .auto_out_7_b_bits_id(bus_auto_out_7_b_bits_id),
    .auto_out_7_b_bits_resp(bus_auto_out_7_b_bits_resp),
    .auto_out_7_ar_ready(bus_auto_out_7_ar_ready),
    .auto_out_7_ar_valid(bus_auto_out_7_ar_valid),
    .auto_out_7_ar_bits_id(bus_auto_out_7_ar_bits_id),
    .auto_out_7_ar_bits_addr(bus_auto_out_7_ar_bits_addr),
    .auto_out_7_ar_bits_size(bus_auto_out_7_ar_bits_size),
    .auto_out_7_r_ready(bus_auto_out_7_r_ready),
    .auto_out_7_r_valid(bus_auto_out_7_r_valid),
    .auto_out_7_r_bits_id(bus_auto_out_7_r_bits_id),
    .auto_out_7_r_bits_data(bus_auto_out_7_r_bits_data),
    .auto_out_7_r_bits_resp(bus_auto_out_7_r_bits_resp),
    .auto_out_7_r_bits_last(bus_auto_out_7_r_bits_last),
    .auto_out_6_aw_ready(bus_auto_out_6_aw_ready),
    .auto_out_6_aw_valid(bus_auto_out_6_aw_valid),
    .auto_out_6_aw_bits_id(bus_auto_out_6_aw_bits_id),
    .auto_out_6_aw_bits_addr(bus_auto_out_6_aw_bits_addr),
    .auto_out_6_aw_bits_size(bus_auto_out_6_aw_bits_size),
    .auto_out_6_w_ready(bus_auto_out_6_w_ready),
    .auto_out_6_w_valid(bus_auto_out_6_w_valid),
    .auto_out_6_w_bits_data(bus_auto_out_6_w_bits_data),
    .auto_out_6_w_bits_strb(bus_auto_out_6_w_bits_strb),
    .auto_out_6_w_bits_last(bus_auto_out_6_w_bits_last),
    .auto_out_6_b_ready(bus_auto_out_6_b_ready),
    .auto_out_6_b_valid(bus_auto_out_6_b_valid),
    .auto_out_6_b_bits_id(bus_auto_out_6_b_bits_id),
    .auto_out_6_b_bits_resp(bus_auto_out_6_b_bits_resp),
    .auto_out_6_ar_ready(bus_auto_out_6_ar_ready),
    .auto_out_6_ar_valid(bus_auto_out_6_ar_valid),
    .auto_out_6_ar_bits_id(bus_auto_out_6_ar_bits_id),
    .auto_out_6_ar_bits_addr(bus_auto_out_6_ar_bits_addr),
    .auto_out_6_ar_bits_size(bus_auto_out_6_ar_bits_size),
    .auto_out_6_r_ready(bus_auto_out_6_r_ready),
    .auto_out_6_r_valid(bus_auto_out_6_r_valid),
    .auto_out_6_r_bits_id(bus_auto_out_6_r_bits_id),
    .auto_out_6_r_bits_data(bus_auto_out_6_r_bits_data),
    .auto_out_6_r_bits_resp(bus_auto_out_6_r_bits_resp),
    .auto_out_6_r_bits_last(bus_auto_out_6_r_bits_last),
    .auto_out_5_aw_ready(bus_auto_out_5_aw_ready),
    .auto_out_5_aw_valid(bus_auto_out_5_aw_valid),
    .auto_out_5_aw_bits_id(bus_auto_out_5_aw_bits_id),
    .auto_out_5_aw_bits_addr(bus_auto_out_5_aw_bits_addr),
    .auto_out_5_aw_bits_size(bus_auto_out_5_aw_bits_size),
    .auto_out_5_w_ready(bus_auto_out_5_w_ready),
    .auto_out_5_w_valid(bus_auto_out_5_w_valid),
    .auto_out_5_w_bits_data(bus_auto_out_5_w_bits_data),
    .auto_out_5_w_bits_strb(bus_auto_out_5_w_bits_strb),
    .auto_out_5_w_bits_last(bus_auto_out_5_w_bits_last),
    .auto_out_5_b_ready(bus_auto_out_5_b_ready),
    .auto_out_5_b_valid(bus_auto_out_5_b_valid),
    .auto_out_5_b_bits_id(bus_auto_out_5_b_bits_id),
    .auto_out_5_b_bits_resp(bus_auto_out_5_b_bits_resp),
    .auto_out_5_ar_ready(bus_auto_out_5_ar_ready),
    .auto_out_5_ar_valid(bus_auto_out_5_ar_valid),
    .auto_out_5_ar_bits_id(bus_auto_out_5_ar_bits_id),
    .auto_out_5_ar_bits_addr(bus_auto_out_5_ar_bits_addr),
    .auto_out_5_ar_bits_size(bus_auto_out_5_ar_bits_size),
    .auto_out_5_r_ready(bus_auto_out_5_r_ready),
    .auto_out_5_r_valid(bus_auto_out_5_r_valid),
    .auto_out_5_r_bits_id(bus_auto_out_5_r_bits_id),
    .auto_out_5_r_bits_data(bus_auto_out_5_r_bits_data),
    .auto_out_5_r_bits_resp(bus_auto_out_5_r_bits_resp),
    .auto_out_5_r_bits_last(bus_auto_out_5_r_bits_last),
    .auto_out_4_aw_ready(bus_auto_out_4_aw_ready),
    .auto_out_4_aw_valid(bus_auto_out_4_aw_valid),
    .auto_out_4_aw_bits_id(bus_auto_out_4_aw_bits_id),
    .auto_out_4_aw_bits_addr(bus_auto_out_4_aw_bits_addr),
    .auto_out_4_aw_bits_size(bus_auto_out_4_aw_bits_size),
    .auto_out_4_w_ready(bus_auto_out_4_w_ready),
    .auto_out_4_w_valid(bus_auto_out_4_w_valid),
    .auto_out_4_w_bits_data(bus_auto_out_4_w_bits_data),
    .auto_out_4_w_bits_strb(bus_auto_out_4_w_bits_strb),
    .auto_out_4_w_bits_last(bus_auto_out_4_w_bits_last),
    .auto_out_4_b_ready(bus_auto_out_4_b_ready),
    .auto_out_4_b_valid(bus_auto_out_4_b_valid),
    .auto_out_4_b_bits_id(bus_auto_out_4_b_bits_id),
    .auto_out_4_b_bits_resp(bus_auto_out_4_b_bits_resp),
    .auto_out_4_ar_ready(bus_auto_out_4_ar_ready),
    .auto_out_4_ar_valid(bus_auto_out_4_ar_valid),
    .auto_out_4_ar_bits_id(bus_auto_out_4_ar_bits_id),
    .auto_out_4_ar_bits_addr(bus_auto_out_4_ar_bits_addr),
    .auto_out_4_ar_bits_size(bus_auto_out_4_ar_bits_size),
    .auto_out_4_r_ready(bus_auto_out_4_r_ready),
    .auto_out_4_r_valid(bus_auto_out_4_r_valid),
    .auto_out_4_r_bits_id(bus_auto_out_4_r_bits_id),
    .auto_out_4_r_bits_data(bus_auto_out_4_r_bits_data),
    .auto_out_4_r_bits_resp(bus_auto_out_4_r_bits_resp),
    .auto_out_4_r_bits_last(bus_auto_out_4_r_bits_last),
    .auto_out_3_aw_ready(bus_auto_out_3_aw_ready),
    .auto_out_3_aw_valid(bus_auto_out_3_aw_valid),
    .auto_out_3_aw_bits_id(bus_auto_out_3_aw_bits_id),
    .auto_out_3_aw_bits_addr(bus_auto_out_3_aw_bits_addr),
    .auto_out_3_aw_bits_size(bus_auto_out_3_aw_bits_size),
    .auto_out_3_w_ready(bus_auto_out_3_w_ready),
    .auto_out_3_w_valid(bus_auto_out_3_w_valid),
    .auto_out_3_w_bits_data(bus_auto_out_3_w_bits_data),
    .auto_out_3_w_bits_strb(bus_auto_out_3_w_bits_strb),
    .auto_out_3_w_bits_last(bus_auto_out_3_w_bits_last),
    .auto_out_3_b_ready(bus_auto_out_3_b_ready),
    .auto_out_3_b_valid(bus_auto_out_3_b_valid),
    .auto_out_3_b_bits_id(bus_auto_out_3_b_bits_id),
    .auto_out_3_b_bits_resp(bus_auto_out_3_b_bits_resp),
    .auto_out_3_ar_ready(bus_auto_out_3_ar_ready),
    .auto_out_3_ar_valid(bus_auto_out_3_ar_valid),
    .auto_out_3_ar_bits_id(bus_auto_out_3_ar_bits_id),
    .auto_out_3_ar_bits_addr(bus_auto_out_3_ar_bits_addr),
    .auto_out_3_ar_bits_size(bus_auto_out_3_ar_bits_size),
    .auto_out_3_r_ready(bus_auto_out_3_r_ready),
    .auto_out_3_r_valid(bus_auto_out_3_r_valid),
    .auto_out_3_r_bits_id(bus_auto_out_3_r_bits_id),
    .auto_out_3_r_bits_data(bus_auto_out_3_r_bits_data),
    .auto_out_3_r_bits_resp(bus_auto_out_3_r_bits_resp),
    .auto_out_3_r_bits_last(bus_auto_out_3_r_bits_last),
    .auto_out_2_aw_ready(bus_auto_out_2_aw_ready),
    .auto_out_2_aw_valid(bus_auto_out_2_aw_valid),
    .auto_out_2_aw_bits_id(bus_auto_out_2_aw_bits_id),
    .auto_out_2_aw_bits_addr(bus_auto_out_2_aw_bits_addr),
    .auto_out_2_aw_bits_size(bus_auto_out_2_aw_bits_size),
    .auto_out_2_w_ready(bus_auto_out_2_w_ready),
    .auto_out_2_w_valid(bus_auto_out_2_w_valid),
    .auto_out_2_w_bits_data(bus_auto_out_2_w_bits_data),
    .auto_out_2_w_bits_strb(bus_auto_out_2_w_bits_strb),
    .auto_out_2_w_bits_last(bus_auto_out_2_w_bits_last),
    .auto_out_2_b_ready(bus_auto_out_2_b_ready),
    .auto_out_2_b_valid(bus_auto_out_2_b_valid),
    .auto_out_2_b_bits_id(bus_auto_out_2_b_bits_id),
    .auto_out_2_b_bits_resp(bus_auto_out_2_b_bits_resp),
    .auto_out_2_ar_ready(bus_auto_out_2_ar_ready),
    .auto_out_2_ar_valid(bus_auto_out_2_ar_valid),
    .auto_out_2_ar_bits_id(bus_auto_out_2_ar_bits_id),
    .auto_out_2_ar_bits_addr(bus_auto_out_2_ar_bits_addr),
    .auto_out_2_ar_bits_size(bus_auto_out_2_ar_bits_size),
    .auto_out_2_r_ready(bus_auto_out_2_r_ready),
    .auto_out_2_r_valid(bus_auto_out_2_r_valid),
    .auto_out_2_r_bits_id(bus_auto_out_2_r_bits_id),
    .auto_out_2_r_bits_data(bus_auto_out_2_r_bits_data),
    .auto_out_2_r_bits_resp(bus_auto_out_2_r_bits_resp),
    .auto_out_2_r_bits_last(bus_auto_out_2_r_bits_last),
    .auto_out_1_aw_ready(bus_auto_out_1_aw_ready),
    .auto_out_1_aw_valid(bus_auto_out_1_aw_valid),
    .auto_out_1_aw_bits_id(bus_auto_out_1_aw_bits_id),
    .auto_out_1_aw_bits_addr(bus_auto_out_1_aw_bits_addr),
    .auto_out_1_aw_bits_size(bus_auto_out_1_aw_bits_size),
    .auto_out_1_w_ready(bus_auto_out_1_w_ready),
    .auto_out_1_w_valid(bus_auto_out_1_w_valid),
    .auto_out_1_w_bits_data(bus_auto_out_1_w_bits_data),
    .auto_out_1_w_bits_strb(bus_auto_out_1_w_bits_strb),
    .auto_out_1_w_bits_last(bus_auto_out_1_w_bits_last),
    .auto_out_1_b_ready(bus_auto_out_1_b_ready),
    .auto_out_1_b_valid(bus_auto_out_1_b_valid),
    .auto_out_1_b_bits_id(bus_auto_out_1_b_bits_id),
    .auto_out_1_b_bits_resp(bus_auto_out_1_b_bits_resp),
    .auto_out_1_ar_ready(bus_auto_out_1_ar_ready),
    .auto_out_1_ar_valid(bus_auto_out_1_ar_valid),
    .auto_out_1_ar_bits_id(bus_auto_out_1_ar_bits_id),
    .auto_out_1_ar_bits_addr(bus_auto_out_1_ar_bits_addr),
    .auto_out_1_ar_bits_size(bus_auto_out_1_ar_bits_size),
    .auto_out_1_r_ready(bus_auto_out_1_r_ready),
    .auto_out_1_r_valid(bus_auto_out_1_r_valid),
    .auto_out_1_r_bits_id(bus_auto_out_1_r_bits_id),
    .auto_out_1_r_bits_data(bus_auto_out_1_r_bits_data),
    .auto_out_1_r_bits_resp(bus_auto_out_1_r_bits_resp),
    .auto_out_1_r_bits_last(bus_auto_out_1_r_bits_last),
    .auto_out_0_aw_ready(bus_auto_out_0_aw_ready),
    .auto_out_0_aw_valid(bus_auto_out_0_aw_valid),
    .auto_out_0_aw_bits_id(bus_auto_out_0_aw_bits_id),
    .auto_out_0_aw_bits_addr(bus_auto_out_0_aw_bits_addr),
    .auto_out_0_aw_bits_size(bus_auto_out_0_aw_bits_size),
    .auto_out_0_w_ready(bus_auto_out_0_w_ready),
    .auto_out_0_w_valid(bus_auto_out_0_w_valid),
    .auto_out_0_w_bits_data(bus_auto_out_0_w_bits_data),
    .auto_out_0_w_bits_strb(bus_auto_out_0_w_bits_strb),
    .auto_out_0_w_bits_last(bus_auto_out_0_w_bits_last),
    .auto_out_0_b_ready(bus_auto_out_0_b_ready),
    .auto_out_0_b_valid(bus_auto_out_0_b_valid),
    .auto_out_0_b_bits_id(bus_auto_out_0_b_bits_id),
    .auto_out_0_b_bits_resp(bus_auto_out_0_b_bits_resp),
    .auto_out_0_ar_ready(bus_auto_out_0_ar_ready),
    .auto_out_0_ar_valid(bus_auto_out_0_ar_valid),
    .auto_out_0_ar_bits_id(bus_auto_out_0_ar_bits_id),
    .auto_out_0_ar_bits_addr(bus_auto_out_0_ar_bits_addr),
    .auto_out_0_ar_bits_size(bus_auto_out_0_ar_bits_size),
    .auto_out_0_r_ready(bus_auto_out_0_r_ready),
    .auto_out_0_r_valid(bus_auto_out_0_r_valid),
    .auto_out_0_r_bits_id(bus_auto_out_0_r_bits_id),
    .auto_out_0_r_bits_data(bus_auto_out_0_r_bits_data),
    .auto_out_0_r_bits_resp(bus_auto_out_0_r_bits_resp),
    .auto_out_0_r_bits_last(bus_auto_out_0_r_bits_last)
  );
  AXI4Buffer axi4buf ( // @[Buffer.scala 58:29]
    .clock(axi4buf_clock),
    .reset(axi4buf_reset),
    .auto_in_aw_ready(axi4buf_auto_in_aw_ready),
    .auto_in_aw_valid(axi4buf_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4buf_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4buf_auto_in_aw_bits_addr),
    .auto_in_aw_bits_size(axi4buf_auto_in_aw_bits_size),
    .auto_in_w_ready(axi4buf_auto_in_w_ready),
    .auto_in_w_valid(axi4buf_auto_in_w_valid),
    .auto_in_w_bits_data(axi4buf_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi4buf_auto_in_w_bits_strb),
    .auto_in_w_bits_last(axi4buf_auto_in_w_bits_last),
    .auto_in_b_ready(axi4buf_auto_in_b_ready),
    .auto_in_b_valid(axi4buf_auto_in_b_valid),
    .auto_in_b_bits_id(axi4buf_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi4buf_auto_in_b_bits_resp),
    .auto_in_ar_ready(axi4buf_auto_in_ar_ready),
    .auto_in_ar_valid(axi4buf_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4buf_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4buf_auto_in_ar_bits_addr),
    .auto_in_ar_bits_size(axi4buf_auto_in_ar_bits_size),
    .auto_in_r_ready(axi4buf_auto_in_r_ready),
    .auto_in_r_valid(axi4buf_auto_in_r_valid),
    .auto_in_r_bits_id(axi4buf_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4buf_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4buf_auto_in_r_bits_resp),
    .auto_in_r_bits_last(axi4buf_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4buf_auto_out_aw_ready),
    .auto_out_aw_valid(axi4buf_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4buf_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4buf_auto_out_aw_bits_addr),
    .auto_out_w_ready(axi4buf_auto_out_w_ready),
    .auto_out_w_valid(axi4buf_auto_out_w_valid),
    .auto_out_w_bits_data(axi4buf_auto_out_w_bits_data),
    .auto_out_w_bits_strb(axi4buf_auto_out_w_bits_strb),
    .auto_out_w_bits_last(axi4buf_auto_out_w_bits_last),
    .auto_out_b_ready(axi4buf_auto_out_b_ready),
    .auto_out_b_valid(axi4buf_auto_out_b_valid),
    .auto_out_b_bits_id(axi4buf_auto_out_b_bits_id),
    .auto_out_b_bits_resp(axi4buf_auto_out_b_bits_resp),
    .auto_out_ar_ready(axi4buf_auto_out_ar_ready),
    .auto_out_ar_valid(axi4buf_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4buf_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4buf_auto_out_ar_bits_addr),
    .auto_out_ar_bits_size(axi4buf_auto_out_ar_bits_size),
    .auto_out_r_ready(axi4buf_auto_out_r_ready),
    .auto_out_r_valid(axi4buf_auto_out_r_valid),
    .auto_out_r_bits_id(axi4buf_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4buf_auto_out_r_bits_data),
    .auto_out_r_bits_resp(axi4buf_auto_out_r_bits_resp),
    .auto_out_r_bits_last(axi4buf_auto_out_r_bits_last)
  );
  AXI4Buffer axi4buf_1 ( // @[Buffer.scala 58:29]
    .clock(axi4buf_1_clock),
    .reset(axi4buf_1_reset),
    .auto_in_aw_ready(axi4buf_1_auto_in_aw_ready),
    .auto_in_aw_valid(axi4buf_1_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4buf_1_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4buf_1_auto_in_aw_bits_addr),
    .auto_in_aw_bits_size(axi4buf_1_auto_in_aw_bits_size),
    .auto_in_w_ready(axi4buf_1_auto_in_w_ready),
    .auto_in_w_valid(axi4buf_1_auto_in_w_valid),
    .auto_in_w_bits_data(axi4buf_1_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi4buf_1_auto_in_w_bits_strb),
    .auto_in_w_bits_last(axi4buf_1_auto_in_w_bits_last),
    .auto_in_b_ready(axi4buf_1_auto_in_b_ready),
    .auto_in_b_valid(axi4buf_1_auto_in_b_valid),
    .auto_in_b_bits_id(axi4buf_1_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi4buf_1_auto_in_b_bits_resp),
    .auto_in_ar_ready(axi4buf_1_auto_in_ar_ready),
    .auto_in_ar_valid(axi4buf_1_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4buf_1_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4buf_1_auto_in_ar_bits_addr),
    .auto_in_ar_bits_size(axi4buf_1_auto_in_ar_bits_size),
    .auto_in_r_ready(axi4buf_1_auto_in_r_ready),
    .auto_in_r_valid(axi4buf_1_auto_in_r_valid),
    .auto_in_r_bits_id(axi4buf_1_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4buf_1_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4buf_1_auto_in_r_bits_resp),
    .auto_in_r_bits_last(axi4buf_1_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4buf_1_auto_out_aw_ready),
    .auto_out_aw_valid(axi4buf_1_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4buf_1_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4buf_1_auto_out_aw_bits_addr),
    .auto_out_w_ready(axi4buf_1_auto_out_w_ready),
    .auto_out_w_valid(axi4buf_1_auto_out_w_valid),
    .auto_out_w_bits_data(axi4buf_1_auto_out_w_bits_data),
    .auto_out_w_bits_strb(axi4buf_1_auto_out_w_bits_strb),
    .auto_out_w_bits_last(axi4buf_1_auto_out_w_bits_last),
    .auto_out_b_ready(axi4buf_1_auto_out_b_ready),
    .auto_out_b_valid(axi4buf_1_auto_out_b_valid),
    .auto_out_b_bits_id(axi4buf_1_auto_out_b_bits_id),
    .auto_out_b_bits_resp(axi4buf_1_auto_out_b_bits_resp),
    .auto_out_ar_ready(axi4buf_1_auto_out_ar_ready),
    .auto_out_ar_valid(axi4buf_1_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4buf_1_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4buf_1_auto_out_ar_bits_addr),
    .auto_out_ar_bits_size(axi4buf_1_auto_out_ar_bits_size),
    .auto_out_r_ready(axi4buf_1_auto_out_r_ready),
    .auto_out_r_valid(axi4buf_1_auto_out_r_valid),
    .auto_out_r_bits_id(axi4buf_1_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4buf_1_auto_out_r_bits_data),
    .auto_out_r_bits_resp(axi4buf_1_auto_out_r_bits_resp),
    .auto_out_r_bits_last(axi4buf_1_auto_out_r_bits_last)
  );
  AXI4Buffer axi4buf_2 ( // @[Buffer.scala 58:29]
    .clock(axi4buf_2_clock),
    .reset(axi4buf_2_reset),
    .auto_in_aw_ready(axi4buf_2_auto_in_aw_ready),
    .auto_in_aw_valid(axi4buf_2_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4buf_2_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4buf_2_auto_in_aw_bits_addr),
    .auto_in_aw_bits_size(axi4buf_2_auto_in_aw_bits_size),
    .auto_in_w_ready(axi4buf_2_auto_in_w_ready),
    .auto_in_w_valid(axi4buf_2_auto_in_w_valid),
    .auto_in_w_bits_data(axi4buf_2_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi4buf_2_auto_in_w_bits_strb),
    .auto_in_w_bits_last(axi4buf_2_auto_in_w_bits_last),
    .auto_in_b_ready(axi4buf_2_auto_in_b_ready),
    .auto_in_b_valid(axi4buf_2_auto_in_b_valid),
    .auto_in_b_bits_id(axi4buf_2_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi4buf_2_auto_in_b_bits_resp),
    .auto_in_ar_ready(axi4buf_2_auto_in_ar_ready),
    .auto_in_ar_valid(axi4buf_2_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4buf_2_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4buf_2_auto_in_ar_bits_addr),
    .auto_in_ar_bits_size(axi4buf_2_auto_in_ar_bits_size),
    .auto_in_r_ready(axi4buf_2_auto_in_r_ready),
    .auto_in_r_valid(axi4buf_2_auto_in_r_valid),
    .auto_in_r_bits_id(axi4buf_2_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4buf_2_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4buf_2_auto_in_r_bits_resp),
    .auto_in_r_bits_last(axi4buf_2_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4buf_2_auto_out_aw_ready),
    .auto_out_aw_valid(axi4buf_2_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4buf_2_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4buf_2_auto_out_aw_bits_addr),
    .auto_out_w_ready(axi4buf_2_auto_out_w_ready),
    .auto_out_w_valid(axi4buf_2_auto_out_w_valid),
    .auto_out_w_bits_data(axi4buf_2_auto_out_w_bits_data),
    .auto_out_w_bits_strb(axi4buf_2_auto_out_w_bits_strb),
    .auto_out_w_bits_last(axi4buf_2_auto_out_w_bits_last),
    .auto_out_b_ready(axi4buf_2_auto_out_b_ready),
    .auto_out_b_valid(axi4buf_2_auto_out_b_valid),
    .auto_out_b_bits_id(axi4buf_2_auto_out_b_bits_id),
    .auto_out_b_bits_resp(axi4buf_2_auto_out_b_bits_resp),
    .auto_out_ar_ready(axi4buf_2_auto_out_ar_ready),
    .auto_out_ar_valid(axi4buf_2_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4buf_2_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4buf_2_auto_out_ar_bits_addr),
    .auto_out_ar_bits_size(axi4buf_2_auto_out_ar_bits_size),
    .auto_out_r_ready(axi4buf_2_auto_out_r_ready),
    .auto_out_r_valid(axi4buf_2_auto_out_r_valid),
    .auto_out_r_bits_id(axi4buf_2_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4buf_2_auto_out_r_bits_data),
    .auto_out_r_bits_resp(axi4buf_2_auto_out_r_bits_resp),
    .auto_out_r_bits_last(axi4buf_2_auto_out_r_bits_last)
  );
  AXI4Buffer axi4buf_3 ( // @[Buffer.scala 58:29]
    .clock(axi4buf_3_clock),
    .reset(axi4buf_3_reset),
    .auto_in_aw_ready(axi4buf_3_auto_in_aw_ready),
    .auto_in_aw_valid(axi4buf_3_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4buf_3_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4buf_3_auto_in_aw_bits_addr),
    .auto_in_aw_bits_size(axi4buf_3_auto_in_aw_bits_size),
    .auto_in_w_ready(axi4buf_3_auto_in_w_ready),
    .auto_in_w_valid(axi4buf_3_auto_in_w_valid),
    .auto_in_w_bits_data(axi4buf_3_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi4buf_3_auto_in_w_bits_strb),
    .auto_in_w_bits_last(axi4buf_3_auto_in_w_bits_last),
    .auto_in_b_ready(axi4buf_3_auto_in_b_ready),
    .auto_in_b_valid(axi4buf_3_auto_in_b_valid),
    .auto_in_b_bits_id(axi4buf_3_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi4buf_3_auto_in_b_bits_resp),
    .auto_in_ar_ready(axi4buf_3_auto_in_ar_ready),
    .auto_in_ar_valid(axi4buf_3_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4buf_3_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4buf_3_auto_in_ar_bits_addr),
    .auto_in_ar_bits_size(axi4buf_3_auto_in_ar_bits_size),
    .auto_in_r_ready(axi4buf_3_auto_in_r_ready),
    .auto_in_r_valid(axi4buf_3_auto_in_r_valid),
    .auto_in_r_bits_id(axi4buf_3_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4buf_3_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4buf_3_auto_in_r_bits_resp),
    .auto_in_r_bits_last(axi4buf_3_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4buf_3_auto_out_aw_ready),
    .auto_out_aw_valid(axi4buf_3_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4buf_3_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4buf_3_auto_out_aw_bits_addr),
    .auto_out_w_ready(axi4buf_3_auto_out_w_ready),
    .auto_out_w_valid(axi4buf_3_auto_out_w_valid),
    .auto_out_w_bits_data(axi4buf_3_auto_out_w_bits_data),
    .auto_out_w_bits_strb(axi4buf_3_auto_out_w_bits_strb),
    .auto_out_w_bits_last(axi4buf_3_auto_out_w_bits_last),
    .auto_out_b_ready(axi4buf_3_auto_out_b_ready),
    .auto_out_b_valid(axi4buf_3_auto_out_b_valid),
    .auto_out_b_bits_id(axi4buf_3_auto_out_b_bits_id),
    .auto_out_b_bits_resp(axi4buf_3_auto_out_b_bits_resp),
    .auto_out_ar_ready(axi4buf_3_auto_out_ar_ready),
    .auto_out_ar_valid(axi4buf_3_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4buf_3_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4buf_3_auto_out_ar_bits_addr),
    .auto_out_ar_bits_size(axi4buf_3_auto_out_ar_bits_size),
    .auto_out_r_ready(axi4buf_3_auto_out_r_ready),
    .auto_out_r_valid(axi4buf_3_auto_out_r_valid),
    .auto_out_r_bits_id(axi4buf_3_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4buf_3_auto_out_r_bits_data),
    .auto_out_r_bits_resp(axi4buf_3_auto_out_r_bits_resp),
    .auto_out_r_bits_last(axi4buf_3_auto_out_r_bits_last)
  );
  AXI4Buffer axi4buf_4 ( // @[Buffer.scala 58:29]
    .clock(axi4buf_4_clock),
    .reset(axi4buf_4_reset),
    .auto_in_aw_ready(axi4buf_4_auto_in_aw_ready),
    .auto_in_aw_valid(axi4buf_4_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4buf_4_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4buf_4_auto_in_aw_bits_addr),
    .auto_in_aw_bits_size(axi4buf_4_auto_in_aw_bits_size),
    .auto_in_w_ready(axi4buf_4_auto_in_w_ready),
    .auto_in_w_valid(axi4buf_4_auto_in_w_valid),
    .auto_in_w_bits_data(axi4buf_4_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi4buf_4_auto_in_w_bits_strb),
    .auto_in_w_bits_last(axi4buf_4_auto_in_w_bits_last),
    .auto_in_b_ready(axi4buf_4_auto_in_b_ready),
    .auto_in_b_valid(axi4buf_4_auto_in_b_valid),
    .auto_in_b_bits_id(axi4buf_4_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi4buf_4_auto_in_b_bits_resp),
    .auto_in_ar_ready(axi4buf_4_auto_in_ar_ready),
    .auto_in_ar_valid(axi4buf_4_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4buf_4_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4buf_4_auto_in_ar_bits_addr),
    .auto_in_ar_bits_size(axi4buf_4_auto_in_ar_bits_size),
    .auto_in_r_ready(axi4buf_4_auto_in_r_ready),
    .auto_in_r_valid(axi4buf_4_auto_in_r_valid),
    .auto_in_r_bits_id(axi4buf_4_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4buf_4_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4buf_4_auto_in_r_bits_resp),
    .auto_in_r_bits_last(axi4buf_4_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4buf_4_auto_out_aw_ready),
    .auto_out_aw_valid(axi4buf_4_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4buf_4_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4buf_4_auto_out_aw_bits_addr),
    .auto_out_w_ready(axi4buf_4_auto_out_w_ready),
    .auto_out_w_valid(axi4buf_4_auto_out_w_valid),
    .auto_out_w_bits_data(axi4buf_4_auto_out_w_bits_data),
    .auto_out_w_bits_strb(axi4buf_4_auto_out_w_bits_strb),
    .auto_out_w_bits_last(axi4buf_4_auto_out_w_bits_last),
    .auto_out_b_ready(axi4buf_4_auto_out_b_ready),
    .auto_out_b_valid(axi4buf_4_auto_out_b_valid),
    .auto_out_b_bits_id(axi4buf_4_auto_out_b_bits_id),
    .auto_out_b_bits_resp(axi4buf_4_auto_out_b_bits_resp),
    .auto_out_ar_ready(axi4buf_4_auto_out_ar_ready),
    .auto_out_ar_valid(axi4buf_4_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4buf_4_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4buf_4_auto_out_ar_bits_addr),
    .auto_out_ar_bits_size(axi4buf_4_auto_out_ar_bits_size),
    .auto_out_r_ready(axi4buf_4_auto_out_r_ready),
    .auto_out_r_valid(axi4buf_4_auto_out_r_valid),
    .auto_out_r_bits_id(axi4buf_4_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4buf_4_auto_out_r_bits_data),
    .auto_out_r_bits_resp(axi4buf_4_auto_out_r_bits_resp),
    .auto_out_r_bits_last(axi4buf_4_auto_out_r_bits_last)
  );
  AXI4Buffer axi4buf_5 ( // @[Buffer.scala 58:29]
    .clock(axi4buf_5_clock),
    .reset(axi4buf_5_reset),
    .auto_in_aw_ready(axi4buf_5_auto_in_aw_ready),
    .auto_in_aw_valid(axi4buf_5_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4buf_5_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4buf_5_auto_in_aw_bits_addr),
    .auto_in_aw_bits_size(axi4buf_5_auto_in_aw_bits_size),
    .auto_in_w_ready(axi4buf_5_auto_in_w_ready),
    .auto_in_w_valid(axi4buf_5_auto_in_w_valid),
    .auto_in_w_bits_data(axi4buf_5_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi4buf_5_auto_in_w_bits_strb),
    .auto_in_w_bits_last(axi4buf_5_auto_in_w_bits_last),
    .auto_in_b_ready(axi4buf_5_auto_in_b_ready),
    .auto_in_b_valid(axi4buf_5_auto_in_b_valid),
    .auto_in_b_bits_id(axi4buf_5_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi4buf_5_auto_in_b_bits_resp),
    .auto_in_ar_ready(axi4buf_5_auto_in_ar_ready),
    .auto_in_ar_valid(axi4buf_5_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4buf_5_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4buf_5_auto_in_ar_bits_addr),
    .auto_in_ar_bits_size(axi4buf_5_auto_in_ar_bits_size),
    .auto_in_r_ready(axi4buf_5_auto_in_r_ready),
    .auto_in_r_valid(axi4buf_5_auto_in_r_valid),
    .auto_in_r_bits_id(axi4buf_5_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4buf_5_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4buf_5_auto_in_r_bits_resp),
    .auto_in_r_bits_last(axi4buf_5_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4buf_5_auto_out_aw_ready),
    .auto_out_aw_valid(axi4buf_5_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4buf_5_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4buf_5_auto_out_aw_bits_addr),
    .auto_out_w_ready(axi4buf_5_auto_out_w_ready),
    .auto_out_w_valid(axi4buf_5_auto_out_w_valid),
    .auto_out_w_bits_data(axi4buf_5_auto_out_w_bits_data),
    .auto_out_w_bits_strb(axi4buf_5_auto_out_w_bits_strb),
    .auto_out_w_bits_last(axi4buf_5_auto_out_w_bits_last),
    .auto_out_b_ready(axi4buf_5_auto_out_b_ready),
    .auto_out_b_valid(axi4buf_5_auto_out_b_valid),
    .auto_out_b_bits_id(axi4buf_5_auto_out_b_bits_id),
    .auto_out_b_bits_resp(axi4buf_5_auto_out_b_bits_resp),
    .auto_out_ar_ready(axi4buf_5_auto_out_ar_ready),
    .auto_out_ar_valid(axi4buf_5_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4buf_5_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4buf_5_auto_out_ar_bits_addr),
    .auto_out_ar_bits_size(axi4buf_5_auto_out_ar_bits_size),
    .auto_out_r_ready(axi4buf_5_auto_out_r_ready),
    .auto_out_r_valid(axi4buf_5_auto_out_r_valid),
    .auto_out_r_bits_id(axi4buf_5_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4buf_5_auto_out_r_bits_data),
    .auto_out_r_bits_resp(axi4buf_5_auto_out_r_bits_resp),
    .auto_out_r_bits_last(axi4buf_5_auto_out_r_bits_last)
  );
  AXI4Buffer axi4buf_6 ( // @[Buffer.scala 58:29]
    .clock(axi4buf_6_clock),
    .reset(axi4buf_6_reset),
    .auto_in_aw_ready(axi4buf_6_auto_in_aw_ready),
    .auto_in_aw_valid(axi4buf_6_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4buf_6_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4buf_6_auto_in_aw_bits_addr),
    .auto_in_aw_bits_size(axi4buf_6_auto_in_aw_bits_size),
    .auto_in_w_ready(axi4buf_6_auto_in_w_ready),
    .auto_in_w_valid(axi4buf_6_auto_in_w_valid),
    .auto_in_w_bits_data(axi4buf_6_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi4buf_6_auto_in_w_bits_strb),
    .auto_in_w_bits_last(axi4buf_6_auto_in_w_bits_last),
    .auto_in_b_ready(axi4buf_6_auto_in_b_ready),
    .auto_in_b_valid(axi4buf_6_auto_in_b_valid),
    .auto_in_b_bits_id(axi4buf_6_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi4buf_6_auto_in_b_bits_resp),
    .auto_in_ar_ready(axi4buf_6_auto_in_ar_ready),
    .auto_in_ar_valid(axi4buf_6_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4buf_6_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4buf_6_auto_in_ar_bits_addr),
    .auto_in_ar_bits_size(axi4buf_6_auto_in_ar_bits_size),
    .auto_in_r_ready(axi4buf_6_auto_in_r_ready),
    .auto_in_r_valid(axi4buf_6_auto_in_r_valid),
    .auto_in_r_bits_id(axi4buf_6_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4buf_6_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4buf_6_auto_in_r_bits_resp),
    .auto_in_r_bits_last(axi4buf_6_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4buf_6_auto_out_aw_ready),
    .auto_out_aw_valid(axi4buf_6_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4buf_6_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4buf_6_auto_out_aw_bits_addr),
    .auto_out_w_ready(axi4buf_6_auto_out_w_ready),
    .auto_out_w_valid(axi4buf_6_auto_out_w_valid),
    .auto_out_w_bits_data(axi4buf_6_auto_out_w_bits_data),
    .auto_out_w_bits_strb(axi4buf_6_auto_out_w_bits_strb),
    .auto_out_w_bits_last(axi4buf_6_auto_out_w_bits_last),
    .auto_out_b_ready(axi4buf_6_auto_out_b_ready),
    .auto_out_b_valid(axi4buf_6_auto_out_b_valid),
    .auto_out_b_bits_id(axi4buf_6_auto_out_b_bits_id),
    .auto_out_b_bits_resp(axi4buf_6_auto_out_b_bits_resp),
    .auto_out_ar_ready(axi4buf_6_auto_out_ar_ready),
    .auto_out_ar_valid(axi4buf_6_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4buf_6_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4buf_6_auto_out_ar_bits_addr),
    .auto_out_ar_bits_size(axi4buf_6_auto_out_ar_bits_size),
    .auto_out_r_ready(axi4buf_6_auto_out_r_ready),
    .auto_out_r_valid(axi4buf_6_auto_out_r_valid),
    .auto_out_r_bits_id(axi4buf_6_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4buf_6_auto_out_r_bits_data),
    .auto_out_r_bits_resp(axi4buf_6_auto_out_r_bits_resp),
    .auto_out_r_bits_last(axi4buf_6_auto_out_r_bits_last)
  );
  AXI4Buffer axi4buf_7 ( // @[Buffer.scala 58:29]
    .clock(axi4buf_7_clock),
    .reset(axi4buf_7_reset),
    .auto_in_aw_ready(axi4buf_7_auto_in_aw_ready),
    .auto_in_aw_valid(axi4buf_7_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4buf_7_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4buf_7_auto_in_aw_bits_addr),
    .auto_in_aw_bits_size(axi4buf_7_auto_in_aw_bits_size),
    .auto_in_w_ready(axi4buf_7_auto_in_w_ready),
    .auto_in_w_valid(axi4buf_7_auto_in_w_valid),
    .auto_in_w_bits_data(axi4buf_7_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi4buf_7_auto_in_w_bits_strb),
    .auto_in_w_bits_last(axi4buf_7_auto_in_w_bits_last),
    .auto_in_b_ready(axi4buf_7_auto_in_b_ready),
    .auto_in_b_valid(axi4buf_7_auto_in_b_valid),
    .auto_in_b_bits_id(axi4buf_7_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi4buf_7_auto_in_b_bits_resp),
    .auto_in_ar_ready(axi4buf_7_auto_in_ar_ready),
    .auto_in_ar_valid(axi4buf_7_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4buf_7_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4buf_7_auto_in_ar_bits_addr),
    .auto_in_ar_bits_size(axi4buf_7_auto_in_ar_bits_size),
    .auto_in_r_ready(axi4buf_7_auto_in_r_ready),
    .auto_in_r_valid(axi4buf_7_auto_in_r_valid),
    .auto_in_r_bits_id(axi4buf_7_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4buf_7_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4buf_7_auto_in_r_bits_resp),
    .auto_in_r_bits_last(axi4buf_7_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4buf_7_auto_out_aw_ready),
    .auto_out_aw_valid(axi4buf_7_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4buf_7_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4buf_7_auto_out_aw_bits_addr),
    .auto_out_w_ready(axi4buf_7_auto_out_w_ready),
    .auto_out_w_valid(axi4buf_7_auto_out_w_valid),
    .auto_out_w_bits_data(axi4buf_7_auto_out_w_bits_data),
    .auto_out_w_bits_strb(axi4buf_7_auto_out_w_bits_strb),
    .auto_out_w_bits_last(axi4buf_7_auto_out_w_bits_last),
    .auto_out_b_ready(axi4buf_7_auto_out_b_ready),
    .auto_out_b_valid(axi4buf_7_auto_out_b_valid),
    .auto_out_b_bits_id(axi4buf_7_auto_out_b_bits_id),
    .auto_out_b_bits_resp(axi4buf_7_auto_out_b_bits_resp),
    .auto_out_ar_ready(axi4buf_7_auto_out_ar_ready),
    .auto_out_ar_valid(axi4buf_7_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4buf_7_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4buf_7_auto_out_ar_bits_addr),
    .auto_out_ar_bits_size(axi4buf_7_auto_out_ar_bits_size),
    .auto_out_r_ready(axi4buf_7_auto_out_r_ready),
    .auto_out_r_valid(axi4buf_7_auto_out_r_valid),
    .auto_out_r_bits_id(axi4buf_7_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4buf_7_auto_out_r_bits_data),
    .auto_out_r_bits_resp(axi4buf_7_auto_out_r_bits_resp),
    .auto_out_r_bits_last(axi4buf_7_auto_out_r_bits_last)
  );
  AXI4Buffer axi4buf_8 ( // @[Buffer.scala 58:29]
    .clock(axi4buf_8_clock),
    .reset(axi4buf_8_reset),
    .auto_in_aw_ready(axi4buf_8_auto_in_aw_ready),
    .auto_in_aw_valid(axi4buf_8_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4buf_8_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4buf_8_auto_in_aw_bits_addr),
    .auto_in_aw_bits_size(axi4buf_8_auto_in_aw_bits_size),
    .auto_in_w_ready(axi4buf_8_auto_in_w_ready),
    .auto_in_w_valid(axi4buf_8_auto_in_w_valid),
    .auto_in_w_bits_data(axi4buf_8_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi4buf_8_auto_in_w_bits_strb),
    .auto_in_w_bits_last(axi4buf_8_auto_in_w_bits_last),
    .auto_in_b_ready(axi4buf_8_auto_in_b_ready),
    .auto_in_b_valid(axi4buf_8_auto_in_b_valid),
    .auto_in_b_bits_id(axi4buf_8_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi4buf_8_auto_in_b_bits_resp),
    .auto_in_ar_ready(axi4buf_8_auto_in_ar_ready),
    .auto_in_ar_valid(axi4buf_8_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4buf_8_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4buf_8_auto_in_ar_bits_addr),
    .auto_in_ar_bits_size(axi4buf_8_auto_in_ar_bits_size),
    .auto_in_r_ready(axi4buf_8_auto_in_r_ready),
    .auto_in_r_valid(axi4buf_8_auto_in_r_valid),
    .auto_in_r_bits_id(axi4buf_8_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4buf_8_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4buf_8_auto_in_r_bits_resp),
    .auto_in_r_bits_last(axi4buf_8_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4buf_8_auto_out_aw_ready),
    .auto_out_aw_valid(axi4buf_8_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4buf_8_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4buf_8_auto_out_aw_bits_addr),
    .auto_out_w_ready(axi4buf_8_auto_out_w_ready),
    .auto_out_w_valid(axi4buf_8_auto_out_w_valid),
    .auto_out_w_bits_data(axi4buf_8_auto_out_w_bits_data),
    .auto_out_w_bits_strb(axi4buf_8_auto_out_w_bits_strb),
    .auto_out_w_bits_last(axi4buf_8_auto_out_w_bits_last),
    .auto_out_b_ready(axi4buf_8_auto_out_b_ready),
    .auto_out_b_valid(axi4buf_8_auto_out_b_valid),
    .auto_out_b_bits_id(axi4buf_8_auto_out_b_bits_id),
    .auto_out_b_bits_resp(axi4buf_8_auto_out_b_bits_resp),
    .auto_out_ar_ready(axi4buf_8_auto_out_ar_ready),
    .auto_out_ar_valid(axi4buf_8_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4buf_8_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4buf_8_auto_out_ar_bits_addr),
    .auto_out_ar_bits_size(axi4buf_8_auto_out_ar_bits_size),
    .auto_out_r_ready(axi4buf_8_auto_out_r_ready),
    .auto_out_r_valid(axi4buf_8_auto_out_r_valid),
    .auto_out_r_bits_id(axi4buf_8_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4buf_8_auto_out_r_bits_data),
    .auto_out_r_bits_resp(axi4buf_8_auto_out_r_bits_resp),
    .auto_out_r_bits_last(axi4buf_8_auto_out_r_bits_last)
  );
  AXI4Buffer axi4buf_9 ( // @[Buffer.scala 58:29]
    .clock(axi4buf_9_clock),
    .reset(axi4buf_9_reset),
    .auto_in_aw_ready(axi4buf_9_auto_in_aw_ready),
    .auto_in_aw_valid(axi4buf_9_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4buf_9_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4buf_9_auto_in_aw_bits_addr),
    .auto_in_aw_bits_size(axi4buf_9_auto_in_aw_bits_size),
    .auto_in_w_ready(axi4buf_9_auto_in_w_ready),
    .auto_in_w_valid(axi4buf_9_auto_in_w_valid),
    .auto_in_w_bits_data(axi4buf_9_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi4buf_9_auto_in_w_bits_strb),
    .auto_in_w_bits_last(axi4buf_9_auto_in_w_bits_last),
    .auto_in_b_ready(axi4buf_9_auto_in_b_ready),
    .auto_in_b_valid(axi4buf_9_auto_in_b_valid),
    .auto_in_b_bits_id(axi4buf_9_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi4buf_9_auto_in_b_bits_resp),
    .auto_in_ar_ready(axi4buf_9_auto_in_ar_ready),
    .auto_in_ar_valid(axi4buf_9_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4buf_9_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4buf_9_auto_in_ar_bits_addr),
    .auto_in_ar_bits_size(axi4buf_9_auto_in_ar_bits_size),
    .auto_in_r_ready(axi4buf_9_auto_in_r_ready),
    .auto_in_r_valid(axi4buf_9_auto_in_r_valid),
    .auto_in_r_bits_id(axi4buf_9_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4buf_9_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4buf_9_auto_in_r_bits_resp),
    .auto_in_r_bits_last(axi4buf_9_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4buf_9_auto_out_aw_ready),
    .auto_out_aw_valid(axi4buf_9_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4buf_9_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4buf_9_auto_out_aw_bits_addr),
    .auto_out_w_ready(axi4buf_9_auto_out_w_ready),
    .auto_out_w_valid(axi4buf_9_auto_out_w_valid),
    .auto_out_w_bits_data(axi4buf_9_auto_out_w_bits_data),
    .auto_out_w_bits_strb(axi4buf_9_auto_out_w_bits_strb),
    .auto_out_w_bits_last(axi4buf_9_auto_out_w_bits_last),
    .auto_out_b_ready(axi4buf_9_auto_out_b_ready),
    .auto_out_b_valid(axi4buf_9_auto_out_b_valid),
    .auto_out_b_bits_id(axi4buf_9_auto_out_b_bits_id),
    .auto_out_b_bits_resp(axi4buf_9_auto_out_b_bits_resp),
    .auto_out_ar_ready(axi4buf_9_auto_out_ar_ready),
    .auto_out_ar_valid(axi4buf_9_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4buf_9_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4buf_9_auto_out_ar_bits_addr),
    .auto_out_ar_bits_size(axi4buf_9_auto_out_ar_bits_size),
    .auto_out_r_ready(axi4buf_9_auto_out_r_ready),
    .auto_out_r_valid(axi4buf_9_auto_out_r_valid),
    .auto_out_r_bits_id(axi4buf_9_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4buf_9_auto_out_r_bits_data),
    .auto_out_r_bits_resp(axi4buf_9_auto_out_r_bits_resp),
    .auto_out_r_bits_last(axi4buf_9_auto_out_r_bits_last)
  );
  AXI4Buffer axi4buf_10 ( // @[Buffer.scala 58:29]
    .clock(axi4buf_10_clock),
    .reset(axi4buf_10_reset),
    .auto_in_aw_ready(axi4buf_10_auto_in_aw_ready),
    .auto_in_aw_valid(axi4buf_10_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4buf_10_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4buf_10_auto_in_aw_bits_addr),
    .auto_in_aw_bits_size(axi4buf_10_auto_in_aw_bits_size),
    .auto_in_w_ready(axi4buf_10_auto_in_w_ready),
    .auto_in_w_valid(axi4buf_10_auto_in_w_valid),
    .auto_in_w_bits_data(axi4buf_10_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi4buf_10_auto_in_w_bits_strb),
    .auto_in_w_bits_last(axi4buf_10_auto_in_w_bits_last),
    .auto_in_b_ready(axi4buf_10_auto_in_b_ready),
    .auto_in_b_valid(axi4buf_10_auto_in_b_valid),
    .auto_in_b_bits_id(axi4buf_10_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi4buf_10_auto_in_b_bits_resp),
    .auto_in_ar_ready(axi4buf_10_auto_in_ar_ready),
    .auto_in_ar_valid(axi4buf_10_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4buf_10_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4buf_10_auto_in_ar_bits_addr),
    .auto_in_ar_bits_size(axi4buf_10_auto_in_ar_bits_size),
    .auto_in_r_ready(axi4buf_10_auto_in_r_ready),
    .auto_in_r_valid(axi4buf_10_auto_in_r_valid),
    .auto_in_r_bits_id(axi4buf_10_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4buf_10_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4buf_10_auto_in_r_bits_resp),
    .auto_in_r_bits_last(axi4buf_10_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4buf_10_auto_out_aw_ready),
    .auto_out_aw_valid(axi4buf_10_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4buf_10_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4buf_10_auto_out_aw_bits_addr),
    .auto_out_w_ready(axi4buf_10_auto_out_w_ready),
    .auto_out_w_valid(axi4buf_10_auto_out_w_valid),
    .auto_out_w_bits_data(axi4buf_10_auto_out_w_bits_data),
    .auto_out_w_bits_strb(axi4buf_10_auto_out_w_bits_strb),
    .auto_out_w_bits_last(axi4buf_10_auto_out_w_bits_last),
    .auto_out_b_ready(axi4buf_10_auto_out_b_ready),
    .auto_out_b_valid(axi4buf_10_auto_out_b_valid),
    .auto_out_b_bits_id(axi4buf_10_auto_out_b_bits_id),
    .auto_out_b_bits_resp(axi4buf_10_auto_out_b_bits_resp),
    .auto_out_ar_ready(axi4buf_10_auto_out_ar_ready),
    .auto_out_ar_valid(axi4buf_10_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4buf_10_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4buf_10_auto_out_ar_bits_addr),
    .auto_out_ar_bits_size(axi4buf_10_auto_out_ar_bits_size),
    .auto_out_r_ready(axi4buf_10_auto_out_r_ready),
    .auto_out_r_valid(axi4buf_10_auto_out_r_valid),
    .auto_out_r_bits_id(axi4buf_10_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4buf_10_auto_out_r_bits_data),
    .auto_out_r_bits_resp(axi4buf_10_auto_out_r_bits_resp),
    .auto_out_r_bits_last(axi4buf_10_auto_out_r_bits_last)
  );
  AXI4Buffer axi4buf_11 ( // @[Buffer.scala 58:29]
    .clock(axi4buf_11_clock),
    .reset(axi4buf_11_reset),
    .auto_in_aw_ready(axi4buf_11_auto_in_aw_ready),
    .auto_in_aw_valid(axi4buf_11_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4buf_11_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4buf_11_auto_in_aw_bits_addr),
    .auto_in_aw_bits_size(axi4buf_11_auto_in_aw_bits_size),
    .auto_in_w_ready(axi4buf_11_auto_in_w_ready),
    .auto_in_w_valid(axi4buf_11_auto_in_w_valid),
    .auto_in_w_bits_data(axi4buf_11_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi4buf_11_auto_in_w_bits_strb),
    .auto_in_w_bits_last(axi4buf_11_auto_in_w_bits_last),
    .auto_in_b_ready(axi4buf_11_auto_in_b_ready),
    .auto_in_b_valid(axi4buf_11_auto_in_b_valid),
    .auto_in_b_bits_id(axi4buf_11_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi4buf_11_auto_in_b_bits_resp),
    .auto_in_ar_ready(axi4buf_11_auto_in_ar_ready),
    .auto_in_ar_valid(axi4buf_11_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4buf_11_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4buf_11_auto_in_ar_bits_addr),
    .auto_in_ar_bits_size(axi4buf_11_auto_in_ar_bits_size),
    .auto_in_r_ready(axi4buf_11_auto_in_r_ready),
    .auto_in_r_valid(axi4buf_11_auto_in_r_valid),
    .auto_in_r_bits_id(axi4buf_11_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4buf_11_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4buf_11_auto_in_r_bits_resp),
    .auto_in_r_bits_last(axi4buf_11_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4buf_11_auto_out_aw_ready),
    .auto_out_aw_valid(axi4buf_11_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4buf_11_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4buf_11_auto_out_aw_bits_addr),
    .auto_out_w_ready(axi4buf_11_auto_out_w_ready),
    .auto_out_w_valid(axi4buf_11_auto_out_w_valid),
    .auto_out_w_bits_data(axi4buf_11_auto_out_w_bits_data),
    .auto_out_w_bits_strb(axi4buf_11_auto_out_w_bits_strb),
    .auto_out_w_bits_last(axi4buf_11_auto_out_w_bits_last),
    .auto_out_b_ready(axi4buf_11_auto_out_b_ready),
    .auto_out_b_valid(axi4buf_11_auto_out_b_valid),
    .auto_out_b_bits_id(axi4buf_11_auto_out_b_bits_id),
    .auto_out_b_bits_resp(axi4buf_11_auto_out_b_bits_resp),
    .auto_out_ar_ready(axi4buf_11_auto_out_ar_ready),
    .auto_out_ar_valid(axi4buf_11_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4buf_11_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4buf_11_auto_out_ar_bits_addr),
    .auto_out_ar_bits_size(axi4buf_11_auto_out_ar_bits_size),
    .auto_out_r_ready(axi4buf_11_auto_out_r_ready),
    .auto_out_r_valid(axi4buf_11_auto_out_r_valid),
    .auto_out_r_bits_id(axi4buf_11_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4buf_11_auto_out_r_bits_data),
    .auto_out_r_bits_resp(axi4buf_11_auto_out_r_bits_resp),
    .auto_out_r_bits_last(axi4buf_11_auto_out_r_bits_last)
  );
  AXI4Buffer axi4buf_12 ( // @[Buffer.scala 58:29]
    .clock(axi4buf_12_clock),
    .reset(axi4buf_12_reset),
    .auto_in_aw_ready(axi4buf_12_auto_in_aw_ready),
    .auto_in_aw_valid(axi4buf_12_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4buf_12_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4buf_12_auto_in_aw_bits_addr),
    .auto_in_aw_bits_size(axi4buf_12_auto_in_aw_bits_size),
    .auto_in_w_ready(axi4buf_12_auto_in_w_ready),
    .auto_in_w_valid(axi4buf_12_auto_in_w_valid),
    .auto_in_w_bits_data(axi4buf_12_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi4buf_12_auto_in_w_bits_strb),
    .auto_in_w_bits_last(axi4buf_12_auto_in_w_bits_last),
    .auto_in_b_ready(axi4buf_12_auto_in_b_ready),
    .auto_in_b_valid(axi4buf_12_auto_in_b_valid),
    .auto_in_b_bits_id(axi4buf_12_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi4buf_12_auto_in_b_bits_resp),
    .auto_in_ar_ready(axi4buf_12_auto_in_ar_ready),
    .auto_in_ar_valid(axi4buf_12_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4buf_12_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4buf_12_auto_in_ar_bits_addr),
    .auto_in_ar_bits_size(axi4buf_12_auto_in_ar_bits_size),
    .auto_in_r_ready(axi4buf_12_auto_in_r_ready),
    .auto_in_r_valid(axi4buf_12_auto_in_r_valid),
    .auto_in_r_bits_id(axi4buf_12_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4buf_12_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4buf_12_auto_in_r_bits_resp),
    .auto_in_r_bits_last(axi4buf_12_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4buf_12_auto_out_aw_ready),
    .auto_out_aw_valid(axi4buf_12_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4buf_12_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4buf_12_auto_out_aw_bits_addr),
    .auto_out_w_ready(axi4buf_12_auto_out_w_ready),
    .auto_out_w_valid(axi4buf_12_auto_out_w_valid),
    .auto_out_w_bits_data(axi4buf_12_auto_out_w_bits_data),
    .auto_out_w_bits_strb(axi4buf_12_auto_out_w_bits_strb),
    .auto_out_w_bits_last(axi4buf_12_auto_out_w_bits_last),
    .auto_out_b_ready(axi4buf_12_auto_out_b_ready),
    .auto_out_b_valid(axi4buf_12_auto_out_b_valid),
    .auto_out_b_bits_id(axi4buf_12_auto_out_b_bits_id),
    .auto_out_b_bits_resp(axi4buf_12_auto_out_b_bits_resp),
    .auto_out_ar_ready(axi4buf_12_auto_out_ar_ready),
    .auto_out_ar_valid(axi4buf_12_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4buf_12_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4buf_12_auto_out_ar_bits_addr),
    .auto_out_ar_bits_size(axi4buf_12_auto_out_ar_bits_size),
    .auto_out_r_ready(axi4buf_12_auto_out_r_ready),
    .auto_out_r_valid(axi4buf_12_auto_out_r_valid),
    .auto_out_r_bits_id(axi4buf_12_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4buf_12_auto_out_r_bits_data),
    .auto_out_r_bits_resp(axi4buf_12_auto_out_r_bits_resp),
    .auto_out_r_bits_last(axi4buf_12_auto_out_r_bits_last)
  );
  AXI4Buffer axi4buf_13 ( // @[Buffer.scala 58:29]
    .clock(axi4buf_13_clock),
    .reset(axi4buf_13_reset),
    .auto_in_aw_ready(axi4buf_13_auto_in_aw_ready),
    .auto_in_aw_valid(axi4buf_13_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4buf_13_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4buf_13_auto_in_aw_bits_addr),
    .auto_in_aw_bits_size(axi4buf_13_auto_in_aw_bits_size),
    .auto_in_w_ready(axi4buf_13_auto_in_w_ready),
    .auto_in_w_valid(axi4buf_13_auto_in_w_valid),
    .auto_in_w_bits_data(axi4buf_13_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi4buf_13_auto_in_w_bits_strb),
    .auto_in_w_bits_last(axi4buf_13_auto_in_w_bits_last),
    .auto_in_b_ready(axi4buf_13_auto_in_b_ready),
    .auto_in_b_valid(axi4buf_13_auto_in_b_valid),
    .auto_in_b_bits_id(axi4buf_13_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi4buf_13_auto_in_b_bits_resp),
    .auto_in_ar_ready(axi4buf_13_auto_in_ar_ready),
    .auto_in_ar_valid(axi4buf_13_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4buf_13_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4buf_13_auto_in_ar_bits_addr),
    .auto_in_ar_bits_size(axi4buf_13_auto_in_ar_bits_size),
    .auto_in_r_ready(axi4buf_13_auto_in_r_ready),
    .auto_in_r_valid(axi4buf_13_auto_in_r_valid),
    .auto_in_r_bits_id(axi4buf_13_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4buf_13_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4buf_13_auto_in_r_bits_resp),
    .auto_in_r_bits_last(axi4buf_13_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4buf_13_auto_out_aw_ready),
    .auto_out_aw_valid(axi4buf_13_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4buf_13_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4buf_13_auto_out_aw_bits_addr),
    .auto_out_w_ready(axi4buf_13_auto_out_w_ready),
    .auto_out_w_valid(axi4buf_13_auto_out_w_valid),
    .auto_out_w_bits_data(axi4buf_13_auto_out_w_bits_data),
    .auto_out_w_bits_strb(axi4buf_13_auto_out_w_bits_strb),
    .auto_out_w_bits_last(axi4buf_13_auto_out_w_bits_last),
    .auto_out_b_ready(axi4buf_13_auto_out_b_ready),
    .auto_out_b_valid(axi4buf_13_auto_out_b_valid),
    .auto_out_b_bits_id(axi4buf_13_auto_out_b_bits_id),
    .auto_out_b_bits_resp(axi4buf_13_auto_out_b_bits_resp),
    .auto_out_ar_ready(axi4buf_13_auto_out_ar_ready),
    .auto_out_ar_valid(axi4buf_13_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4buf_13_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4buf_13_auto_out_ar_bits_addr),
    .auto_out_ar_bits_size(axi4buf_13_auto_out_ar_bits_size),
    .auto_out_r_ready(axi4buf_13_auto_out_r_ready),
    .auto_out_r_valid(axi4buf_13_auto_out_r_valid),
    .auto_out_r_bits_id(axi4buf_13_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4buf_13_auto_out_r_bits_data),
    .auto_out_r_bits_resp(axi4buf_13_auto_out_r_bits_resp),
    .auto_out_r_bits_last(axi4buf_13_auto_out_r_bits_last)
  );
  AXI4Buffer axi4buf_14 ( // @[Buffer.scala 58:29]
    .clock(axi4buf_14_clock),
    .reset(axi4buf_14_reset),
    .auto_in_aw_ready(axi4buf_14_auto_in_aw_ready),
    .auto_in_aw_valid(axi4buf_14_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4buf_14_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4buf_14_auto_in_aw_bits_addr),
    .auto_in_aw_bits_size(axi4buf_14_auto_in_aw_bits_size),
    .auto_in_w_ready(axi4buf_14_auto_in_w_ready),
    .auto_in_w_valid(axi4buf_14_auto_in_w_valid),
    .auto_in_w_bits_data(axi4buf_14_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi4buf_14_auto_in_w_bits_strb),
    .auto_in_w_bits_last(axi4buf_14_auto_in_w_bits_last),
    .auto_in_b_ready(axi4buf_14_auto_in_b_ready),
    .auto_in_b_valid(axi4buf_14_auto_in_b_valid),
    .auto_in_b_bits_id(axi4buf_14_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi4buf_14_auto_in_b_bits_resp),
    .auto_in_ar_ready(axi4buf_14_auto_in_ar_ready),
    .auto_in_ar_valid(axi4buf_14_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4buf_14_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4buf_14_auto_in_ar_bits_addr),
    .auto_in_ar_bits_size(axi4buf_14_auto_in_ar_bits_size),
    .auto_in_r_ready(axi4buf_14_auto_in_r_ready),
    .auto_in_r_valid(axi4buf_14_auto_in_r_valid),
    .auto_in_r_bits_id(axi4buf_14_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4buf_14_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4buf_14_auto_in_r_bits_resp),
    .auto_in_r_bits_last(axi4buf_14_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4buf_14_auto_out_aw_ready),
    .auto_out_aw_valid(axi4buf_14_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4buf_14_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4buf_14_auto_out_aw_bits_addr),
    .auto_out_w_ready(axi4buf_14_auto_out_w_ready),
    .auto_out_w_valid(axi4buf_14_auto_out_w_valid),
    .auto_out_w_bits_data(axi4buf_14_auto_out_w_bits_data),
    .auto_out_w_bits_strb(axi4buf_14_auto_out_w_bits_strb),
    .auto_out_w_bits_last(axi4buf_14_auto_out_w_bits_last),
    .auto_out_b_ready(axi4buf_14_auto_out_b_ready),
    .auto_out_b_valid(axi4buf_14_auto_out_b_valid),
    .auto_out_b_bits_id(axi4buf_14_auto_out_b_bits_id),
    .auto_out_b_bits_resp(axi4buf_14_auto_out_b_bits_resp),
    .auto_out_ar_ready(axi4buf_14_auto_out_ar_ready),
    .auto_out_ar_valid(axi4buf_14_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4buf_14_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4buf_14_auto_out_ar_bits_addr),
    .auto_out_ar_bits_size(axi4buf_14_auto_out_ar_bits_size),
    .auto_out_r_ready(axi4buf_14_auto_out_r_ready),
    .auto_out_r_valid(axi4buf_14_auto_out_r_valid),
    .auto_out_r_bits_id(axi4buf_14_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4buf_14_auto_out_r_bits_data),
    .auto_out_r_bits_resp(axi4buf_14_auto_out_r_bits_resp),
    .auto_out_r_bits_last(axi4buf_14_auto_out_r_bits_last)
  );
  AXI4Buffer axi4buf_15 ( // @[Buffer.scala 58:29]
    .clock(axi4buf_15_clock),
    .reset(axi4buf_15_reset),
    .auto_in_aw_ready(axi4buf_15_auto_in_aw_ready),
    .auto_in_aw_valid(axi4buf_15_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4buf_15_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4buf_15_auto_in_aw_bits_addr),
    .auto_in_aw_bits_size(axi4buf_15_auto_in_aw_bits_size),
    .auto_in_w_ready(axi4buf_15_auto_in_w_ready),
    .auto_in_w_valid(axi4buf_15_auto_in_w_valid),
    .auto_in_w_bits_data(axi4buf_15_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi4buf_15_auto_in_w_bits_strb),
    .auto_in_w_bits_last(axi4buf_15_auto_in_w_bits_last),
    .auto_in_b_ready(axi4buf_15_auto_in_b_ready),
    .auto_in_b_valid(axi4buf_15_auto_in_b_valid),
    .auto_in_b_bits_id(axi4buf_15_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi4buf_15_auto_in_b_bits_resp),
    .auto_in_ar_ready(axi4buf_15_auto_in_ar_ready),
    .auto_in_ar_valid(axi4buf_15_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4buf_15_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4buf_15_auto_in_ar_bits_addr),
    .auto_in_ar_bits_size(axi4buf_15_auto_in_ar_bits_size),
    .auto_in_r_ready(axi4buf_15_auto_in_r_ready),
    .auto_in_r_valid(axi4buf_15_auto_in_r_valid),
    .auto_in_r_bits_id(axi4buf_15_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4buf_15_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4buf_15_auto_in_r_bits_resp),
    .auto_in_r_bits_last(axi4buf_15_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4buf_15_auto_out_aw_ready),
    .auto_out_aw_valid(axi4buf_15_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4buf_15_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4buf_15_auto_out_aw_bits_addr),
    .auto_out_w_ready(axi4buf_15_auto_out_w_ready),
    .auto_out_w_valid(axi4buf_15_auto_out_w_valid),
    .auto_out_w_bits_data(axi4buf_15_auto_out_w_bits_data),
    .auto_out_w_bits_strb(axi4buf_15_auto_out_w_bits_strb),
    .auto_out_w_bits_last(axi4buf_15_auto_out_w_bits_last),
    .auto_out_b_ready(axi4buf_15_auto_out_b_ready),
    .auto_out_b_valid(axi4buf_15_auto_out_b_valid),
    .auto_out_b_bits_id(axi4buf_15_auto_out_b_bits_id),
    .auto_out_b_bits_resp(axi4buf_15_auto_out_b_bits_resp),
    .auto_out_ar_ready(axi4buf_15_auto_out_ar_ready),
    .auto_out_ar_valid(axi4buf_15_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4buf_15_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4buf_15_auto_out_ar_bits_addr),
    .auto_out_ar_bits_size(axi4buf_15_auto_out_ar_bits_size),
    .auto_out_r_ready(axi4buf_15_auto_out_r_ready),
    .auto_out_r_valid(axi4buf_15_auto_out_r_valid),
    .auto_out_r_bits_id(axi4buf_15_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4buf_15_auto_out_r_bits_data),
    .auto_out_r_bits_resp(axi4buf_15_auto_out_r_bits_resp),
    .auto_out_r_bits_last(axi4buf_15_auto_out_r_bits_last)
  );
  AXI4Buffer axi4buf_16 ( // @[Buffer.scala 58:29]
    .clock(axi4buf_16_clock),
    .reset(axi4buf_16_reset),
    .auto_in_aw_ready(axi4buf_16_auto_in_aw_ready),
    .auto_in_aw_valid(axi4buf_16_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4buf_16_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4buf_16_auto_in_aw_bits_addr),
    .auto_in_aw_bits_size(axi4buf_16_auto_in_aw_bits_size),
    .auto_in_w_ready(axi4buf_16_auto_in_w_ready),
    .auto_in_w_valid(axi4buf_16_auto_in_w_valid),
    .auto_in_w_bits_data(axi4buf_16_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi4buf_16_auto_in_w_bits_strb),
    .auto_in_w_bits_last(axi4buf_16_auto_in_w_bits_last),
    .auto_in_b_ready(axi4buf_16_auto_in_b_ready),
    .auto_in_b_valid(axi4buf_16_auto_in_b_valid),
    .auto_in_b_bits_id(axi4buf_16_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi4buf_16_auto_in_b_bits_resp),
    .auto_in_ar_ready(axi4buf_16_auto_in_ar_ready),
    .auto_in_ar_valid(axi4buf_16_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4buf_16_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4buf_16_auto_in_ar_bits_addr),
    .auto_in_ar_bits_size(axi4buf_16_auto_in_ar_bits_size),
    .auto_in_r_ready(axi4buf_16_auto_in_r_ready),
    .auto_in_r_valid(axi4buf_16_auto_in_r_valid),
    .auto_in_r_bits_id(axi4buf_16_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4buf_16_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4buf_16_auto_in_r_bits_resp),
    .auto_in_r_bits_last(axi4buf_16_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4buf_16_auto_out_aw_ready),
    .auto_out_aw_valid(axi4buf_16_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4buf_16_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4buf_16_auto_out_aw_bits_addr),
    .auto_out_w_ready(axi4buf_16_auto_out_w_ready),
    .auto_out_w_valid(axi4buf_16_auto_out_w_valid),
    .auto_out_w_bits_data(axi4buf_16_auto_out_w_bits_data),
    .auto_out_w_bits_strb(axi4buf_16_auto_out_w_bits_strb),
    .auto_out_w_bits_last(axi4buf_16_auto_out_w_bits_last),
    .auto_out_b_ready(axi4buf_16_auto_out_b_ready),
    .auto_out_b_valid(axi4buf_16_auto_out_b_valid),
    .auto_out_b_bits_id(axi4buf_16_auto_out_b_bits_id),
    .auto_out_b_bits_resp(axi4buf_16_auto_out_b_bits_resp),
    .auto_out_ar_ready(axi4buf_16_auto_out_ar_ready),
    .auto_out_ar_valid(axi4buf_16_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4buf_16_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4buf_16_auto_out_ar_bits_addr),
    .auto_out_ar_bits_size(axi4buf_16_auto_out_ar_bits_size),
    .auto_out_r_ready(axi4buf_16_auto_out_r_ready),
    .auto_out_r_valid(axi4buf_16_auto_out_r_valid),
    .auto_out_r_bits_id(axi4buf_16_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4buf_16_auto_out_r_bits_data),
    .auto_out_r_bits_resp(axi4buf_16_auto_out_r_bits_resp),
    .auto_out_r_bits_last(axi4buf_16_auto_out_r_bits_last)
  );
  AXI4Buffer axi4buf_17 ( // @[Buffer.scala 58:29]
    .clock(axi4buf_17_clock),
    .reset(axi4buf_17_reset),
    .auto_in_aw_ready(axi4buf_17_auto_in_aw_ready),
    .auto_in_aw_valid(axi4buf_17_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4buf_17_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4buf_17_auto_in_aw_bits_addr),
    .auto_in_aw_bits_size(axi4buf_17_auto_in_aw_bits_size),
    .auto_in_w_ready(axi4buf_17_auto_in_w_ready),
    .auto_in_w_valid(axi4buf_17_auto_in_w_valid),
    .auto_in_w_bits_data(axi4buf_17_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi4buf_17_auto_in_w_bits_strb),
    .auto_in_w_bits_last(axi4buf_17_auto_in_w_bits_last),
    .auto_in_b_ready(axi4buf_17_auto_in_b_ready),
    .auto_in_b_valid(axi4buf_17_auto_in_b_valid),
    .auto_in_b_bits_id(axi4buf_17_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi4buf_17_auto_in_b_bits_resp),
    .auto_in_ar_ready(axi4buf_17_auto_in_ar_ready),
    .auto_in_ar_valid(axi4buf_17_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4buf_17_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4buf_17_auto_in_ar_bits_addr),
    .auto_in_ar_bits_size(axi4buf_17_auto_in_ar_bits_size),
    .auto_in_r_ready(axi4buf_17_auto_in_r_ready),
    .auto_in_r_valid(axi4buf_17_auto_in_r_valid),
    .auto_in_r_bits_id(axi4buf_17_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4buf_17_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4buf_17_auto_in_r_bits_resp),
    .auto_in_r_bits_last(axi4buf_17_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4buf_17_auto_out_aw_ready),
    .auto_out_aw_valid(axi4buf_17_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4buf_17_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4buf_17_auto_out_aw_bits_addr),
    .auto_out_w_ready(axi4buf_17_auto_out_w_ready),
    .auto_out_w_valid(axi4buf_17_auto_out_w_valid),
    .auto_out_w_bits_data(axi4buf_17_auto_out_w_bits_data),
    .auto_out_w_bits_strb(axi4buf_17_auto_out_w_bits_strb),
    .auto_out_w_bits_last(axi4buf_17_auto_out_w_bits_last),
    .auto_out_b_ready(axi4buf_17_auto_out_b_ready),
    .auto_out_b_valid(axi4buf_17_auto_out_b_valid),
    .auto_out_b_bits_id(axi4buf_17_auto_out_b_bits_id),
    .auto_out_b_bits_resp(axi4buf_17_auto_out_b_bits_resp),
    .auto_out_ar_ready(axi4buf_17_auto_out_ar_ready),
    .auto_out_ar_valid(axi4buf_17_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4buf_17_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4buf_17_auto_out_ar_bits_addr),
    .auto_out_ar_bits_size(axi4buf_17_auto_out_ar_bits_size),
    .auto_out_r_ready(axi4buf_17_auto_out_r_ready),
    .auto_out_r_valid(axi4buf_17_auto_out_r_valid),
    .auto_out_r_bits_id(axi4buf_17_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4buf_17_auto_out_r_bits_data),
    .auto_out_r_bits_resp(axi4buf_17_auto_out_r_bits_resp),
    .auto_out_r_bits_last(axi4buf_17_auto_out_r_bits_last)
  );
  AXI4Buffer axi4buf_18 ( // @[Buffer.scala 58:29]
    .clock(axi4buf_18_clock),
    .reset(axi4buf_18_reset),
    .auto_in_aw_ready(axi4buf_18_auto_in_aw_ready),
    .auto_in_aw_valid(axi4buf_18_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4buf_18_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4buf_18_auto_in_aw_bits_addr),
    .auto_in_aw_bits_size(axi4buf_18_auto_in_aw_bits_size),
    .auto_in_w_ready(axi4buf_18_auto_in_w_ready),
    .auto_in_w_valid(axi4buf_18_auto_in_w_valid),
    .auto_in_w_bits_data(axi4buf_18_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi4buf_18_auto_in_w_bits_strb),
    .auto_in_w_bits_last(axi4buf_18_auto_in_w_bits_last),
    .auto_in_b_ready(axi4buf_18_auto_in_b_ready),
    .auto_in_b_valid(axi4buf_18_auto_in_b_valid),
    .auto_in_b_bits_id(axi4buf_18_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi4buf_18_auto_in_b_bits_resp),
    .auto_in_ar_ready(axi4buf_18_auto_in_ar_ready),
    .auto_in_ar_valid(axi4buf_18_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4buf_18_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4buf_18_auto_in_ar_bits_addr),
    .auto_in_ar_bits_size(axi4buf_18_auto_in_ar_bits_size),
    .auto_in_r_ready(axi4buf_18_auto_in_r_ready),
    .auto_in_r_valid(axi4buf_18_auto_in_r_valid),
    .auto_in_r_bits_id(axi4buf_18_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4buf_18_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4buf_18_auto_in_r_bits_resp),
    .auto_in_r_bits_last(axi4buf_18_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4buf_18_auto_out_aw_ready),
    .auto_out_aw_valid(axi4buf_18_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4buf_18_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4buf_18_auto_out_aw_bits_addr),
    .auto_out_w_ready(axi4buf_18_auto_out_w_ready),
    .auto_out_w_valid(axi4buf_18_auto_out_w_valid),
    .auto_out_w_bits_data(axi4buf_18_auto_out_w_bits_data),
    .auto_out_w_bits_strb(axi4buf_18_auto_out_w_bits_strb),
    .auto_out_w_bits_last(axi4buf_18_auto_out_w_bits_last),
    .auto_out_b_ready(axi4buf_18_auto_out_b_ready),
    .auto_out_b_valid(axi4buf_18_auto_out_b_valid),
    .auto_out_b_bits_id(axi4buf_18_auto_out_b_bits_id),
    .auto_out_b_bits_resp(axi4buf_18_auto_out_b_bits_resp),
    .auto_out_ar_ready(axi4buf_18_auto_out_ar_ready),
    .auto_out_ar_valid(axi4buf_18_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4buf_18_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4buf_18_auto_out_ar_bits_addr),
    .auto_out_ar_bits_size(axi4buf_18_auto_out_ar_bits_size),
    .auto_out_r_ready(axi4buf_18_auto_out_r_ready),
    .auto_out_r_valid(axi4buf_18_auto_out_r_valid),
    .auto_out_r_bits_id(axi4buf_18_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4buf_18_auto_out_r_bits_data),
    .auto_out_r_bits_resp(axi4buf_18_auto_out_r_bits_resp),
    .auto_out_r_bits_last(axi4buf_18_auto_out_r_bits_last)
  );
  AXI4Buffer axi4buf_19 ( // @[Buffer.scala 58:29]
    .clock(axi4buf_19_clock),
    .reset(axi4buf_19_reset),
    .auto_in_aw_ready(axi4buf_19_auto_in_aw_ready),
    .auto_in_aw_valid(axi4buf_19_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4buf_19_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4buf_19_auto_in_aw_bits_addr),
    .auto_in_aw_bits_size(axi4buf_19_auto_in_aw_bits_size),
    .auto_in_w_ready(axi4buf_19_auto_in_w_ready),
    .auto_in_w_valid(axi4buf_19_auto_in_w_valid),
    .auto_in_w_bits_data(axi4buf_19_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi4buf_19_auto_in_w_bits_strb),
    .auto_in_w_bits_last(axi4buf_19_auto_in_w_bits_last),
    .auto_in_b_ready(axi4buf_19_auto_in_b_ready),
    .auto_in_b_valid(axi4buf_19_auto_in_b_valid),
    .auto_in_b_bits_id(axi4buf_19_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi4buf_19_auto_in_b_bits_resp),
    .auto_in_ar_ready(axi4buf_19_auto_in_ar_ready),
    .auto_in_ar_valid(axi4buf_19_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4buf_19_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4buf_19_auto_in_ar_bits_addr),
    .auto_in_ar_bits_size(axi4buf_19_auto_in_ar_bits_size),
    .auto_in_r_ready(axi4buf_19_auto_in_r_ready),
    .auto_in_r_valid(axi4buf_19_auto_in_r_valid),
    .auto_in_r_bits_id(axi4buf_19_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4buf_19_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4buf_19_auto_in_r_bits_resp),
    .auto_in_r_bits_last(axi4buf_19_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4buf_19_auto_out_aw_ready),
    .auto_out_aw_valid(axi4buf_19_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4buf_19_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4buf_19_auto_out_aw_bits_addr),
    .auto_out_w_ready(axi4buf_19_auto_out_w_ready),
    .auto_out_w_valid(axi4buf_19_auto_out_w_valid),
    .auto_out_w_bits_data(axi4buf_19_auto_out_w_bits_data),
    .auto_out_w_bits_strb(axi4buf_19_auto_out_w_bits_strb),
    .auto_out_w_bits_last(axi4buf_19_auto_out_w_bits_last),
    .auto_out_b_ready(axi4buf_19_auto_out_b_ready),
    .auto_out_b_valid(axi4buf_19_auto_out_b_valid),
    .auto_out_b_bits_id(axi4buf_19_auto_out_b_bits_id),
    .auto_out_b_bits_resp(axi4buf_19_auto_out_b_bits_resp),
    .auto_out_ar_ready(axi4buf_19_auto_out_ar_ready),
    .auto_out_ar_valid(axi4buf_19_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4buf_19_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4buf_19_auto_out_ar_bits_addr),
    .auto_out_ar_bits_size(axi4buf_19_auto_out_ar_bits_size),
    .auto_out_r_ready(axi4buf_19_auto_out_r_ready),
    .auto_out_r_valid(axi4buf_19_auto_out_r_valid),
    .auto_out_r_bits_id(axi4buf_19_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4buf_19_auto_out_r_bits_data),
    .auto_out_r_bits_resp(axi4buf_19_auto_out_r_bits_resp),
    .auto_out_r_bits_last(axi4buf_19_auto_out_r_bits_last)
  );
  AXI4Buffer axi4buf_20 ( // @[Buffer.scala 58:29]
    .clock(axi4buf_20_clock),
    .reset(axi4buf_20_reset),
    .auto_in_aw_ready(axi4buf_20_auto_in_aw_ready),
    .auto_in_aw_valid(axi4buf_20_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4buf_20_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4buf_20_auto_in_aw_bits_addr),
    .auto_in_aw_bits_size(axi4buf_20_auto_in_aw_bits_size),
    .auto_in_w_ready(axi4buf_20_auto_in_w_ready),
    .auto_in_w_valid(axi4buf_20_auto_in_w_valid),
    .auto_in_w_bits_data(axi4buf_20_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi4buf_20_auto_in_w_bits_strb),
    .auto_in_w_bits_last(axi4buf_20_auto_in_w_bits_last),
    .auto_in_b_ready(axi4buf_20_auto_in_b_ready),
    .auto_in_b_valid(axi4buf_20_auto_in_b_valid),
    .auto_in_b_bits_id(axi4buf_20_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi4buf_20_auto_in_b_bits_resp),
    .auto_in_ar_ready(axi4buf_20_auto_in_ar_ready),
    .auto_in_ar_valid(axi4buf_20_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4buf_20_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4buf_20_auto_in_ar_bits_addr),
    .auto_in_ar_bits_size(axi4buf_20_auto_in_ar_bits_size),
    .auto_in_r_ready(axi4buf_20_auto_in_r_ready),
    .auto_in_r_valid(axi4buf_20_auto_in_r_valid),
    .auto_in_r_bits_id(axi4buf_20_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4buf_20_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4buf_20_auto_in_r_bits_resp),
    .auto_in_r_bits_last(axi4buf_20_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4buf_20_auto_out_aw_ready),
    .auto_out_aw_valid(axi4buf_20_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4buf_20_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4buf_20_auto_out_aw_bits_addr),
    .auto_out_w_ready(axi4buf_20_auto_out_w_ready),
    .auto_out_w_valid(axi4buf_20_auto_out_w_valid),
    .auto_out_w_bits_data(axi4buf_20_auto_out_w_bits_data),
    .auto_out_w_bits_strb(axi4buf_20_auto_out_w_bits_strb),
    .auto_out_w_bits_last(axi4buf_20_auto_out_w_bits_last),
    .auto_out_b_ready(axi4buf_20_auto_out_b_ready),
    .auto_out_b_valid(axi4buf_20_auto_out_b_valid),
    .auto_out_b_bits_id(axi4buf_20_auto_out_b_bits_id),
    .auto_out_b_bits_resp(axi4buf_20_auto_out_b_bits_resp),
    .auto_out_ar_ready(axi4buf_20_auto_out_ar_ready),
    .auto_out_ar_valid(axi4buf_20_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4buf_20_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4buf_20_auto_out_ar_bits_addr),
    .auto_out_ar_bits_size(axi4buf_20_auto_out_ar_bits_size),
    .auto_out_r_ready(axi4buf_20_auto_out_r_ready),
    .auto_out_r_valid(axi4buf_20_auto_out_r_valid),
    .auto_out_r_bits_id(axi4buf_20_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4buf_20_auto_out_r_bits_data),
    .auto_out_r_bits_resp(axi4buf_20_auto_out_r_bits_resp),
    .auto_out_r_bits_last(axi4buf_20_auto_out_r_bits_last)
  );
  AXI4StreamBuffer buffer ( // @[Buffer.scala 29:28]
    .clock(buffer_clock),
    .reset(buffer_reset),
    .auto_in_ready(buffer_auto_in_ready),
    .auto_in_valid(buffer_auto_in_valid),
    .auto_in_bits_data(buffer_auto_in_bits_data),
    .auto_in_bits_last(buffer_auto_in_bits_last),
    .auto_out_ready(buffer_auto_out_ready),
    .auto_out_valid(buffer_auto_out_valid),
    .auto_out_bits_data(buffer_auto_out_bits_data),
    .auto_out_bits_last(buffer_auto_out_bits_last)
  );
  AXI4StreamBuffer_1 buffer_1 ( // @[Buffer.scala 29:28]
    .clock(buffer_1_clock),
    .reset(buffer_1_reset),
    .auto_in_ready(buffer_1_auto_in_ready),
    .auto_in_valid(buffer_1_auto_in_valid),
    .auto_in_bits_data(buffer_1_auto_in_bits_data),
    .auto_in_bits_last(buffer_1_auto_in_bits_last),
    .auto_out_ready(buffer_1_auto_out_ready),
    .auto_out_valid(buffer_1_auto_out_valid),
    .auto_out_bits_data(buffer_1_auto_out_bits_data),
    .auto_out_bits_last(buffer_1_auto_out_bits_last)
  );
  AXI4StreamBuffer_2 buffer_2 ( // @[Buffer.scala 29:28]
    .clock(buffer_2_clock),
    .reset(buffer_2_reset),
    .auto_in_ready(buffer_2_auto_in_ready),
    .auto_in_valid(buffer_2_auto_in_valid),
    .auto_in_bits_data(buffer_2_auto_in_bits_data),
    .auto_in_bits_last(buffer_2_auto_in_bits_last),
    .auto_out_ready(buffer_2_auto_out_ready),
    .auto_out_valid(buffer_2_auto_out_valid),
    .auto_out_bits_data(buffer_2_auto_out_bits_data),
    .auto_out_bits_last(buffer_2_auto_out_bits_last)
  );
  AXI4StreamBuffer_1 buffer_3 ( // @[Buffer.scala 29:28]
    .clock(buffer_3_clock),
    .reset(buffer_3_reset),
    .auto_in_ready(buffer_3_auto_in_ready),
    .auto_in_valid(buffer_3_auto_in_valid),
    .auto_in_bits_data(buffer_3_auto_in_bits_data),
    .auto_in_bits_last(buffer_3_auto_in_bits_last),
    .auto_out_ready(buffer_3_auto_out_ready),
    .auto_out_valid(buffer_3_auto_out_valid),
    .auto_out_bits_data(buffer_3_auto_out_bits_data),
    .auto_out_bits_last(buffer_3_auto_out_bits_last)
  );
  AXI4StreamBuffer_4 buffer_4 ( // @[Buffer.scala 29:28]
    .clock(buffer_4_clock),
    .reset(buffer_4_reset),
    .auto_in_ready(buffer_4_auto_in_ready),
    .auto_in_valid(buffer_4_auto_in_valid),
    .auto_in_bits_data(buffer_4_auto_in_bits_data),
    .auto_in_bits_last(buffer_4_auto_in_bits_last),
    .auto_out_ready(buffer_4_auto_out_ready),
    .auto_out_valid(buffer_4_auto_out_valid),
    .auto_out_bits_data(buffer_4_auto_out_bits_data),
    .auto_out_bits_last(buffer_4_auto_out_bits_last)
  );
  AXI4StreamBuffer_5 buffer_5 ( // @[Buffer.scala 29:28]
    .clock(buffer_5_clock),
    .reset(buffer_5_reset),
    .auto_in_ready(buffer_5_auto_in_ready),
    .auto_in_valid(buffer_5_auto_in_valid),
    .auto_in_bits_data(buffer_5_auto_in_bits_data),
    .auto_in_bits_last(buffer_5_auto_in_bits_last),
    .auto_out_ready(buffer_5_auto_out_ready),
    .auto_out_valid(buffer_5_auto_out_valid),
    .auto_out_bits_data(buffer_5_auto_out_bits_data),
    .auto_out_bits_last(buffer_5_auto_out_bits_last)
  );
  AXI4StreamBuffer_5 buffer_6 ( // @[Buffer.scala 29:28]
    .clock(buffer_6_clock),
    .reset(buffer_6_reset),
    .auto_in_ready(buffer_6_auto_in_ready),
    .auto_in_valid(buffer_6_auto_in_valid),
    .auto_in_bits_data(buffer_6_auto_in_bits_data),
    .auto_in_bits_last(buffer_6_auto_in_bits_last),
    .auto_out_ready(buffer_6_auto_out_ready),
    .auto_out_valid(buffer_6_auto_out_valid),
    .auto_out_bits_data(buffer_6_auto_out_bits_data),
    .auto_out_bits_last(buffer_6_auto_out_bits_last)
  );
  AXI4StreamBuffer_5 buffer_7 ( // @[Buffer.scala 29:28]
    .clock(buffer_7_clock),
    .reset(buffer_7_reset),
    .auto_in_ready(buffer_7_auto_in_ready),
    .auto_in_valid(buffer_7_auto_in_valid),
    .auto_in_bits_data(buffer_7_auto_in_bits_data),
    .auto_in_bits_last(buffer_7_auto_in_bits_last),
    .auto_out_ready(buffer_7_auto_out_ready),
    .auto_out_valid(buffer_7_auto_out_valid),
    .auto_out_bits_data(buffer_7_auto_out_bits_data),
    .auto_out_bits_last(buffer_7_auto_out_bits_last)
  );
  AXI4StreamBuffer_5 buffer_8 ( // @[Buffer.scala 29:28]
    .clock(buffer_8_clock),
    .reset(buffer_8_reset),
    .auto_in_ready(buffer_8_auto_in_ready),
    .auto_in_valid(buffer_8_auto_in_valid),
    .auto_in_bits_data(buffer_8_auto_in_bits_data),
    .auto_in_bits_last(buffer_8_auto_in_bits_last),
    .auto_out_ready(buffer_8_auto_out_ready),
    .auto_out_valid(buffer_8_auto_out_valid),
    .auto_out_bits_data(buffer_8_auto_out_bits_data),
    .auto_out_bits_last(buffer_8_auto_out_bits_last)
  );
  AXI4StreamBuffer_9 buffer_9 ( // @[Buffer.scala 29:28]
    .clock(buffer_9_clock),
    .reset(buffer_9_reset),
    .auto_in_ready(buffer_9_auto_in_ready),
    .auto_in_valid(buffer_9_auto_in_valid),
    .auto_in_bits_data(buffer_9_auto_in_bits_data),
    .auto_in_bits_last(buffer_9_auto_in_bits_last),
    .auto_out_ready(buffer_9_auto_out_ready),
    .auto_out_valid(buffer_9_auto_out_valid),
    .auto_out_bits_data(buffer_9_auto_out_bits_data),
    .auto_out_bits_last(buffer_9_auto_out_bits_last)
  );
  BundleBridgeToAXI4 converter ( // @[Node.scala 65:31]
    .auto_in_aw_ready(converter_auto_in_aw_ready),
    .auto_in_aw_valid(converter_auto_in_aw_valid),
    .auto_in_aw_bits_id(converter_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(converter_auto_in_aw_bits_addr),
    .auto_in_aw_bits_size(converter_auto_in_aw_bits_size),
    .auto_in_w_ready(converter_auto_in_w_ready),
    .auto_in_w_valid(converter_auto_in_w_valid),
    .auto_in_w_bits_data(converter_auto_in_w_bits_data),
    .auto_in_w_bits_strb(converter_auto_in_w_bits_strb),
    .auto_in_w_bits_last(converter_auto_in_w_bits_last),
    .auto_in_b_ready(converter_auto_in_b_ready),
    .auto_in_b_valid(converter_auto_in_b_valid),
    .auto_in_b_bits_resp(converter_auto_in_b_bits_resp),
    .auto_in_ar_ready(converter_auto_in_ar_ready),
    .auto_in_ar_valid(converter_auto_in_ar_valid),
    .auto_in_ar_bits_id(converter_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(converter_auto_in_ar_bits_addr),
    .auto_in_ar_bits_size(converter_auto_in_ar_bits_size),
    .auto_in_r_ready(converter_auto_in_r_ready),
    .auto_in_r_valid(converter_auto_in_r_valid),
    .auto_in_r_bits_data(converter_auto_in_r_bits_data),
    .auto_in_r_bits_resp(converter_auto_in_r_bits_resp),
    .auto_in_r_bits_last(converter_auto_in_r_bits_last),
    .auto_out_aw_ready(converter_auto_out_aw_ready),
    .auto_out_aw_valid(converter_auto_out_aw_valid),
    .auto_out_aw_bits_id(converter_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(converter_auto_out_aw_bits_addr),
    .auto_out_aw_bits_size(converter_auto_out_aw_bits_size),
    .auto_out_w_ready(converter_auto_out_w_ready),
    .auto_out_w_valid(converter_auto_out_w_valid),
    .auto_out_w_bits_data(converter_auto_out_w_bits_data),
    .auto_out_w_bits_strb(converter_auto_out_w_bits_strb),
    .auto_out_w_bits_last(converter_auto_out_w_bits_last),
    .auto_out_b_ready(converter_auto_out_b_ready),
    .auto_out_b_valid(converter_auto_out_b_valid),
    .auto_out_b_bits_resp(converter_auto_out_b_bits_resp),
    .auto_out_ar_ready(converter_auto_out_ar_ready),
    .auto_out_ar_valid(converter_auto_out_ar_valid),
    .auto_out_ar_bits_id(converter_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(converter_auto_out_ar_bits_addr),
    .auto_out_ar_bits_size(converter_auto_out_ar_bits_size),
    .auto_out_r_ready(converter_auto_out_r_ready),
    .auto_out_r_valid(converter_auto_out_r_valid),
    .auto_out_r_bits_data(converter_auto_out_r_bits_data),
    .auto_out_r_bits_resp(converter_auto_out_r_bits_resp),
    .auto_out_r_bits_last(converter_auto_out_r_bits_last)
  );
  AXI4StreamToBundleBridge converter_1 ( // @[Nodes.scala 165:31]
    .auto_in_ready(converter_1_auto_in_ready),
    .auto_in_valid(converter_1_auto_in_valid),
    .auto_in_bits_data(converter_1_auto_in_bits_data),
    .auto_in_bits_last(converter_1_auto_in_bits_last),
    .auto_out_ready(converter_1_auto_out_ready),
    .auto_out_valid(converter_1_auto_out_valid),
    .auto_out_bits_data(converter_1_auto_out_bits_data),
    .auto_out_bits_last(converter_1_auto_out_bits_last)
  );
  AXI4StreamToBundleBridge converter_2 ( // @[Nodes.scala 201:31]
    .auto_in_ready(converter_2_auto_in_ready),
    .auto_in_valid(converter_2_auto_in_valid),
    .auto_in_bits_data(converter_2_auto_in_bits_data),
    .auto_in_bits_last(converter_2_auto_in_bits_last),
    .auto_out_ready(converter_2_auto_out_ready),
    .auto_out_valid(converter_2_auto_out_valid),
    .auto_out_bits_data(converter_2_auto_out_bits_data),
    .auto_out_bits_last(converter_2_auto_out_bits_last)
  );
  assign ioMem_0_aw_ready = converter_auto_in_aw_ready; // @[Nodes.scala 624:60]
  assign ioMem_0_w_ready = converter_auto_in_w_ready; // @[Nodes.scala 624:60]
  assign ioMem_0_b_valid = converter_auto_in_b_valid; // @[Nodes.scala 624:60]
  assign ioMem_0_b_bits_id = 1'h0; // @[Nodes.scala 624:60]
  assign ioMem_0_b_bits_resp = converter_auto_in_b_bits_resp; // @[Nodes.scala 624:60]
  assign ioMem_0_ar_ready = converter_auto_in_ar_ready; // @[Nodes.scala 624:60]
  assign ioMem_0_r_valid = converter_auto_in_r_valid; // @[Nodes.scala 624:60]
  assign ioMem_0_r_bits_id = 1'h0; // @[Nodes.scala 624:60]
  assign ioMem_0_r_bits_data = converter_auto_in_r_bits_data; // @[Nodes.scala 624:60]
  assign ioMem_0_r_bits_resp = converter_auto_in_r_bits_resp; // @[Nodes.scala 624:60]
  assign ioMem_0_r_bits_last = converter_auto_in_r_bits_last; // @[Nodes.scala 624:60]
  assign outStream_0_valid = converter_1_auto_out_valid; // @[Nodes.scala 649:56]
  assign outStream_0_bits_data = converter_1_auto_out_bits_data; // @[Nodes.scala 649:56]
  assign outStream_0_bits_last = converter_1_auto_out_bits_last; // @[Nodes.scala 649:56]
  assign inStream_0_ready = converter_2_auto_in_ready; // @[Nodes.scala 624:60]
  assign int_0 = uart_int_0; // @[SpectrometerTestWithoutLA.scala 206:9]
  assign uTx = uart_io_txd; // @[SpectrometerTestWithoutLA.scala 212:9]
  assign widthAdapter_clock = clock;
  assign widthAdapter_reset = reset;
  assign widthAdapter_auto_in_valid = in_queue_auto_out_out_valid; // @[LazyModule.scala 167:31]
  assign widthAdapter_auto_in_bits_data = in_queue_auto_out_out_bits_data; // @[LazyModule.scala 167:31]
  assign widthAdapter_auto_in_bits_last = in_queue_auto_out_out_bits_last; // @[LazyModule.scala 167:31]
  assign widthAdapter_auto_out_ready = in_split_auto_stream_in_ready; // @[LazyModule.scala 167:57]
  assign in_split_clock = clock;
  assign in_split_reset = reset;
  assign in_split_auto_mem_in_aw_valid = axi4buf_auto_out_aw_valid; // @[LazyModule.scala 167:31]
  assign in_split_auto_mem_in_aw_bits_id = axi4buf_auto_out_aw_bits_id; // @[LazyModule.scala 167:31]
  assign in_split_auto_mem_in_aw_bits_addr = axi4buf_auto_out_aw_bits_addr; // @[LazyModule.scala 167:31]
  assign in_split_auto_mem_in_w_valid = axi4buf_auto_out_w_valid; // @[LazyModule.scala 167:31]
  assign in_split_auto_mem_in_w_bits_data = axi4buf_auto_out_w_bits_data; // @[LazyModule.scala 167:31]
  assign in_split_auto_mem_in_w_bits_strb = axi4buf_auto_out_w_bits_strb; // @[LazyModule.scala 167:31]
  assign in_split_auto_mem_in_b_ready = axi4buf_auto_out_b_ready; // @[LazyModule.scala 167:31]
  assign in_split_auto_mem_in_ar_valid = axi4buf_auto_out_ar_valid; // @[LazyModule.scala 167:31]
  assign in_split_auto_mem_in_ar_bits_id = axi4buf_auto_out_ar_bits_id; // @[LazyModule.scala 167:31]
  assign in_split_auto_mem_in_ar_bits_addr = axi4buf_auto_out_ar_bits_addr; // @[LazyModule.scala 167:31]
  assign in_split_auto_mem_in_ar_bits_size = axi4buf_auto_out_ar_bits_size; // @[LazyModule.scala 167:31]
  assign in_split_auto_mem_in_r_ready = axi4buf_auto_out_r_ready; // @[LazyModule.scala 167:31]
  assign in_split_auto_stream_in_valid = widthAdapter_auto_out_valid; // @[LazyModule.scala 167:57]
  assign in_split_auto_stream_in_bits_data = widthAdapter_auto_out_bits_data; // @[LazyModule.scala 167:57]
  assign in_split_auto_stream_in_bits_last = widthAdapter_auto_out_bits_last; // @[LazyModule.scala 167:57]
  assign in_split_auto_stream_out_4_ready = buffer_7_auto_in_ready; // @[LazyModule.scala 167:57]
  assign in_split_auto_stream_out_3_ready = mag_mux_0_auto_stream_in_1_ready; // @[LazyModule.scala 167:57]
  assign in_split_auto_stream_out_2_ready = fft_mux_0_auto_stream_in_1_ready; // @[LazyModule.scala 167:57]
  assign in_split_auto_stream_out_1_ready = nco_mux_0_auto_stream_in_1_ready; // @[LazyModule.scala 167:57]
  assign in_split_auto_stream_out_0_ready = plfg_mux_0_auto_stream_in_1_ready; // @[LazyModule.scala 167:57]
  assign in_queue_clock = clock;
  assign in_queue_reset = reset;
  assign in_queue_auto_out_out_ready = widthAdapter_auto_in_ready; // @[LazyModule.scala 167:31]
  assign in_queue_auto_in_in_valid = converter_2_auto_out_valid; // @[LazyModule.scala 167:31]
  assign in_queue_auto_in_in_bits_data = converter_2_auto_out_bits_data; // @[LazyModule.scala 167:31]
  assign in_queue_auto_in_in_bits_last = converter_2_auto_out_bits_last; // @[LazyModule.scala 167:31]
  assign plfg_clock = clock;
  assign plfg_reset = reset;
  assign plfg_auto_mem_in_aw_valid = axi4buf_1_auto_out_aw_valid; // @[LazyModule.scala 167:31]
  assign plfg_auto_mem_in_aw_bits_id = axi4buf_1_auto_out_aw_bits_id; // @[LazyModule.scala 167:31]
  assign plfg_auto_mem_in_aw_bits_addr = axi4buf_1_auto_out_aw_bits_addr; // @[LazyModule.scala 167:31]
  assign plfg_auto_mem_in_w_valid = axi4buf_1_auto_out_w_valid; // @[LazyModule.scala 167:31]
  assign plfg_auto_mem_in_w_bits_data = axi4buf_1_auto_out_w_bits_data; // @[LazyModule.scala 167:31]
  assign plfg_auto_mem_in_w_bits_strb = axi4buf_1_auto_out_w_bits_strb; // @[LazyModule.scala 167:31]
  assign plfg_auto_mem_in_w_bits_last = axi4buf_1_auto_out_w_bits_last; // @[LazyModule.scala 167:31]
  assign plfg_auto_mem_in_b_ready = axi4buf_1_auto_out_b_ready; // @[LazyModule.scala 167:31]
  assign plfg_auto_mem_in_ar_valid = axi4buf_1_auto_out_ar_valid; // @[LazyModule.scala 167:31]
  assign plfg_auto_mem_in_ar_bits_id = axi4buf_1_auto_out_ar_bits_id; // @[LazyModule.scala 167:31]
  assign plfg_auto_mem_in_ar_bits_addr = axi4buf_1_auto_out_ar_bits_addr; // @[LazyModule.scala 167:31]
  assign plfg_auto_mem_in_ar_bits_size = axi4buf_1_auto_out_ar_bits_size; // @[LazyModule.scala 167:31]
  assign plfg_auto_mem_in_r_ready = axi4buf_1_auto_out_r_ready; // @[LazyModule.scala 167:31]
  assign plfg_auto_stream_out_ready = plfg_split_auto_stream_in_ready; // @[LazyModule.scala 167:57]
  assign plfg_split_clock = clock;
  assign plfg_split_reset = reset;
  assign plfg_split_auto_mem_in_aw_valid = axi4buf_2_auto_out_aw_valid; // @[LazyModule.scala 167:31]
  assign plfg_split_auto_mem_in_aw_bits_id = axi4buf_2_auto_out_aw_bits_id; // @[LazyModule.scala 167:31]
  assign plfg_split_auto_mem_in_aw_bits_addr = axi4buf_2_auto_out_aw_bits_addr; // @[LazyModule.scala 167:31]
  assign plfg_split_auto_mem_in_w_valid = axi4buf_2_auto_out_w_valid; // @[LazyModule.scala 167:31]
  assign plfg_split_auto_mem_in_w_bits_data = axi4buf_2_auto_out_w_bits_data; // @[LazyModule.scala 167:31]
  assign plfg_split_auto_mem_in_w_bits_strb = axi4buf_2_auto_out_w_bits_strb; // @[LazyModule.scala 167:31]
  assign plfg_split_auto_mem_in_b_ready = axi4buf_2_auto_out_b_ready; // @[LazyModule.scala 167:31]
  assign plfg_split_auto_mem_in_ar_valid = axi4buf_2_auto_out_ar_valid; // @[LazyModule.scala 167:31]
  assign plfg_split_auto_mem_in_ar_bits_id = axi4buf_2_auto_out_ar_bits_id; // @[LazyModule.scala 167:31]
  assign plfg_split_auto_mem_in_ar_bits_addr = axi4buf_2_auto_out_ar_bits_addr; // @[LazyModule.scala 167:31]
  assign plfg_split_auto_mem_in_ar_bits_size = axi4buf_2_auto_out_ar_bits_size; // @[LazyModule.scala 167:31]
  assign plfg_split_auto_mem_in_r_ready = axi4buf_2_auto_out_r_ready; // @[LazyModule.scala 167:31]
  assign plfg_split_auto_stream_in_valid = plfg_auto_stream_out_valid; // @[LazyModule.scala 167:57]
  assign plfg_split_auto_stream_in_bits_data = plfg_auto_stream_out_bits_data; // @[LazyModule.scala 167:57]
  assign plfg_split_auto_stream_in_bits_last = plfg_auto_stream_out_bits_last; // @[LazyModule.scala 167:57]
  assign plfg_split_auto_stream_out_1_ready = plfg_mux_0_auto_stream_in_0_ready; // @[LazyModule.scala 167:57]
  assign plfg_split_auto_stream_out_0_ready = plfg_mux_1_auto_stream_in_ready; // @[LazyModule.scala 167:57]
  assign plfg_mux_0_clock = clock;
  assign plfg_mux_0_reset = reset;
  assign plfg_mux_0_auto_register_in_aw_valid = axi4buf_3_auto_out_aw_valid; // @[LazyModule.scala 167:31]
  assign plfg_mux_0_auto_register_in_aw_bits_id = axi4buf_3_auto_out_aw_bits_id; // @[LazyModule.scala 167:31]
  assign plfg_mux_0_auto_register_in_aw_bits_addr = axi4buf_3_auto_out_aw_bits_addr; // @[LazyModule.scala 167:31]
  assign plfg_mux_0_auto_register_in_w_valid = axi4buf_3_auto_out_w_valid; // @[LazyModule.scala 167:31]
  assign plfg_mux_0_auto_register_in_w_bits_data = axi4buf_3_auto_out_w_bits_data; // @[LazyModule.scala 167:31]
  assign plfg_mux_0_auto_register_in_w_bits_strb = axi4buf_3_auto_out_w_bits_strb; // @[LazyModule.scala 167:31]
  assign plfg_mux_0_auto_register_in_b_ready = axi4buf_3_auto_out_b_ready; // @[LazyModule.scala 167:31]
  assign plfg_mux_0_auto_register_in_ar_valid = axi4buf_3_auto_out_ar_valid; // @[LazyModule.scala 167:31]
  assign plfg_mux_0_auto_register_in_ar_bits_id = axi4buf_3_auto_out_ar_bits_id; // @[LazyModule.scala 167:31]
  assign plfg_mux_0_auto_register_in_ar_bits_addr = axi4buf_3_auto_out_ar_bits_addr; // @[LazyModule.scala 167:31]
  assign plfg_mux_0_auto_register_in_ar_bits_size = axi4buf_3_auto_out_ar_bits_size; // @[LazyModule.scala 167:31]
  assign plfg_mux_0_auto_register_in_r_ready = axi4buf_3_auto_out_r_ready; // @[LazyModule.scala 167:31]
  assign plfg_mux_0_auto_stream_in_2_valid = uRx_split_auto_stream_out_0_valid; // @[LazyModule.scala 167:31]
  assign plfg_mux_0_auto_stream_in_2_bits_data = uRx_split_auto_stream_out_0_bits_data; // @[LazyModule.scala 167:31]
  assign plfg_mux_0_auto_stream_in_2_bits_last = uRx_split_auto_stream_out_0_bits_last; // @[LazyModule.scala 167:31]
  assign plfg_mux_0_auto_stream_in_1_valid = in_split_auto_stream_out_0_valid; // @[LazyModule.scala 167:57]
  assign plfg_mux_0_auto_stream_in_1_bits_data = in_split_auto_stream_out_0_bits_data; // @[LazyModule.scala 167:57]
  assign plfg_mux_0_auto_stream_in_1_bits_last = in_split_auto_stream_out_0_bits_last; // @[LazyModule.scala 167:57]
  assign plfg_mux_0_auto_stream_in_0_valid = plfg_split_auto_stream_out_1_valid; // @[LazyModule.scala 167:57]
  assign plfg_mux_0_auto_stream_in_0_bits_data = plfg_split_auto_stream_out_1_bits_data; // @[LazyModule.scala 167:57]
  assign plfg_mux_0_auto_stream_in_0_bits_last = plfg_split_auto_stream_out_1_bits_last; // @[LazyModule.scala 167:57]
  assign plfg_mux_0_auto_stream_out_0_ready = nco_auto_freq_in_ready; // @[LazyModule.scala 167:57]
  assign plfg_mux_1_clock = clock;
  assign plfg_mux_1_reset = reset;
  assign plfg_mux_1_auto_register_in_aw_valid = axi4buf_4_auto_out_aw_valid; // @[LazyModule.scala 167:31]
  assign plfg_mux_1_auto_register_in_aw_bits_id = axi4buf_4_auto_out_aw_bits_id; // @[LazyModule.scala 167:31]
  assign plfg_mux_1_auto_register_in_aw_bits_addr = axi4buf_4_auto_out_aw_bits_addr; // @[LazyModule.scala 167:31]
  assign plfg_mux_1_auto_register_in_w_valid = axi4buf_4_auto_out_w_valid; // @[LazyModule.scala 167:31]
  assign plfg_mux_1_auto_register_in_w_bits_data = axi4buf_4_auto_out_w_bits_data; // @[LazyModule.scala 167:31]
  assign plfg_mux_1_auto_register_in_w_bits_strb = axi4buf_4_auto_out_w_bits_strb; // @[LazyModule.scala 167:31]
  assign plfg_mux_1_auto_register_in_b_ready = axi4buf_4_auto_out_b_ready; // @[LazyModule.scala 167:31]
  assign plfg_mux_1_auto_register_in_ar_valid = axi4buf_4_auto_out_ar_valid; // @[LazyModule.scala 167:31]
  assign plfg_mux_1_auto_register_in_ar_bits_id = axi4buf_4_auto_out_ar_bits_id; // @[LazyModule.scala 167:31]
  assign plfg_mux_1_auto_register_in_ar_bits_addr = axi4buf_4_auto_out_ar_bits_addr; // @[LazyModule.scala 167:31]
  assign plfg_mux_1_auto_register_in_ar_bits_size = axi4buf_4_auto_out_ar_bits_size; // @[LazyModule.scala 167:31]
  assign plfg_mux_1_auto_register_in_r_ready = axi4buf_4_auto_out_r_ready; // @[LazyModule.scala 167:31]
  assign plfg_mux_1_auto_stream_in_valid = plfg_split_auto_stream_out_0_valid; // @[LazyModule.scala 167:57]
  assign plfg_mux_1_auto_stream_in_bits_data = plfg_split_auto_stream_out_0_bits_data; // @[LazyModule.scala 167:57]
  assign plfg_mux_1_auto_stream_in_bits_last = plfg_split_auto_stream_out_0_bits_last; // @[LazyModule.scala 167:57]
  assign plfg_mux_1_auto_stream_out_1_ready = buffer_6_auto_in_ready; // @[LazyModule.scala 167:57]
  assign nco_clock = clock;
  assign nco_reset = reset;
  assign nco_auto_stream_out_ready = nco_split_auto_stream_in_ready; // @[LazyModule.scala 167:57]
  assign nco_auto_freq_in_valid = plfg_mux_0_auto_stream_out_0_valid; // @[LazyModule.scala 167:57]
  assign nco_auto_freq_in_bits_data = plfg_mux_0_auto_stream_out_0_bits_data; // @[LazyModule.scala 167:57]
  assign nco_auto_freq_in_bits_last = plfg_mux_0_auto_stream_out_0_bits_last; // @[LazyModule.scala 167:57]
  assign nco_split_clock = clock;
  assign nco_split_reset = reset;
  assign nco_split_auto_mem_in_aw_valid = axi4buf_6_auto_out_aw_valid; // @[LazyModule.scala 167:31]
  assign nco_split_auto_mem_in_aw_bits_id = axi4buf_6_auto_out_aw_bits_id; // @[LazyModule.scala 167:31]
  assign nco_split_auto_mem_in_aw_bits_addr = axi4buf_6_auto_out_aw_bits_addr; // @[LazyModule.scala 167:31]
  assign nco_split_auto_mem_in_w_valid = axi4buf_6_auto_out_w_valid; // @[LazyModule.scala 167:31]
  assign nco_split_auto_mem_in_w_bits_data = axi4buf_6_auto_out_w_bits_data; // @[LazyModule.scala 167:31]
  assign nco_split_auto_mem_in_w_bits_strb = axi4buf_6_auto_out_w_bits_strb; // @[LazyModule.scala 167:31]
  assign nco_split_auto_mem_in_b_ready = axi4buf_6_auto_out_b_ready; // @[LazyModule.scala 167:31]
  assign nco_split_auto_mem_in_ar_valid = axi4buf_6_auto_out_ar_valid; // @[LazyModule.scala 167:31]
  assign nco_split_auto_mem_in_ar_bits_id = axi4buf_6_auto_out_ar_bits_id; // @[LazyModule.scala 167:31]
  assign nco_split_auto_mem_in_ar_bits_addr = axi4buf_6_auto_out_ar_bits_addr; // @[LazyModule.scala 167:31]
  assign nco_split_auto_mem_in_ar_bits_size = axi4buf_6_auto_out_ar_bits_size; // @[LazyModule.scala 167:31]
  assign nco_split_auto_mem_in_r_ready = axi4buf_6_auto_out_r_ready; // @[LazyModule.scala 167:31]
  assign nco_split_auto_stream_in_valid = nco_auto_stream_out_valid; // @[LazyModule.scala 167:57]
  assign nco_split_auto_stream_in_bits_data = nco_auto_stream_out_bits_data; // @[LazyModule.scala 167:57]
  assign nco_split_auto_stream_in_bits_last = nco_auto_stream_out_bits_last; // @[LazyModule.scala 167:57]
  assign nco_split_auto_stream_out_1_ready = nco_mux_0_auto_stream_in_0_ready; // @[LazyModule.scala 167:57]
  assign nco_split_auto_stream_out_0_ready = nco_mux_1_auto_stream_in_ready; // @[LazyModule.scala 167:57]
  assign nco_mux_0_clock = clock;
  assign nco_mux_0_reset = reset;
  assign nco_mux_0_auto_register_in_aw_valid = axi4buf_7_auto_out_aw_valid; // @[LazyModule.scala 167:31]
  assign nco_mux_0_auto_register_in_aw_bits_id = axi4buf_7_auto_out_aw_bits_id; // @[LazyModule.scala 167:31]
  assign nco_mux_0_auto_register_in_aw_bits_addr = axi4buf_7_auto_out_aw_bits_addr; // @[LazyModule.scala 167:31]
  assign nco_mux_0_auto_register_in_w_valid = axi4buf_7_auto_out_w_valid; // @[LazyModule.scala 167:31]
  assign nco_mux_0_auto_register_in_w_bits_data = axi4buf_7_auto_out_w_bits_data; // @[LazyModule.scala 167:31]
  assign nco_mux_0_auto_register_in_w_bits_strb = axi4buf_7_auto_out_w_bits_strb; // @[LazyModule.scala 167:31]
  assign nco_mux_0_auto_register_in_b_ready = axi4buf_7_auto_out_b_ready; // @[LazyModule.scala 167:31]
  assign nco_mux_0_auto_register_in_ar_valid = axi4buf_7_auto_out_ar_valid; // @[LazyModule.scala 167:31]
  assign nco_mux_0_auto_register_in_ar_bits_id = axi4buf_7_auto_out_ar_bits_id; // @[LazyModule.scala 167:31]
  assign nco_mux_0_auto_register_in_ar_bits_addr = axi4buf_7_auto_out_ar_bits_addr; // @[LazyModule.scala 167:31]
  assign nco_mux_0_auto_register_in_ar_bits_size = axi4buf_7_auto_out_ar_bits_size; // @[LazyModule.scala 167:31]
  assign nco_mux_0_auto_register_in_r_ready = axi4buf_7_auto_out_r_ready; // @[LazyModule.scala 167:31]
  assign nco_mux_0_auto_stream_in_2_valid = uRx_split_auto_stream_out_1_valid; // @[LazyModule.scala 167:31]
  assign nco_mux_0_auto_stream_in_2_bits_data = uRx_split_auto_stream_out_1_bits_data; // @[LazyModule.scala 167:31]
  assign nco_mux_0_auto_stream_in_2_bits_last = uRx_split_auto_stream_out_1_bits_last; // @[LazyModule.scala 167:31]
  assign nco_mux_0_auto_stream_in_1_valid = in_split_auto_stream_out_1_valid; // @[LazyModule.scala 167:57]
  assign nco_mux_0_auto_stream_in_1_bits_data = in_split_auto_stream_out_1_bits_data; // @[LazyModule.scala 167:57]
  assign nco_mux_0_auto_stream_in_1_bits_last = in_split_auto_stream_out_1_bits_last; // @[LazyModule.scala 167:57]
  assign nco_mux_0_auto_stream_in_0_valid = nco_split_auto_stream_out_1_valid; // @[LazyModule.scala 167:57]
  assign nco_mux_0_auto_stream_in_0_bits_data = nco_split_auto_stream_out_1_bits_data; // @[LazyModule.scala 167:57]
  assign nco_mux_0_auto_stream_in_0_bits_last = nco_split_auto_stream_out_1_bits_last; // @[LazyModule.scala 167:57]
  assign nco_mux_0_auto_stream_out_0_ready = buffer_auto_in_ready; // @[LazyModule.scala 167:57]
  assign nco_mux_1_clock = clock;
  assign nco_mux_1_reset = reset;
  assign nco_mux_1_auto_register_in_aw_valid = axi4buf_8_auto_out_aw_valid; // @[LazyModule.scala 167:31]
  assign nco_mux_1_auto_register_in_aw_bits_id = axi4buf_8_auto_out_aw_bits_id; // @[LazyModule.scala 167:31]
  assign nco_mux_1_auto_register_in_aw_bits_addr = axi4buf_8_auto_out_aw_bits_addr; // @[LazyModule.scala 167:31]
  assign nco_mux_1_auto_register_in_w_valid = axi4buf_8_auto_out_w_valid; // @[LazyModule.scala 167:31]
  assign nco_mux_1_auto_register_in_w_bits_data = axi4buf_8_auto_out_w_bits_data; // @[LazyModule.scala 167:31]
  assign nco_mux_1_auto_register_in_w_bits_strb = axi4buf_8_auto_out_w_bits_strb; // @[LazyModule.scala 167:31]
  assign nco_mux_1_auto_register_in_b_ready = axi4buf_8_auto_out_b_ready; // @[LazyModule.scala 167:31]
  assign nco_mux_1_auto_register_in_ar_valid = axi4buf_8_auto_out_ar_valid; // @[LazyModule.scala 167:31]
  assign nco_mux_1_auto_register_in_ar_bits_id = axi4buf_8_auto_out_ar_bits_id; // @[LazyModule.scala 167:31]
  assign nco_mux_1_auto_register_in_ar_bits_addr = axi4buf_8_auto_out_ar_bits_addr; // @[LazyModule.scala 167:31]
  assign nco_mux_1_auto_register_in_ar_bits_size = axi4buf_8_auto_out_ar_bits_size; // @[LazyModule.scala 167:31]
  assign nco_mux_1_auto_register_in_r_ready = axi4buf_8_auto_out_r_ready; // @[LazyModule.scala 167:31]
  assign nco_mux_1_auto_stream_in_valid = nco_split_auto_stream_out_0_valid; // @[LazyModule.scala 167:57]
  assign nco_mux_1_auto_stream_in_bits_data = nco_split_auto_stream_out_0_bits_data; // @[LazyModule.scala 167:57]
  assign nco_mux_1_auto_stream_in_bits_last = nco_split_auto_stream_out_0_bits_last; // @[LazyModule.scala 167:57]
  assign nco_mux_1_auto_stream_out_1_ready = buffer_5_auto_in_ready; // @[LazyModule.scala 167:57]
  assign fft_clock = clock;
  assign fft_reset = reset;
  assign fft_auto_mem_in_aw_valid = axi4buf_9_auto_out_aw_valid; // @[LazyModule.scala 167:31]
  assign fft_auto_mem_in_aw_bits_id = axi4buf_9_auto_out_aw_bits_id; // @[LazyModule.scala 167:31]
  assign fft_auto_mem_in_aw_bits_addr = axi4buf_9_auto_out_aw_bits_addr; // @[LazyModule.scala 167:31]
  assign fft_auto_mem_in_w_valid = axi4buf_9_auto_out_w_valid; // @[LazyModule.scala 167:31]
  assign fft_auto_mem_in_w_bits_data = axi4buf_9_auto_out_w_bits_data; // @[LazyModule.scala 167:31]
  assign fft_auto_mem_in_w_bits_strb = axi4buf_9_auto_out_w_bits_strb; // @[LazyModule.scala 167:31]
  assign fft_auto_mem_in_b_ready = axi4buf_9_auto_out_b_ready; // @[LazyModule.scala 167:31]
  assign fft_auto_mem_in_ar_valid = axi4buf_9_auto_out_ar_valid; // @[LazyModule.scala 167:31]
  assign fft_auto_mem_in_ar_bits_id = axi4buf_9_auto_out_ar_bits_id; // @[LazyModule.scala 167:31]
  assign fft_auto_mem_in_ar_bits_addr = axi4buf_9_auto_out_ar_bits_addr; // @[LazyModule.scala 167:31]
  assign fft_auto_mem_in_ar_bits_size = axi4buf_9_auto_out_ar_bits_size; // @[LazyModule.scala 167:31]
  assign fft_auto_mem_in_r_ready = axi4buf_9_auto_out_r_ready; // @[LazyModule.scala 167:31]
  assign fft_auto_stream_in_valid = buffer_auto_out_valid; // @[LazyModule.scala 167:31]
  assign fft_auto_stream_in_bits_data = buffer_auto_out_bits_data; // @[LazyModule.scala 167:31]
  assign fft_auto_stream_in_bits_last = buffer_auto_out_bits_last; // @[LazyModule.scala 167:31]
  assign fft_auto_stream_out_ready = fft_split_auto_stream_in_ready; // @[LazyModule.scala 167:57]
  assign fft_split_clock = clock;
  assign fft_split_reset = reset;
  assign fft_split_auto_mem_in_aw_valid = axi4buf_10_auto_out_aw_valid; // @[LazyModule.scala 167:31]
  assign fft_split_auto_mem_in_aw_bits_id = axi4buf_10_auto_out_aw_bits_id; // @[LazyModule.scala 167:31]
  assign fft_split_auto_mem_in_aw_bits_addr = axi4buf_10_auto_out_aw_bits_addr; // @[LazyModule.scala 167:31]
  assign fft_split_auto_mem_in_w_valid = axi4buf_10_auto_out_w_valid; // @[LazyModule.scala 167:31]
  assign fft_split_auto_mem_in_w_bits_data = axi4buf_10_auto_out_w_bits_data; // @[LazyModule.scala 167:31]
  assign fft_split_auto_mem_in_w_bits_strb = axi4buf_10_auto_out_w_bits_strb; // @[LazyModule.scala 167:31]
  assign fft_split_auto_mem_in_b_ready = axi4buf_10_auto_out_b_ready; // @[LazyModule.scala 167:31]
  assign fft_split_auto_mem_in_ar_valid = axi4buf_10_auto_out_ar_valid; // @[LazyModule.scala 167:31]
  assign fft_split_auto_mem_in_ar_bits_id = axi4buf_10_auto_out_ar_bits_id; // @[LazyModule.scala 167:31]
  assign fft_split_auto_mem_in_ar_bits_addr = axi4buf_10_auto_out_ar_bits_addr; // @[LazyModule.scala 167:31]
  assign fft_split_auto_mem_in_ar_bits_size = axi4buf_10_auto_out_ar_bits_size; // @[LazyModule.scala 167:31]
  assign fft_split_auto_mem_in_r_ready = axi4buf_10_auto_out_r_ready; // @[LazyModule.scala 167:31]
  assign fft_split_auto_stream_in_valid = fft_auto_stream_out_valid; // @[LazyModule.scala 167:57]
  assign fft_split_auto_stream_in_bits_data = fft_auto_stream_out_bits_data; // @[LazyModule.scala 167:57]
  assign fft_split_auto_stream_in_bits_last = fft_auto_stream_out_bits_last; // @[LazyModule.scala 167:57]
  assign fft_split_auto_stream_out_1_ready = fft_mux_0_auto_stream_in_0_ready; // @[LazyModule.scala 167:57]
  assign fft_split_auto_stream_out_0_ready = fft_mux_1_auto_stream_in_ready; // @[LazyModule.scala 167:57]
  assign fft_mux_0_clock = clock;
  assign fft_mux_0_reset = reset;
  assign fft_mux_0_auto_register_in_aw_valid = axi4buf_11_auto_out_aw_valid; // @[LazyModule.scala 167:31]
  assign fft_mux_0_auto_register_in_aw_bits_id = axi4buf_11_auto_out_aw_bits_id; // @[LazyModule.scala 167:31]
  assign fft_mux_0_auto_register_in_aw_bits_addr = axi4buf_11_auto_out_aw_bits_addr; // @[LazyModule.scala 167:31]
  assign fft_mux_0_auto_register_in_w_valid = axi4buf_11_auto_out_w_valid; // @[LazyModule.scala 167:31]
  assign fft_mux_0_auto_register_in_w_bits_data = axi4buf_11_auto_out_w_bits_data; // @[LazyModule.scala 167:31]
  assign fft_mux_0_auto_register_in_w_bits_strb = axi4buf_11_auto_out_w_bits_strb; // @[LazyModule.scala 167:31]
  assign fft_mux_0_auto_register_in_b_ready = axi4buf_11_auto_out_b_ready; // @[LazyModule.scala 167:31]
  assign fft_mux_0_auto_register_in_ar_valid = axi4buf_11_auto_out_ar_valid; // @[LazyModule.scala 167:31]
  assign fft_mux_0_auto_register_in_ar_bits_id = axi4buf_11_auto_out_ar_bits_id; // @[LazyModule.scala 167:31]
  assign fft_mux_0_auto_register_in_ar_bits_addr = axi4buf_11_auto_out_ar_bits_addr; // @[LazyModule.scala 167:31]
  assign fft_mux_0_auto_register_in_ar_bits_size = axi4buf_11_auto_out_ar_bits_size; // @[LazyModule.scala 167:31]
  assign fft_mux_0_auto_register_in_r_ready = axi4buf_11_auto_out_r_ready; // @[LazyModule.scala 167:31]
  assign fft_mux_0_auto_stream_in_2_valid = uRx_split_auto_stream_out_2_valid; // @[LazyModule.scala 167:31]
  assign fft_mux_0_auto_stream_in_2_bits_data = uRx_split_auto_stream_out_2_bits_data; // @[LazyModule.scala 167:31]
  assign fft_mux_0_auto_stream_in_2_bits_last = uRx_split_auto_stream_out_2_bits_last; // @[LazyModule.scala 167:31]
  assign fft_mux_0_auto_stream_in_1_valid = in_split_auto_stream_out_2_valid; // @[LazyModule.scala 167:57]
  assign fft_mux_0_auto_stream_in_1_bits_data = in_split_auto_stream_out_2_bits_data; // @[LazyModule.scala 167:57]
  assign fft_mux_0_auto_stream_in_1_bits_last = in_split_auto_stream_out_2_bits_last; // @[LazyModule.scala 167:57]
  assign fft_mux_0_auto_stream_in_0_valid = fft_split_auto_stream_out_1_valid; // @[LazyModule.scala 167:57]
  assign fft_mux_0_auto_stream_in_0_bits_data = fft_split_auto_stream_out_1_bits_data; // @[LazyModule.scala 167:57]
  assign fft_mux_0_auto_stream_in_0_bits_last = fft_split_auto_stream_out_1_bits_last; // @[LazyModule.scala 167:57]
  assign fft_mux_0_auto_stream_out_0_ready = buffer_1_auto_in_ready; // @[LazyModule.scala 167:57]
  assign fft_mux_1_clock = clock;
  assign fft_mux_1_reset = reset;
  assign fft_mux_1_auto_register_in_aw_valid = axi4buf_12_auto_out_aw_valid; // @[LazyModule.scala 167:31]
  assign fft_mux_1_auto_register_in_aw_bits_id = axi4buf_12_auto_out_aw_bits_id; // @[LazyModule.scala 167:31]
  assign fft_mux_1_auto_register_in_aw_bits_addr = axi4buf_12_auto_out_aw_bits_addr; // @[LazyModule.scala 167:31]
  assign fft_mux_1_auto_register_in_w_valid = axi4buf_12_auto_out_w_valid; // @[LazyModule.scala 167:31]
  assign fft_mux_1_auto_register_in_w_bits_data = axi4buf_12_auto_out_w_bits_data; // @[LazyModule.scala 167:31]
  assign fft_mux_1_auto_register_in_w_bits_strb = axi4buf_12_auto_out_w_bits_strb; // @[LazyModule.scala 167:31]
  assign fft_mux_1_auto_register_in_b_ready = axi4buf_12_auto_out_b_ready; // @[LazyModule.scala 167:31]
  assign fft_mux_1_auto_register_in_ar_valid = axi4buf_12_auto_out_ar_valid; // @[LazyModule.scala 167:31]
  assign fft_mux_1_auto_register_in_ar_bits_id = axi4buf_12_auto_out_ar_bits_id; // @[LazyModule.scala 167:31]
  assign fft_mux_1_auto_register_in_ar_bits_addr = axi4buf_12_auto_out_ar_bits_addr; // @[LazyModule.scala 167:31]
  assign fft_mux_1_auto_register_in_ar_bits_size = axi4buf_12_auto_out_ar_bits_size; // @[LazyModule.scala 167:31]
  assign fft_mux_1_auto_register_in_r_ready = axi4buf_12_auto_out_r_ready; // @[LazyModule.scala 167:31]
  assign fft_mux_1_auto_stream_in_valid = fft_split_auto_stream_out_0_valid; // @[LazyModule.scala 167:57]
  assign fft_mux_1_auto_stream_in_bits_data = fft_split_auto_stream_out_0_bits_data; // @[LazyModule.scala 167:57]
  assign fft_mux_1_auto_stream_in_bits_last = fft_split_auto_stream_out_0_bits_last; // @[LazyModule.scala 167:57]
  assign fft_mux_1_auto_stream_out_1_ready = buffer_4_auto_in_ready; // @[LazyModule.scala 167:57]
  assign mag_clock = clock;
  assign mag_reset = reset;
  assign mag_auto_mem_in_aw_valid = axi4buf_13_auto_out_aw_valid; // @[LazyModule.scala 167:31]
  assign mag_auto_mem_in_aw_bits_id = axi4buf_13_auto_out_aw_bits_id; // @[LazyModule.scala 167:31]
  assign mag_auto_mem_in_aw_bits_addr = axi4buf_13_auto_out_aw_bits_addr; // @[LazyModule.scala 167:31]
  assign mag_auto_mem_in_w_valid = axi4buf_13_auto_out_w_valid; // @[LazyModule.scala 167:31]
  assign mag_auto_mem_in_w_bits_data = axi4buf_13_auto_out_w_bits_data; // @[LazyModule.scala 167:31]
  assign mag_auto_mem_in_w_bits_strb = axi4buf_13_auto_out_w_bits_strb; // @[LazyModule.scala 167:31]
  assign mag_auto_mem_in_b_ready = axi4buf_13_auto_out_b_ready; // @[LazyModule.scala 167:31]
  assign mag_auto_mem_in_ar_valid = axi4buf_13_auto_out_ar_valid; // @[LazyModule.scala 167:31]
  assign mag_auto_mem_in_ar_bits_id = axi4buf_13_auto_out_ar_bits_id; // @[LazyModule.scala 167:31]
  assign mag_auto_mem_in_ar_bits_addr = axi4buf_13_auto_out_ar_bits_addr; // @[LazyModule.scala 167:31]
  assign mag_auto_mem_in_ar_bits_size = axi4buf_13_auto_out_ar_bits_size; // @[LazyModule.scala 167:31]
  assign mag_auto_mem_in_r_ready = axi4buf_13_auto_out_r_ready; // @[LazyModule.scala 167:31]
  assign mag_auto_stream_in_valid = buffer_1_auto_out_valid; // @[LazyModule.scala 167:31]
  assign mag_auto_stream_in_bits_data = buffer_1_auto_out_bits_data; // @[LazyModule.scala 167:31]
  assign mag_auto_stream_in_bits_last = buffer_1_auto_out_bits_last; // @[LazyModule.scala 167:31]
  assign mag_auto_stream_out_ready = mag_split_auto_stream_in_ready; // @[LazyModule.scala 167:57]
  assign mag_split_clock = clock;
  assign mag_split_reset = reset;
  assign mag_split_auto_mem_in_aw_valid = axi4buf_14_auto_out_aw_valid; // @[LazyModule.scala 167:31]
  assign mag_split_auto_mem_in_aw_bits_id = axi4buf_14_auto_out_aw_bits_id; // @[LazyModule.scala 167:31]
  assign mag_split_auto_mem_in_aw_bits_addr = axi4buf_14_auto_out_aw_bits_addr; // @[LazyModule.scala 167:31]
  assign mag_split_auto_mem_in_w_valid = axi4buf_14_auto_out_w_valid; // @[LazyModule.scala 167:31]
  assign mag_split_auto_mem_in_w_bits_data = axi4buf_14_auto_out_w_bits_data; // @[LazyModule.scala 167:31]
  assign mag_split_auto_mem_in_w_bits_strb = axi4buf_14_auto_out_w_bits_strb; // @[LazyModule.scala 167:31]
  assign mag_split_auto_mem_in_b_ready = axi4buf_14_auto_out_b_ready; // @[LazyModule.scala 167:31]
  assign mag_split_auto_mem_in_ar_valid = axi4buf_14_auto_out_ar_valid; // @[LazyModule.scala 167:31]
  assign mag_split_auto_mem_in_ar_bits_id = axi4buf_14_auto_out_ar_bits_id; // @[LazyModule.scala 167:31]
  assign mag_split_auto_mem_in_ar_bits_addr = axi4buf_14_auto_out_ar_bits_addr; // @[LazyModule.scala 167:31]
  assign mag_split_auto_mem_in_ar_bits_size = axi4buf_14_auto_out_ar_bits_size; // @[LazyModule.scala 167:31]
  assign mag_split_auto_mem_in_r_ready = axi4buf_14_auto_out_r_ready; // @[LazyModule.scala 167:31]
  assign mag_split_auto_stream_in_valid = mag_auto_stream_out_valid; // @[LazyModule.scala 167:57]
  assign mag_split_auto_stream_in_bits_data = mag_auto_stream_out_bits_data; // @[LazyModule.scala 167:57]
  assign mag_split_auto_stream_in_bits_last = mag_auto_stream_out_bits_last; // @[LazyModule.scala 167:57]
  assign mag_split_auto_stream_out_1_ready = mag_mux_0_auto_stream_in_0_ready; // @[LazyModule.scala 167:57]
  assign mag_split_auto_stream_out_0_ready = mag_mux_1_auto_stream_in_ready; // @[LazyModule.scala 167:57]
  assign mag_mux_0_clock = clock;
  assign mag_mux_0_reset = reset;
  assign mag_mux_0_auto_register_in_aw_valid = axi4buf_15_auto_out_aw_valid; // @[LazyModule.scala 167:31]
  assign mag_mux_0_auto_register_in_aw_bits_id = axi4buf_15_auto_out_aw_bits_id; // @[LazyModule.scala 167:31]
  assign mag_mux_0_auto_register_in_aw_bits_addr = axi4buf_15_auto_out_aw_bits_addr; // @[LazyModule.scala 167:31]
  assign mag_mux_0_auto_register_in_w_valid = axi4buf_15_auto_out_w_valid; // @[LazyModule.scala 167:31]
  assign mag_mux_0_auto_register_in_w_bits_data = axi4buf_15_auto_out_w_bits_data; // @[LazyModule.scala 167:31]
  assign mag_mux_0_auto_register_in_w_bits_strb = axi4buf_15_auto_out_w_bits_strb; // @[LazyModule.scala 167:31]
  assign mag_mux_0_auto_register_in_b_ready = axi4buf_15_auto_out_b_ready; // @[LazyModule.scala 167:31]
  assign mag_mux_0_auto_register_in_ar_valid = axi4buf_15_auto_out_ar_valid; // @[LazyModule.scala 167:31]
  assign mag_mux_0_auto_register_in_ar_bits_id = axi4buf_15_auto_out_ar_bits_id; // @[LazyModule.scala 167:31]
  assign mag_mux_0_auto_register_in_ar_bits_addr = axi4buf_15_auto_out_ar_bits_addr; // @[LazyModule.scala 167:31]
  assign mag_mux_0_auto_register_in_ar_bits_size = axi4buf_15_auto_out_ar_bits_size; // @[LazyModule.scala 167:31]
  assign mag_mux_0_auto_register_in_r_ready = axi4buf_15_auto_out_r_ready; // @[LazyModule.scala 167:31]
  assign mag_mux_0_auto_stream_in_2_valid = uRx_split_auto_stream_out_3_valid; // @[LazyModule.scala 167:31]
  assign mag_mux_0_auto_stream_in_2_bits_data = uRx_split_auto_stream_out_3_bits_data; // @[LazyModule.scala 167:31]
  assign mag_mux_0_auto_stream_in_2_bits_last = uRx_split_auto_stream_out_3_bits_last; // @[LazyModule.scala 167:31]
  assign mag_mux_0_auto_stream_in_1_valid = in_split_auto_stream_out_3_valid; // @[LazyModule.scala 167:57]
  assign mag_mux_0_auto_stream_in_1_bits_data = in_split_auto_stream_out_3_bits_data; // @[LazyModule.scala 167:57]
  assign mag_mux_0_auto_stream_in_1_bits_last = in_split_auto_stream_out_3_bits_last; // @[LazyModule.scala 167:57]
  assign mag_mux_0_auto_stream_in_0_valid = mag_split_auto_stream_out_1_valid; // @[LazyModule.scala 167:57]
  assign mag_mux_0_auto_stream_in_0_bits_data = mag_split_auto_stream_out_1_bits_data; // @[LazyModule.scala 167:57]
  assign mag_mux_0_auto_stream_in_0_bits_last = mag_split_auto_stream_out_1_bits_last; // @[LazyModule.scala 167:57]
  assign mag_mux_0_auto_stream_out_0_ready = buffer_2_auto_in_ready; // @[LazyModule.scala 167:57]
  assign mag_mux_1_clock = clock;
  assign mag_mux_1_reset = reset;
  assign mag_mux_1_auto_register_in_aw_valid = axi4buf_16_auto_out_aw_valid; // @[LazyModule.scala 167:31]
  assign mag_mux_1_auto_register_in_aw_bits_id = axi4buf_16_auto_out_aw_bits_id; // @[LazyModule.scala 167:31]
  assign mag_mux_1_auto_register_in_aw_bits_addr = axi4buf_16_auto_out_aw_bits_addr; // @[LazyModule.scala 167:31]
  assign mag_mux_1_auto_register_in_w_valid = axi4buf_16_auto_out_w_valid; // @[LazyModule.scala 167:31]
  assign mag_mux_1_auto_register_in_w_bits_data = axi4buf_16_auto_out_w_bits_data; // @[LazyModule.scala 167:31]
  assign mag_mux_1_auto_register_in_w_bits_strb = axi4buf_16_auto_out_w_bits_strb; // @[LazyModule.scala 167:31]
  assign mag_mux_1_auto_register_in_b_ready = axi4buf_16_auto_out_b_ready; // @[LazyModule.scala 167:31]
  assign mag_mux_1_auto_register_in_ar_valid = axi4buf_16_auto_out_ar_valid; // @[LazyModule.scala 167:31]
  assign mag_mux_1_auto_register_in_ar_bits_id = axi4buf_16_auto_out_ar_bits_id; // @[LazyModule.scala 167:31]
  assign mag_mux_1_auto_register_in_ar_bits_addr = axi4buf_16_auto_out_ar_bits_addr; // @[LazyModule.scala 167:31]
  assign mag_mux_1_auto_register_in_ar_bits_size = axi4buf_16_auto_out_ar_bits_size; // @[LazyModule.scala 167:31]
  assign mag_mux_1_auto_register_in_r_ready = axi4buf_16_auto_out_r_ready; // @[LazyModule.scala 167:31]
  assign mag_mux_1_auto_stream_in_valid = mag_split_auto_stream_out_0_valid; // @[LazyModule.scala 167:57]
  assign mag_mux_1_auto_stream_in_bits_data = mag_split_auto_stream_out_0_bits_data; // @[LazyModule.scala 167:57]
  assign mag_mux_1_auto_stream_in_bits_last = mag_split_auto_stream_out_0_bits_last; // @[LazyModule.scala 167:57]
  assign mag_mux_1_auto_stream_out_1_ready = buffer_3_auto_in_ready; // @[LazyModule.scala 167:57]
  assign acc_clock = clock;
  assign acc_reset = reset;
  assign acc_auto_bus_in_aw_valid = bus_auto_out_21_aw_valid; // @[LazyModule.scala 167:31]
  assign acc_auto_bus_in_aw_bits_id = bus_auto_out_21_aw_bits_id; // @[LazyModule.scala 167:31]
  assign acc_auto_bus_in_aw_bits_addr = bus_auto_out_21_aw_bits_addr; // @[LazyModule.scala 167:31]
  assign acc_auto_bus_in_aw_bits_size = bus_auto_out_21_aw_bits_size; // @[LazyModule.scala 167:31]
  assign acc_auto_bus_in_w_valid = bus_auto_out_21_w_valid; // @[LazyModule.scala 167:31]
  assign acc_auto_bus_in_w_bits_data = bus_auto_out_21_w_bits_data; // @[LazyModule.scala 167:31]
  assign acc_auto_bus_in_w_bits_strb = bus_auto_out_21_w_bits_strb; // @[LazyModule.scala 167:31]
  assign acc_auto_bus_in_w_bits_last = bus_auto_out_21_w_bits_last; // @[LazyModule.scala 167:31]
  assign acc_auto_bus_in_b_ready = bus_auto_out_21_b_ready; // @[LazyModule.scala 167:31]
  assign acc_auto_bus_in_ar_valid = bus_auto_out_21_ar_valid; // @[LazyModule.scala 167:31]
  assign acc_auto_bus_in_ar_bits_id = bus_auto_out_21_ar_bits_id; // @[LazyModule.scala 167:31]
  assign acc_auto_bus_in_ar_bits_addr = bus_auto_out_21_ar_bits_addr; // @[LazyModule.scala 167:31]
  assign acc_auto_bus_in_ar_bits_size = bus_auto_out_21_ar_bits_size; // @[LazyModule.scala 167:31]
  assign acc_auto_bus_in_r_ready = bus_auto_out_21_r_ready; // @[LazyModule.scala 167:31]
  assign acc_auto_dspQueue_stream_out_ready = widthAdapter_1_auto_in_ready; // @[LazyModule.scala 167:57]
  assign acc_auto_accumulator_slave_in_valid = buffer_2_auto_out_valid; // @[LazyModule.scala 167:31]
  assign acc_auto_accumulator_slave_in_bits_data = buffer_2_auto_out_bits_data; // @[LazyModule.scala 167:31]
  assign acc_auto_accumulator_slave_in_bits_last = buffer_2_auto_out_bits_last; // @[LazyModule.scala 167:31]
  assign widthAdapter_1_clock = clock;
  assign widthAdapter_1_reset = reset;
  assign widthAdapter_1_auto_in_valid = acc_auto_dspQueue_stream_out_valid; // @[LazyModule.scala 167:57]
  assign widthAdapter_1_auto_in_bits_data = acc_auto_dspQueue_stream_out_bits_data; // @[LazyModule.scala 167:57]
  assign widthAdapter_1_auto_in_bits_last = acc_auto_dspQueue_stream_out_bits_last; // @[LazyModule.scala 167:57]
  assign widthAdapter_1_auto_out_ready = acc_queue_auto_in_in_ready; // @[LazyModule.scala 167:57]
  assign acc_queue_clock = clock;
  assign acc_queue_reset = reset;
  assign acc_queue_auto_out_out_ready = out_mux_auto_stream_in_0_ready; // @[LazyModule.scala 167:57]
  assign acc_queue_auto_in_in_valid = widthAdapter_1_auto_out_valid; // @[LazyModule.scala 167:57]
  assign acc_queue_auto_in_in_bits_data = widthAdapter_1_auto_out_bits_data; // @[LazyModule.scala 167:57]
  assign acc_queue_auto_in_in_bits_last = widthAdapter_1_auto_out_bits_last; // @[LazyModule.scala 167:57]
  assign out_mux_clock = clock;
  assign out_mux_reset = reset;
  assign out_mux_auto_register_in_aw_valid = axi4buf_17_auto_out_aw_valid; // @[LazyModule.scala 167:31]
  assign out_mux_auto_register_in_aw_bits_id = axi4buf_17_auto_out_aw_bits_id; // @[LazyModule.scala 167:31]
  assign out_mux_auto_register_in_aw_bits_addr = axi4buf_17_auto_out_aw_bits_addr; // @[LazyModule.scala 167:31]
  assign out_mux_auto_register_in_w_valid = axi4buf_17_auto_out_w_valid; // @[LazyModule.scala 167:31]
  assign out_mux_auto_register_in_w_bits_data = axi4buf_17_auto_out_w_bits_data; // @[LazyModule.scala 167:31]
  assign out_mux_auto_register_in_w_bits_strb = axi4buf_17_auto_out_w_bits_strb; // @[LazyModule.scala 167:31]
  assign out_mux_auto_register_in_b_ready = axi4buf_17_auto_out_b_ready; // @[LazyModule.scala 167:31]
  assign out_mux_auto_register_in_ar_valid = axi4buf_17_auto_out_ar_valid; // @[LazyModule.scala 167:31]
  assign out_mux_auto_register_in_ar_bits_id = axi4buf_17_auto_out_ar_bits_id; // @[LazyModule.scala 167:31]
  assign out_mux_auto_register_in_ar_bits_addr = axi4buf_17_auto_out_ar_bits_addr; // @[LazyModule.scala 167:31]
  assign out_mux_auto_register_in_ar_bits_size = axi4buf_17_auto_out_ar_bits_size; // @[LazyModule.scala 167:31]
  assign out_mux_auto_register_in_r_ready = axi4buf_17_auto_out_r_ready; // @[LazyModule.scala 167:31]
  assign out_mux_auto_stream_in_6_valid = buffer_8_auto_out_valid; // @[LazyModule.scala 167:31]
  assign out_mux_auto_stream_in_6_bits_data = buffer_8_auto_out_bits_data; // @[LazyModule.scala 167:31]
  assign out_mux_auto_stream_in_6_bits_last = buffer_8_auto_out_bits_last; // @[LazyModule.scala 167:31]
  assign out_mux_auto_stream_in_5_valid = buffer_7_auto_out_valid; // @[LazyModule.scala 167:31]
  assign out_mux_auto_stream_in_5_bits_data = buffer_7_auto_out_bits_data; // @[LazyModule.scala 167:31]
  assign out_mux_auto_stream_in_5_bits_last = buffer_7_auto_out_bits_last; // @[LazyModule.scala 167:31]
  assign out_mux_auto_stream_in_4_valid = buffer_6_auto_out_valid; // @[LazyModule.scala 167:31]
  assign out_mux_auto_stream_in_4_bits_data = buffer_6_auto_out_bits_data; // @[LazyModule.scala 167:31]
  assign out_mux_auto_stream_in_4_bits_last = buffer_6_auto_out_bits_last; // @[LazyModule.scala 167:31]
  assign out_mux_auto_stream_in_3_valid = buffer_5_auto_out_valid; // @[LazyModule.scala 167:31]
  assign out_mux_auto_stream_in_3_bits_data = buffer_5_auto_out_bits_data; // @[LazyModule.scala 167:31]
  assign out_mux_auto_stream_in_3_bits_last = buffer_5_auto_out_bits_last; // @[LazyModule.scala 167:31]
  assign out_mux_auto_stream_in_2_valid = buffer_4_auto_out_valid; // @[LazyModule.scala 167:31]
  assign out_mux_auto_stream_in_2_bits_data = buffer_4_auto_out_bits_data; // @[LazyModule.scala 167:31]
  assign out_mux_auto_stream_in_2_bits_last = buffer_4_auto_out_bits_last; // @[LazyModule.scala 167:31]
  assign out_mux_auto_stream_in_1_valid = buffer_3_auto_out_valid; // @[LazyModule.scala 167:31]
  assign out_mux_auto_stream_in_1_bits_data = buffer_3_auto_out_bits_data; // @[LazyModule.scala 167:31]
  assign out_mux_auto_stream_in_1_bits_last = buffer_3_auto_out_bits_last; // @[LazyModule.scala 167:31]
  assign out_mux_auto_stream_in_0_valid = acc_queue_auto_out_out_valid; // @[LazyModule.scala 167:57]
  assign out_mux_auto_stream_in_0_bits_data = acc_queue_auto_out_out_bits_data; // @[LazyModule.scala 167:57]
  assign out_mux_auto_stream_in_0_bits_last = acc_queue_auto_out_out_bits_last; // @[LazyModule.scala 167:57]
  assign out_mux_auto_stream_out_1_ready = uTx_queue_auto_in_in_ready; // @[LazyModule.scala 167:57]
  assign out_mux_auto_stream_out_0_ready = buffer_9_auto_in_ready; // @[LazyModule.scala 167:57]
  assign out_split_clock = clock;
  assign out_split_reset = reset;
  assign out_split_auto_mem_in_aw_valid = axi4buf_18_auto_out_aw_valid; // @[LazyModule.scala 167:31]
  assign out_split_auto_mem_in_aw_bits_id = axi4buf_18_auto_out_aw_bits_id; // @[LazyModule.scala 167:31]
  assign out_split_auto_mem_in_aw_bits_addr = axi4buf_18_auto_out_aw_bits_addr; // @[LazyModule.scala 167:31]
  assign out_split_auto_mem_in_w_valid = axi4buf_18_auto_out_w_valid; // @[LazyModule.scala 167:31]
  assign out_split_auto_mem_in_w_bits_data = axi4buf_18_auto_out_w_bits_data; // @[LazyModule.scala 167:31]
  assign out_split_auto_mem_in_w_bits_strb = axi4buf_18_auto_out_w_bits_strb; // @[LazyModule.scala 167:31]
  assign out_split_auto_mem_in_b_ready = axi4buf_18_auto_out_b_ready; // @[LazyModule.scala 167:31]
  assign out_split_auto_mem_in_ar_valid = axi4buf_18_auto_out_ar_valid; // @[LazyModule.scala 167:31]
  assign out_split_auto_mem_in_ar_bits_id = axi4buf_18_auto_out_ar_bits_id; // @[LazyModule.scala 167:31]
  assign out_split_auto_mem_in_ar_bits_addr = axi4buf_18_auto_out_ar_bits_addr; // @[LazyModule.scala 167:31]
  assign out_split_auto_mem_in_ar_bits_size = axi4buf_18_auto_out_ar_bits_size; // @[LazyModule.scala 167:31]
  assign out_split_auto_mem_in_r_ready = axi4buf_18_auto_out_r_ready; // @[LazyModule.scala 167:31]
  assign out_split_auto_stream_in_valid = out_queue_auto_out_out_valid; // @[LazyModule.scala 167:31]
  assign out_split_auto_stream_in_bits_data = out_queue_auto_out_out_bits_data; // @[LazyModule.scala 167:31]
  assign out_split_auto_stream_in_bits_last = out_queue_auto_out_out_bits_last; // @[LazyModule.scala 167:31]
  assign out_split_auto_stream_out_ready = widthAdapter_2_auto_in_ready; // @[LazyModule.scala 167:57]
  assign out_queue_clock = clock;
  assign out_queue_reset = reset;
  assign out_queue_auto_out_out_ready = out_split_auto_stream_in_ready; // @[LazyModule.scala 167:31]
  assign out_queue_auto_in_in_valid = buffer_9_auto_out_valid; // @[LazyModule.scala 167:31]
  assign out_queue_auto_in_in_bits_data = buffer_9_auto_out_bits_data; // @[LazyModule.scala 167:31]
  assign out_queue_auto_in_in_bits_last = buffer_9_auto_out_bits_last; // @[LazyModule.scala 167:31]
  assign widthAdapter_2_clock = clock;
  assign widthAdapter_2_reset = reset;
  assign widthAdapter_2_auto_in_valid = out_split_auto_stream_out_valid; // @[LazyModule.scala 167:57]
  assign widthAdapter_2_auto_in_bits_data = out_split_auto_stream_out_bits_data; // @[LazyModule.scala 167:57]
  assign widthAdapter_2_auto_in_bits_last = out_split_auto_stream_out_bits_last; // @[LazyModule.scala 167:57]
  assign widthAdapter_2_auto_out_ready = converter_1_auto_in_ready; // @[LazyModule.scala 167:57]
  assign uTx_queue_clock = clock;
  assign uTx_queue_reset = reset;
  assign uTx_queue_auto_out_out_ready = widthAdapter_3_auto_in_ready; // @[LazyModule.scala 167:57]
  assign uTx_queue_auto_in_in_valid = out_mux_auto_stream_out_1_valid; // @[LazyModule.scala 167:57]
  assign uTx_queue_auto_in_in_bits_data = out_mux_auto_stream_out_1_bits_data; // @[LazyModule.scala 167:57]
  assign uTx_queue_auto_in_in_bits_last = out_mux_auto_stream_out_1_bits_last; // @[LazyModule.scala 167:57]
  assign widthAdapter_3_clock = clock;
  assign widthAdapter_3_reset = reset;
  assign widthAdapter_3_auto_in_valid = uTx_queue_auto_out_out_valid; // @[LazyModule.scala 167:57]
  assign widthAdapter_3_auto_in_bits_data = uTx_queue_auto_out_out_bits_data; // @[LazyModule.scala 167:57]
  assign widthAdapter_3_auto_in_bits_last = uTx_queue_auto_out_out_bits_last; // @[LazyModule.scala 167:57]
  assign widthAdapter_3_auto_out_ready = uart_auto_in_in_ready; // @[LazyModule.scala 167:57]
  assign widthAdapter_4_clock = clock;
  assign widthAdapter_4_reset = reset;
  assign widthAdapter_4_auto_in_valid = uart_auto_out_out_valid; // @[LazyModule.scala 167:31]
  assign widthAdapter_4_auto_in_bits_data = uart_auto_out_out_bits_data; // @[LazyModule.scala 167:31]
  assign widthAdapter_4_auto_in_bits_last = 1'h0; // @[LazyModule.scala 167:31]
  assign widthAdapter_4_auto_out_ready = uRx_split_auto_stream_in_ready; // @[LazyModule.scala 167:57]
  assign uRx_split_clock = clock;
  assign uRx_split_reset = reset;
  assign uRx_split_auto_mem_in_aw_valid = axi4buf_20_auto_out_aw_valid; // @[LazyModule.scala 167:31]
  assign uRx_split_auto_mem_in_aw_bits_id = axi4buf_20_auto_out_aw_bits_id; // @[LazyModule.scala 167:31]
  assign uRx_split_auto_mem_in_aw_bits_addr = axi4buf_20_auto_out_aw_bits_addr; // @[LazyModule.scala 167:31]
  assign uRx_split_auto_mem_in_w_valid = axi4buf_20_auto_out_w_valid; // @[LazyModule.scala 167:31]
  assign uRx_split_auto_mem_in_w_bits_data = axi4buf_20_auto_out_w_bits_data; // @[LazyModule.scala 167:31]
  assign uRx_split_auto_mem_in_w_bits_strb = axi4buf_20_auto_out_w_bits_strb; // @[LazyModule.scala 167:31]
  assign uRx_split_auto_mem_in_b_ready = axi4buf_20_auto_out_b_ready; // @[LazyModule.scala 167:31]
  assign uRx_split_auto_mem_in_ar_valid = axi4buf_20_auto_out_ar_valid; // @[LazyModule.scala 167:31]
  assign uRx_split_auto_mem_in_ar_bits_id = axi4buf_20_auto_out_ar_bits_id; // @[LazyModule.scala 167:31]
  assign uRx_split_auto_mem_in_ar_bits_addr = axi4buf_20_auto_out_ar_bits_addr; // @[LazyModule.scala 167:31]
  assign uRx_split_auto_mem_in_ar_bits_size = axi4buf_20_auto_out_ar_bits_size; // @[LazyModule.scala 167:31]
  assign uRx_split_auto_mem_in_r_ready = axi4buf_20_auto_out_r_ready; // @[LazyModule.scala 167:31]
  assign uRx_split_auto_stream_in_valid = widthAdapter_4_auto_out_valid; // @[LazyModule.scala 167:57]
  assign uRx_split_auto_stream_in_bits_data = widthAdapter_4_auto_out_bits_data; // @[LazyModule.scala 167:57]
  assign uRx_split_auto_stream_in_bits_last = widthAdapter_4_auto_out_bits_last; // @[LazyModule.scala 167:57]
  assign uRx_split_auto_stream_out_4_ready = buffer_8_auto_in_ready; // @[LazyModule.scala 167:57]
  assign uRx_split_auto_stream_out_3_ready = mag_mux_0_auto_stream_in_2_ready; // @[LazyModule.scala 167:31]
  assign uRx_split_auto_stream_out_2_ready = fft_mux_0_auto_stream_in_2_ready; // @[LazyModule.scala 167:31]
  assign uRx_split_auto_stream_out_1_ready = nco_mux_0_auto_stream_in_2_ready; // @[LazyModule.scala 167:31]
  assign uRx_split_auto_stream_out_0_ready = plfg_mux_0_auto_stream_in_2_ready; // @[LazyModule.scala 167:31]
  assign uart_clock = clock;
  assign uart_reset = reset;
  assign uart_auto_mem_in_aw_valid = axi4buf_19_auto_out_aw_valid; // @[LazyModule.scala 167:31]
  assign uart_auto_mem_in_aw_bits_id = axi4buf_19_auto_out_aw_bits_id; // @[LazyModule.scala 167:31]
  assign uart_auto_mem_in_aw_bits_addr = axi4buf_19_auto_out_aw_bits_addr; // @[LazyModule.scala 167:31]
  assign uart_auto_mem_in_w_valid = axi4buf_19_auto_out_w_valid; // @[LazyModule.scala 167:31]
  assign uart_auto_mem_in_w_bits_data = axi4buf_19_auto_out_w_bits_data; // @[LazyModule.scala 167:31]
  assign uart_auto_mem_in_w_bits_strb = axi4buf_19_auto_out_w_bits_strb; // @[LazyModule.scala 167:31]
  assign uart_auto_mem_in_b_ready = axi4buf_19_auto_out_b_ready; // @[LazyModule.scala 167:31]
  assign uart_auto_mem_in_ar_valid = axi4buf_19_auto_out_ar_valid; // @[LazyModule.scala 167:31]
  assign uart_auto_mem_in_ar_bits_id = axi4buf_19_auto_out_ar_bits_id; // @[LazyModule.scala 167:31]
  assign uart_auto_mem_in_ar_bits_addr = axi4buf_19_auto_out_ar_bits_addr; // @[LazyModule.scala 167:31]
  assign uart_auto_mem_in_ar_bits_size = axi4buf_19_auto_out_ar_bits_size; // @[LazyModule.scala 167:31]
  assign uart_auto_mem_in_r_ready = axi4buf_19_auto_out_r_ready; // @[LazyModule.scala 167:31]
  assign uart_auto_in_in_valid = widthAdapter_3_auto_out_valid; // @[LazyModule.scala 167:57]
  assign uart_auto_in_in_bits_data = widthAdapter_3_auto_out_bits_data; // @[LazyModule.scala 167:57]
  assign uart_auto_out_out_ready = widthAdapter_4_auto_in_ready; // @[LazyModule.scala 167:31]
  assign uart_io_rxd = uRx; // @[SpectrometerTestWithoutLA.scala 213:24]
  assign bus_clock = clock;
  assign bus_reset = reset;
  assign bus_auto_in_aw_valid = converter_auto_out_aw_valid; // @[LazyModule.scala 167:31]
  assign bus_auto_in_aw_bits_id = converter_auto_out_aw_bits_id; // @[LazyModule.scala 167:31]
  assign bus_auto_in_aw_bits_addr = converter_auto_out_aw_bits_addr; // @[LazyModule.scala 167:31]
  assign bus_auto_in_aw_bits_size = converter_auto_out_aw_bits_size; // @[LazyModule.scala 167:31]
  assign bus_auto_in_w_valid = converter_auto_out_w_valid; // @[LazyModule.scala 167:31]
  assign bus_auto_in_w_bits_data = converter_auto_out_w_bits_data; // @[LazyModule.scala 167:31]
  assign bus_auto_in_w_bits_strb = converter_auto_out_w_bits_strb; // @[LazyModule.scala 167:31]
  assign bus_auto_in_w_bits_last = converter_auto_out_w_bits_last; // @[LazyModule.scala 167:31]
  assign bus_auto_in_b_ready = converter_auto_out_b_ready; // @[LazyModule.scala 167:31]
  assign bus_auto_in_ar_valid = converter_auto_out_ar_valid; // @[LazyModule.scala 167:31]
  assign bus_auto_in_ar_bits_id = converter_auto_out_ar_bits_id; // @[LazyModule.scala 167:31]
  assign bus_auto_in_ar_bits_addr = converter_auto_out_ar_bits_addr; // @[LazyModule.scala 167:31]
  assign bus_auto_in_ar_bits_size = converter_auto_out_ar_bits_size; // @[LazyModule.scala 167:31]
  assign bus_auto_in_r_ready = converter_auto_out_r_ready; // @[LazyModule.scala 167:31]
  assign bus_auto_out_21_aw_ready = acc_auto_bus_in_aw_ready; // @[LazyModule.scala 167:31]
  assign bus_auto_out_21_w_ready = acc_auto_bus_in_w_ready; // @[LazyModule.scala 167:31]
  assign bus_auto_out_21_b_valid = acc_auto_bus_in_b_valid; // @[LazyModule.scala 167:31]
  assign bus_auto_out_21_b_bits_resp = acc_auto_bus_in_b_bits_resp; // @[LazyModule.scala 167:31]
  assign bus_auto_out_21_ar_ready = acc_auto_bus_in_ar_ready; // @[LazyModule.scala 167:31]
  assign bus_auto_out_21_r_valid = acc_auto_bus_in_r_valid; // @[LazyModule.scala 167:31]
  assign bus_auto_out_21_r_bits_data = acc_auto_bus_in_r_bits_data; // @[LazyModule.scala 167:31]
  assign bus_auto_out_21_r_bits_resp = acc_auto_bus_in_r_bits_resp; // @[LazyModule.scala 167:31]
  assign bus_auto_out_21_r_bits_last = acc_auto_bus_in_r_bits_last; // @[LazyModule.scala 167:31]
  assign bus_auto_out_20_aw_ready = axi4buf_20_auto_in_aw_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_20_w_ready = axi4buf_20_auto_in_w_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_20_b_valid = axi4buf_20_auto_in_b_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_20_b_bits_id = axi4buf_20_auto_in_b_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_20_b_bits_resp = axi4buf_20_auto_in_b_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_20_ar_ready = axi4buf_20_auto_in_ar_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_20_r_valid = axi4buf_20_auto_in_r_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_20_r_bits_id = axi4buf_20_auto_in_r_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_20_r_bits_data = axi4buf_20_auto_in_r_bits_data; // @[LazyModule.scala 167:57]
  assign bus_auto_out_20_r_bits_resp = axi4buf_20_auto_in_r_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_20_r_bits_last = axi4buf_20_auto_in_r_bits_last; // @[LazyModule.scala 167:57]
  assign bus_auto_out_19_aw_ready = axi4buf_19_auto_in_aw_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_19_w_ready = axi4buf_19_auto_in_w_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_19_b_valid = axi4buf_19_auto_in_b_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_19_b_bits_id = axi4buf_19_auto_in_b_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_19_b_bits_resp = axi4buf_19_auto_in_b_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_19_ar_ready = axi4buf_19_auto_in_ar_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_19_r_valid = axi4buf_19_auto_in_r_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_19_r_bits_id = axi4buf_19_auto_in_r_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_19_r_bits_data = axi4buf_19_auto_in_r_bits_data; // @[LazyModule.scala 167:57]
  assign bus_auto_out_19_r_bits_resp = axi4buf_19_auto_in_r_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_19_r_bits_last = axi4buf_19_auto_in_r_bits_last; // @[LazyModule.scala 167:57]
  assign bus_auto_out_18_aw_ready = axi4buf_18_auto_in_aw_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_18_w_ready = axi4buf_18_auto_in_w_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_18_b_valid = axi4buf_18_auto_in_b_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_18_b_bits_id = axi4buf_18_auto_in_b_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_18_b_bits_resp = axi4buf_18_auto_in_b_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_18_ar_ready = axi4buf_18_auto_in_ar_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_18_r_valid = axi4buf_18_auto_in_r_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_18_r_bits_id = axi4buf_18_auto_in_r_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_18_r_bits_data = axi4buf_18_auto_in_r_bits_data; // @[LazyModule.scala 167:57]
  assign bus_auto_out_18_r_bits_resp = axi4buf_18_auto_in_r_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_18_r_bits_last = axi4buf_18_auto_in_r_bits_last; // @[LazyModule.scala 167:57]
  assign bus_auto_out_17_aw_ready = axi4buf_17_auto_in_aw_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_17_w_ready = axi4buf_17_auto_in_w_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_17_b_valid = axi4buf_17_auto_in_b_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_17_b_bits_id = axi4buf_17_auto_in_b_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_17_b_bits_resp = axi4buf_17_auto_in_b_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_17_ar_ready = axi4buf_17_auto_in_ar_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_17_r_valid = axi4buf_17_auto_in_r_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_17_r_bits_id = axi4buf_17_auto_in_r_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_17_r_bits_data = axi4buf_17_auto_in_r_bits_data; // @[LazyModule.scala 167:57]
  assign bus_auto_out_17_r_bits_resp = axi4buf_17_auto_in_r_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_17_r_bits_last = axi4buf_17_auto_in_r_bits_last; // @[LazyModule.scala 167:57]
  assign bus_auto_out_16_aw_ready = axi4buf_16_auto_in_aw_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_16_w_ready = axi4buf_16_auto_in_w_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_16_b_valid = axi4buf_16_auto_in_b_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_16_b_bits_id = axi4buf_16_auto_in_b_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_16_b_bits_resp = axi4buf_16_auto_in_b_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_16_ar_ready = axi4buf_16_auto_in_ar_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_16_r_valid = axi4buf_16_auto_in_r_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_16_r_bits_id = axi4buf_16_auto_in_r_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_16_r_bits_data = axi4buf_16_auto_in_r_bits_data; // @[LazyModule.scala 167:57]
  assign bus_auto_out_16_r_bits_resp = axi4buf_16_auto_in_r_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_16_r_bits_last = axi4buf_16_auto_in_r_bits_last; // @[LazyModule.scala 167:57]
  assign bus_auto_out_15_aw_ready = axi4buf_15_auto_in_aw_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_15_w_ready = axi4buf_15_auto_in_w_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_15_b_valid = axi4buf_15_auto_in_b_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_15_b_bits_id = axi4buf_15_auto_in_b_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_15_b_bits_resp = axi4buf_15_auto_in_b_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_15_ar_ready = axi4buf_15_auto_in_ar_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_15_r_valid = axi4buf_15_auto_in_r_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_15_r_bits_id = axi4buf_15_auto_in_r_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_15_r_bits_data = axi4buf_15_auto_in_r_bits_data; // @[LazyModule.scala 167:57]
  assign bus_auto_out_15_r_bits_resp = axi4buf_15_auto_in_r_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_15_r_bits_last = axi4buf_15_auto_in_r_bits_last; // @[LazyModule.scala 167:57]
  assign bus_auto_out_14_aw_ready = axi4buf_14_auto_in_aw_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_14_w_ready = axi4buf_14_auto_in_w_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_14_b_valid = axi4buf_14_auto_in_b_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_14_b_bits_id = axi4buf_14_auto_in_b_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_14_b_bits_resp = axi4buf_14_auto_in_b_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_14_ar_ready = axi4buf_14_auto_in_ar_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_14_r_valid = axi4buf_14_auto_in_r_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_14_r_bits_id = axi4buf_14_auto_in_r_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_14_r_bits_data = axi4buf_14_auto_in_r_bits_data; // @[LazyModule.scala 167:57]
  assign bus_auto_out_14_r_bits_resp = axi4buf_14_auto_in_r_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_14_r_bits_last = axi4buf_14_auto_in_r_bits_last; // @[LazyModule.scala 167:57]
  assign bus_auto_out_13_aw_ready = axi4buf_13_auto_in_aw_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_13_w_ready = axi4buf_13_auto_in_w_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_13_b_valid = axi4buf_13_auto_in_b_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_13_b_bits_id = axi4buf_13_auto_in_b_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_13_b_bits_resp = axi4buf_13_auto_in_b_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_13_ar_ready = axi4buf_13_auto_in_ar_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_13_r_valid = axi4buf_13_auto_in_r_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_13_r_bits_id = axi4buf_13_auto_in_r_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_13_r_bits_data = axi4buf_13_auto_in_r_bits_data; // @[LazyModule.scala 167:57]
  assign bus_auto_out_13_r_bits_resp = axi4buf_13_auto_in_r_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_13_r_bits_last = axi4buf_13_auto_in_r_bits_last; // @[LazyModule.scala 167:57]
  assign bus_auto_out_12_aw_ready = axi4buf_12_auto_in_aw_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_12_w_ready = axi4buf_12_auto_in_w_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_12_b_valid = axi4buf_12_auto_in_b_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_12_b_bits_id = axi4buf_12_auto_in_b_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_12_b_bits_resp = axi4buf_12_auto_in_b_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_12_ar_ready = axi4buf_12_auto_in_ar_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_12_r_valid = axi4buf_12_auto_in_r_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_12_r_bits_id = axi4buf_12_auto_in_r_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_12_r_bits_data = axi4buf_12_auto_in_r_bits_data; // @[LazyModule.scala 167:57]
  assign bus_auto_out_12_r_bits_resp = axi4buf_12_auto_in_r_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_12_r_bits_last = axi4buf_12_auto_in_r_bits_last; // @[LazyModule.scala 167:57]
  assign bus_auto_out_11_aw_ready = axi4buf_11_auto_in_aw_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_11_w_ready = axi4buf_11_auto_in_w_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_11_b_valid = axi4buf_11_auto_in_b_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_11_b_bits_id = axi4buf_11_auto_in_b_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_11_b_bits_resp = axi4buf_11_auto_in_b_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_11_ar_ready = axi4buf_11_auto_in_ar_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_11_r_valid = axi4buf_11_auto_in_r_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_11_r_bits_id = axi4buf_11_auto_in_r_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_11_r_bits_data = axi4buf_11_auto_in_r_bits_data; // @[LazyModule.scala 167:57]
  assign bus_auto_out_11_r_bits_resp = axi4buf_11_auto_in_r_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_11_r_bits_last = axi4buf_11_auto_in_r_bits_last; // @[LazyModule.scala 167:57]
  assign bus_auto_out_10_aw_ready = axi4buf_10_auto_in_aw_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_10_w_ready = axi4buf_10_auto_in_w_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_10_b_valid = axi4buf_10_auto_in_b_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_10_b_bits_id = axi4buf_10_auto_in_b_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_10_b_bits_resp = axi4buf_10_auto_in_b_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_10_ar_ready = axi4buf_10_auto_in_ar_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_10_r_valid = axi4buf_10_auto_in_r_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_10_r_bits_id = axi4buf_10_auto_in_r_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_10_r_bits_data = axi4buf_10_auto_in_r_bits_data; // @[LazyModule.scala 167:57]
  assign bus_auto_out_10_r_bits_resp = axi4buf_10_auto_in_r_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_10_r_bits_last = axi4buf_10_auto_in_r_bits_last; // @[LazyModule.scala 167:57]
  assign bus_auto_out_9_aw_ready = axi4buf_9_auto_in_aw_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_9_w_ready = axi4buf_9_auto_in_w_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_9_b_valid = axi4buf_9_auto_in_b_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_9_b_bits_id = axi4buf_9_auto_in_b_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_9_b_bits_resp = axi4buf_9_auto_in_b_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_9_ar_ready = axi4buf_9_auto_in_ar_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_9_r_valid = axi4buf_9_auto_in_r_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_9_r_bits_id = axi4buf_9_auto_in_r_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_9_r_bits_data = axi4buf_9_auto_in_r_bits_data; // @[LazyModule.scala 167:57]
  assign bus_auto_out_9_r_bits_resp = axi4buf_9_auto_in_r_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_9_r_bits_last = axi4buf_9_auto_in_r_bits_last; // @[LazyModule.scala 167:57]
  assign bus_auto_out_8_aw_ready = axi4buf_8_auto_in_aw_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_8_w_ready = axi4buf_8_auto_in_w_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_8_b_valid = axi4buf_8_auto_in_b_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_8_b_bits_id = axi4buf_8_auto_in_b_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_8_b_bits_resp = axi4buf_8_auto_in_b_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_8_ar_ready = axi4buf_8_auto_in_ar_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_8_r_valid = axi4buf_8_auto_in_r_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_8_r_bits_id = axi4buf_8_auto_in_r_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_8_r_bits_data = axi4buf_8_auto_in_r_bits_data; // @[LazyModule.scala 167:57]
  assign bus_auto_out_8_r_bits_resp = axi4buf_8_auto_in_r_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_8_r_bits_last = axi4buf_8_auto_in_r_bits_last; // @[LazyModule.scala 167:57]
  assign bus_auto_out_7_aw_ready = axi4buf_7_auto_in_aw_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_7_w_ready = axi4buf_7_auto_in_w_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_7_b_valid = axi4buf_7_auto_in_b_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_7_b_bits_id = axi4buf_7_auto_in_b_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_7_b_bits_resp = axi4buf_7_auto_in_b_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_7_ar_ready = axi4buf_7_auto_in_ar_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_7_r_valid = axi4buf_7_auto_in_r_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_7_r_bits_id = axi4buf_7_auto_in_r_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_7_r_bits_data = axi4buf_7_auto_in_r_bits_data; // @[LazyModule.scala 167:57]
  assign bus_auto_out_7_r_bits_resp = axi4buf_7_auto_in_r_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_7_r_bits_last = axi4buf_7_auto_in_r_bits_last; // @[LazyModule.scala 167:57]
  assign bus_auto_out_6_aw_ready = axi4buf_6_auto_in_aw_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_6_w_ready = axi4buf_6_auto_in_w_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_6_b_valid = axi4buf_6_auto_in_b_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_6_b_bits_id = axi4buf_6_auto_in_b_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_6_b_bits_resp = axi4buf_6_auto_in_b_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_6_ar_ready = axi4buf_6_auto_in_ar_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_6_r_valid = axi4buf_6_auto_in_r_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_6_r_bits_id = axi4buf_6_auto_in_r_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_6_r_bits_data = axi4buf_6_auto_in_r_bits_data; // @[LazyModule.scala 167:57]
  assign bus_auto_out_6_r_bits_resp = axi4buf_6_auto_in_r_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_6_r_bits_last = axi4buf_6_auto_in_r_bits_last; // @[LazyModule.scala 167:57]
  assign bus_auto_out_5_aw_ready = axi4buf_5_auto_in_aw_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_5_w_ready = axi4buf_5_auto_in_w_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_5_b_valid = axi4buf_5_auto_in_b_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_5_b_bits_id = axi4buf_5_auto_in_b_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_5_b_bits_resp = axi4buf_5_auto_in_b_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_5_ar_ready = axi4buf_5_auto_in_ar_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_5_r_valid = axi4buf_5_auto_in_r_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_5_r_bits_id = axi4buf_5_auto_in_r_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_5_r_bits_data = axi4buf_5_auto_in_r_bits_data; // @[LazyModule.scala 167:57]
  assign bus_auto_out_5_r_bits_resp = axi4buf_5_auto_in_r_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_5_r_bits_last = axi4buf_5_auto_in_r_bits_last; // @[LazyModule.scala 167:57]
  assign bus_auto_out_4_aw_ready = axi4buf_4_auto_in_aw_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_4_w_ready = axi4buf_4_auto_in_w_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_4_b_valid = axi4buf_4_auto_in_b_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_4_b_bits_id = axi4buf_4_auto_in_b_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_4_b_bits_resp = axi4buf_4_auto_in_b_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_4_ar_ready = axi4buf_4_auto_in_ar_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_4_r_valid = axi4buf_4_auto_in_r_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_4_r_bits_id = axi4buf_4_auto_in_r_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_4_r_bits_data = axi4buf_4_auto_in_r_bits_data; // @[LazyModule.scala 167:57]
  assign bus_auto_out_4_r_bits_resp = axi4buf_4_auto_in_r_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_4_r_bits_last = axi4buf_4_auto_in_r_bits_last; // @[LazyModule.scala 167:57]
  assign bus_auto_out_3_aw_ready = axi4buf_3_auto_in_aw_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_3_w_ready = axi4buf_3_auto_in_w_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_3_b_valid = axi4buf_3_auto_in_b_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_3_b_bits_id = axi4buf_3_auto_in_b_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_3_b_bits_resp = axi4buf_3_auto_in_b_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_3_ar_ready = axi4buf_3_auto_in_ar_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_3_r_valid = axi4buf_3_auto_in_r_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_3_r_bits_id = axi4buf_3_auto_in_r_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_3_r_bits_data = axi4buf_3_auto_in_r_bits_data; // @[LazyModule.scala 167:57]
  assign bus_auto_out_3_r_bits_resp = axi4buf_3_auto_in_r_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_3_r_bits_last = axi4buf_3_auto_in_r_bits_last; // @[LazyModule.scala 167:57]
  assign bus_auto_out_2_aw_ready = axi4buf_2_auto_in_aw_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_2_w_ready = axi4buf_2_auto_in_w_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_2_b_valid = axi4buf_2_auto_in_b_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_2_b_bits_id = axi4buf_2_auto_in_b_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_2_b_bits_resp = axi4buf_2_auto_in_b_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_2_ar_ready = axi4buf_2_auto_in_ar_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_2_r_valid = axi4buf_2_auto_in_r_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_2_r_bits_id = axi4buf_2_auto_in_r_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_2_r_bits_data = axi4buf_2_auto_in_r_bits_data; // @[LazyModule.scala 167:57]
  assign bus_auto_out_2_r_bits_resp = axi4buf_2_auto_in_r_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_2_r_bits_last = axi4buf_2_auto_in_r_bits_last; // @[LazyModule.scala 167:57]
  assign bus_auto_out_1_aw_ready = axi4buf_1_auto_in_aw_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_1_w_ready = axi4buf_1_auto_in_w_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_1_b_valid = axi4buf_1_auto_in_b_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_1_b_bits_id = axi4buf_1_auto_in_b_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_1_b_bits_resp = axi4buf_1_auto_in_b_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_1_ar_ready = axi4buf_1_auto_in_ar_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_1_r_valid = axi4buf_1_auto_in_r_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_1_r_bits_id = axi4buf_1_auto_in_r_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_1_r_bits_data = axi4buf_1_auto_in_r_bits_data; // @[LazyModule.scala 167:57]
  assign bus_auto_out_1_r_bits_resp = axi4buf_1_auto_in_r_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_1_r_bits_last = axi4buf_1_auto_in_r_bits_last; // @[LazyModule.scala 167:57]
  assign bus_auto_out_0_aw_ready = axi4buf_auto_in_aw_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_0_w_ready = axi4buf_auto_in_w_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_0_b_valid = axi4buf_auto_in_b_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_0_b_bits_id = axi4buf_auto_in_b_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_0_b_bits_resp = axi4buf_auto_in_b_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_0_ar_ready = axi4buf_auto_in_ar_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_0_r_valid = axi4buf_auto_in_r_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_0_r_bits_id = axi4buf_auto_in_r_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_0_r_bits_data = axi4buf_auto_in_r_bits_data; // @[LazyModule.scala 167:57]
  assign bus_auto_out_0_r_bits_resp = axi4buf_auto_in_r_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_0_r_bits_last = axi4buf_auto_in_r_bits_last; // @[LazyModule.scala 167:57]
  assign axi4buf_clock = clock;
  assign axi4buf_reset = reset;
  assign axi4buf_auto_in_aw_valid = bus_auto_out_0_aw_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_auto_in_aw_bits_id = bus_auto_out_0_aw_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_auto_in_aw_bits_addr = bus_auto_out_0_aw_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_auto_in_aw_bits_size = bus_auto_out_0_aw_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_auto_in_w_valid = bus_auto_out_0_w_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_auto_in_w_bits_data = bus_auto_out_0_w_bits_data; // @[LazyModule.scala 167:57]
  assign axi4buf_auto_in_w_bits_strb = bus_auto_out_0_w_bits_strb; // @[LazyModule.scala 167:57]
  assign axi4buf_auto_in_w_bits_last = bus_auto_out_0_w_bits_last; // @[LazyModule.scala 167:57]
  assign axi4buf_auto_in_b_ready = bus_auto_out_0_b_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_auto_in_ar_valid = bus_auto_out_0_ar_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_auto_in_ar_bits_id = bus_auto_out_0_ar_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_auto_in_ar_bits_addr = bus_auto_out_0_ar_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_auto_in_ar_bits_size = bus_auto_out_0_ar_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_auto_in_r_ready = bus_auto_out_0_r_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_auto_out_aw_ready = in_split_auto_mem_in_aw_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_auto_out_w_ready = in_split_auto_mem_in_w_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_auto_out_b_valid = in_split_auto_mem_in_b_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_auto_out_b_bits_id = in_split_auto_mem_in_b_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_auto_out_b_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_auto_out_ar_ready = in_split_auto_mem_in_ar_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_auto_out_r_valid = in_split_auto_mem_in_r_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_auto_out_r_bits_id = in_split_auto_mem_in_r_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_auto_out_r_bits_data = in_split_auto_mem_in_r_bits_data; // @[LazyModule.scala 167:31]
  assign axi4buf_auto_out_r_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_auto_out_r_bits_last = 1'h1; // @[LazyModule.scala 167:31]
  assign axi4buf_1_clock = clock;
  assign axi4buf_1_reset = reset;
  assign axi4buf_1_auto_in_aw_valid = bus_auto_out_1_aw_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_1_auto_in_aw_bits_id = bus_auto_out_1_aw_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_1_auto_in_aw_bits_addr = bus_auto_out_1_aw_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_1_auto_in_aw_bits_size = bus_auto_out_1_aw_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_1_auto_in_w_valid = bus_auto_out_1_w_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_1_auto_in_w_bits_data = bus_auto_out_1_w_bits_data; // @[LazyModule.scala 167:57]
  assign axi4buf_1_auto_in_w_bits_strb = bus_auto_out_1_w_bits_strb; // @[LazyModule.scala 167:57]
  assign axi4buf_1_auto_in_w_bits_last = bus_auto_out_1_w_bits_last; // @[LazyModule.scala 167:57]
  assign axi4buf_1_auto_in_b_ready = bus_auto_out_1_b_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_1_auto_in_ar_valid = bus_auto_out_1_ar_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_1_auto_in_ar_bits_id = bus_auto_out_1_ar_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_1_auto_in_ar_bits_addr = bus_auto_out_1_ar_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_1_auto_in_ar_bits_size = bus_auto_out_1_ar_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_1_auto_in_r_ready = bus_auto_out_1_r_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_1_auto_out_aw_ready = plfg_auto_mem_in_aw_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_1_auto_out_w_ready = plfg_auto_mem_in_w_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_1_auto_out_b_valid = plfg_auto_mem_in_b_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_1_auto_out_b_bits_id = 1'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_1_auto_out_b_bits_resp = plfg_auto_mem_in_b_bits_resp; // @[LazyModule.scala 167:31]
  assign axi4buf_1_auto_out_ar_ready = plfg_auto_mem_in_ar_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_1_auto_out_r_valid = plfg_auto_mem_in_r_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_1_auto_out_r_bits_id = 1'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_1_auto_out_r_bits_data = plfg_auto_mem_in_r_bits_data; // @[LazyModule.scala 167:31]
  assign axi4buf_1_auto_out_r_bits_resp = plfg_auto_mem_in_r_bits_resp; // @[LazyModule.scala 167:31]
  assign axi4buf_1_auto_out_r_bits_last = plfg_auto_mem_in_r_bits_last; // @[LazyModule.scala 167:31]
  assign axi4buf_2_clock = clock;
  assign axi4buf_2_reset = reset;
  assign axi4buf_2_auto_in_aw_valid = bus_auto_out_2_aw_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_2_auto_in_aw_bits_id = bus_auto_out_2_aw_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_2_auto_in_aw_bits_addr = bus_auto_out_2_aw_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_2_auto_in_aw_bits_size = bus_auto_out_2_aw_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_2_auto_in_w_valid = bus_auto_out_2_w_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_2_auto_in_w_bits_data = bus_auto_out_2_w_bits_data; // @[LazyModule.scala 167:57]
  assign axi4buf_2_auto_in_w_bits_strb = bus_auto_out_2_w_bits_strb; // @[LazyModule.scala 167:57]
  assign axi4buf_2_auto_in_w_bits_last = bus_auto_out_2_w_bits_last; // @[LazyModule.scala 167:57]
  assign axi4buf_2_auto_in_b_ready = bus_auto_out_2_b_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_2_auto_in_ar_valid = bus_auto_out_2_ar_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_2_auto_in_ar_bits_id = bus_auto_out_2_ar_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_2_auto_in_ar_bits_addr = bus_auto_out_2_ar_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_2_auto_in_ar_bits_size = bus_auto_out_2_ar_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_2_auto_in_r_ready = bus_auto_out_2_r_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_2_auto_out_aw_ready = plfg_split_auto_mem_in_aw_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_2_auto_out_w_ready = plfg_split_auto_mem_in_w_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_2_auto_out_b_valid = plfg_split_auto_mem_in_b_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_2_auto_out_b_bits_id = plfg_split_auto_mem_in_b_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_2_auto_out_b_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_2_auto_out_ar_ready = plfg_split_auto_mem_in_ar_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_2_auto_out_r_valid = plfg_split_auto_mem_in_r_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_2_auto_out_r_bits_id = plfg_split_auto_mem_in_r_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_2_auto_out_r_bits_data = plfg_split_auto_mem_in_r_bits_data; // @[LazyModule.scala 167:31]
  assign axi4buf_2_auto_out_r_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_2_auto_out_r_bits_last = 1'h1; // @[LazyModule.scala 167:31]
  assign axi4buf_3_clock = clock;
  assign axi4buf_3_reset = reset;
  assign axi4buf_3_auto_in_aw_valid = bus_auto_out_3_aw_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_3_auto_in_aw_bits_id = bus_auto_out_3_aw_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_3_auto_in_aw_bits_addr = bus_auto_out_3_aw_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_3_auto_in_aw_bits_size = bus_auto_out_3_aw_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_3_auto_in_w_valid = bus_auto_out_3_w_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_3_auto_in_w_bits_data = bus_auto_out_3_w_bits_data; // @[LazyModule.scala 167:57]
  assign axi4buf_3_auto_in_w_bits_strb = bus_auto_out_3_w_bits_strb; // @[LazyModule.scala 167:57]
  assign axi4buf_3_auto_in_w_bits_last = bus_auto_out_3_w_bits_last; // @[LazyModule.scala 167:57]
  assign axi4buf_3_auto_in_b_ready = bus_auto_out_3_b_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_3_auto_in_ar_valid = bus_auto_out_3_ar_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_3_auto_in_ar_bits_id = bus_auto_out_3_ar_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_3_auto_in_ar_bits_addr = bus_auto_out_3_ar_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_3_auto_in_ar_bits_size = bus_auto_out_3_ar_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_3_auto_in_r_ready = bus_auto_out_3_r_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_3_auto_out_aw_ready = plfg_mux_0_auto_register_in_aw_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_3_auto_out_w_ready = plfg_mux_0_auto_register_in_w_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_3_auto_out_b_valid = plfg_mux_0_auto_register_in_b_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_3_auto_out_b_bits_id = plfg_mux_0_auto_register_in_b_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_3_auto_out_b_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_3_auto_out_ar_ready = plfg_mux_0_auto_register_in_ar_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_3_auto_out_r_valid = plfg_mux_0_auto_register_in_r_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_3_auto_out_r_bits_id = plfg_mux_0_auto_register_in_r_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_3_auto_out_r_bits_data = plfg_mux_0_auto_register_in_r_bits_data; // @[LazyModule.scala 167:31]
  assign axi4buf_3_auto_out_r_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_3_auto_out_r_bits_last = 1'h1; // @[LazyModule.scala 167:31]
  assign axi4buf_4_clock = clock;
  assign axi4buf_4_reset = reset;
  assign axi4buf_4_auto_in_aw_valid = bus_auto_out_4_aw_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_4_auto_in_aw_bits_id = bus_auto_out_4_aw_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_4_auto_in_aw_bits_addr = bus_auto_out_4_aw_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_4_auto_in_aw_bits_size = bus_auto_out_4_aw_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_4_auto_in_w_valid = bus_auto_out_4_w_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_4_auto_in_w_bits_data = bus_auto_out_4_w_bits_data; // @[LazyModule.scala 167:57]
  assign axi4buf_4_auto_in_w_bits_strb = bus_auto_out_4_w_bits_strb; // @[LazyModule.scala 167:57]
  assign axi4buf_4_auto_in_w_bits_last = bus_auto_out_4_w_bits_last; // @[LazyModule.scala 167:57]
  assign axi4buf_4_auto_in_b_ready = bus_auto_out_4_b_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_4_auto_in_ar_valid = bus_auto_out_4_ar_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_4_auto_in_ar_bits_id = bus_auto_out_4_ar_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_4_auto_in_ar_bits_addr = bus_auto_out_4_ar_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_4_auto_in_ar_bits_size = bus_auto_out_4_ar_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_4_auto_in_r_ready = bus_auto_out_4_r_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_4_auto_out_aw_ready = plfg_mux_1_auto_register_in_aw_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_4_auto_out_w_ready = plfg_mux_1_auto_register_in_w_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_4_auto_out_b_valid = plfg_mux_1_auto_register_in_b_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_4_auto_out_b_bits_id = plfg_mux_1_auto_register_in_b_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_4_auto_out_b_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_4_auto_out_ar_ready = plfg_mux_1_auto_register_in_ar_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_4_auto_out_r_valid = plfg_mux_1_auto_register_in_r_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_4_auto_out_r_bits_id = plfg_mux_1_auto_register_in_r_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_4_auto_out_r_bits_data = plfg_mux_1_auto_register_in_r_bits_data; // @[LazyModule.scala 167:31]
  assign axi4buf_4_auto_out_r_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_4_auto_out_r_bits_last = 1'h1; // @[LazyModule.scala 167:31]
  assign axi4buf_5_clock = clock;
  assign axi4buf_5_reset = reset;
  assign axi4buf_5_auto_in_aw_valid = bus_auto_out_5_aw_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_5_auto_in_aw_bits_id = bus_auto_out_5_aw_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_5_auto_in_aw_bits_addr = bus_auto_out_5_aw_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_5_auto_in_aw_bits_size = bus_auto_out_5_aw_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_5_auto_in_w_valid = bus_auto_out_5_w_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_5_auto_in_w_bits_data = bus_auto_out_5_w_bits_data; // @[LazyModule.scala 167:57]
  assign axi4buf_5_auto_in_w_bits_strb = bus_auto_out_5_w_bits_strb; // @[LazyModule.scala 167:57]
  assign axi4buf_5_auto_in_w_bits_last = bus_auto_out_5_w_bits_last; // @[LazyModule.scala 167:57]
  assign axi4buf_5_auto_in_b_ready = bus_auto_out_5_b_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_5_auto_in_ar_valid = bus_auto_out_5_ar_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_5_auto_in_ar_bits_id = bus_auto_out_5_ar_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_5_auto_in_ar_bits_addr = bus_auto_out_5_ar_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_5_auto_in_ar_bits_size = bus_auto_out_5_ar_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_5_auto_in_r_ready = bus_auto_out_5_r_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_5_auto_out_aw_ready = 1'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_5_auto_out_w_ready = 1'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_5_auto_out_b_valid = 1'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_5_auto_out_b_bits_id = 1'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_5_auto_out_b_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_5_auto_out_ar_ready = 1'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_5_auto_out_r_valid = 1'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_5_auto_out_r_bits_id = 1'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_5_auto_out_r_bits_data = 32'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_5_auto_out_r_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_5_auto_out_r_bits_last = 1'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_6_clock = clock;
  assign axi4buf_6_reset = reset;
  assign axi4buf_6_auto_in_aw_valid = bus_auto_out_6_aw_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_6_auto_in_aw_bits_id = bus_auto_out_6_aw_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_6_auto_in_aw_bits_addr = bus_auto_out_6_aw_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_6_auto_in_aw_bits_size = bus_auto_out_6_aw_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_6_auto_in_w_valid = bus_auto_out_6_w_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_6_auto_in_w_bits_data = bus_auto_out_6_w_bits_data; // @[LazyModule.scala 167:57]
  assign axi4buf_6_auto_in_w_bits_strb = bus_auto_out_6_w_bits_strb; // @[LazyModule.scala 167:57]
  assign axi4buf_6_auto_in_w_bits_last = bus_auto_out_6_w_bits_last; // @[LazyModule.scala 167:57]
  assign axi4buf_6_auto_in_b_ready = bus_auto_out_6_b_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_6_auto_in_ar_valid = bus_auto_out_6_ar_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_6_auto_in_ar_bits_id = bus_auto_out_6_ar_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_6_auto_in_ar_bits_addr = bus_auto_out_6_ar_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_6_auto_in_ar_bits_size = bus_auto_out_6_ar_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_6_auto_in_r_ready = bus_auto_out_6_r_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_6_auto_out_aw_ready = nco_split_auto_mem_in_aw_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_6_auto_out_w_ready = nco_split_auto_mem_in_w_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_6_auto_out_b_valid = nco_split_auto_mem_in_b_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_6_auto_out_b_bits_id = nco_split_auto_mem_in_b_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_6_auto_out_b_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_6_auto_out_ar_ready = nco_split_auto_mem_in_ar_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_6_auto_out_r_valid = nco_split_auto_mem_in_r_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_6_auto_out_r_bits_id = nco_split_auto_mem_in_r_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_6_auto_out_r_bits_data = nco_split_auto_mem_in_r_bits_data; // @[LazyModule.scala 167:31]
  assign axi4buf_6_auto_out_r_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_6_auto_out_r_bits_last = 1'h1; // @[LazyModule.scala 167:31]
  assign axi4buf_7_clock = clock;
  assign axi4buf_7_reset = reset;
  assign axi4buf_7_auto_in_aw_valid = bus_auto_out_7_aw_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_7_auto_in_aw_bits_id = bus_auto_out_7_aw_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_7_auto_in_aw_bits_addr = bus_auto_out_7_aw_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_7_auto_in_aw_bits_size = bus_auto_out_7_aw_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_7_auto_in_w_valid = bus_auto_out_7_w_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_7_auto_in_w_bits_data = bus_auto_out_7_w_bits_data; // @[LazyModule.scala 167:57]
  assign axi4buf_7_auto_in_w_bits_strb = bus_auto_out_7_w_bits_strb; // @[LazyModule.scala 167:57]
  assign axi4buf_7_auto_in_w_bits_last = bus_auto_out_7_w_bits_last; // @[LazyModule.scala 167:57]
  assign axi4buf_7_auto_in_b_ready = bus_auto_out_7_b_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_7_auto_in_ar_valid = bus_auto_out_7_ar_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_7_auto_in_ar_bits_id = bus_auto_out_7_ar_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_7_auto_in_ar_bits_addr = bus_auto_out_7_ar_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_7_auto_in_ar_bits_size = bus_auto_out_7_ar_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_7_auto_in_r_ready = bus_auto_out_7_r_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_7_auto_out_aw_ready = nco_mux_0_auto_register_in_aw_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_7_auto_out_w_ready = nco_mux_0_auto_register_in_w_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_7_auto_out_b_valid = nco_mux_0_auto_register_in_b_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_7_auto_out_b_bits_id = nco_mux_0_auto_register_in_b_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_7_auto_out_b_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_7_auto_out_ar_ready = nco_mux_0_auto_register_in_ar_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_7_auto_out_r_valid = nco_mux_0_auto_register_in_r_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_7_auto_out_r_bits_id = nco_mux_0_auto_register_in_r_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_7_auto_out_r_bits_data = nco_mux_0_auto_register_in_r_bits_data; // @[LazyModule.scala 167:31]
  assign axi4buf_7_auto_out_r_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_7_auto_out_r_bits_last = 1'h1; // @[LazyModule.scala 167:31]
  assign axi4buf_8_clock = clock;
  assign axi4buf_8_reset = reset;
  assign axi4buf_8_auto_in_aw_valid = bus_auto_out_8_aw_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_8_auto_in_aw_bits_id = bus_auto_out_8_aw_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_8_auto_in_aw_bits_addr = bus_auto_out_8_aw_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_8_auto_in_aw_bits_size = bus_auto_out_8_aw_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_8_auto_in_w_valid = bus_auto_out_8_w_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_8_auto_in_w_bits_data = bus_auto_out_8_w_bits_data; // @[LazyModule.scala 167:57]
  assign axi4buf_8_auto_in_w_bits_strb = bus_auto_out_8_w_bits_strb; // @[LazyModule.scala 167:57]
  assign axi4buf_8_auto_in_w_bits_last = bus_auto_out_8_w_bits_last; // @[LazyModule.scala 167:57]
  assign axi4buf_8_auto_in_b_ready = bus_auto_out_8_b_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_8_auto_in_ar_valid = bus_auto_out_8_ar_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_8_auto_in_ar_bits_id = bus_auto_out_8_ar_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_8_auto_in_ar_bits_addr = bus_auto_out_8_ar_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_8_auto_in_ar_bits_size = bus_auto_out_8_ar_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_8_auto_in_r_ready = bus_auto_out_8_r_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_8_auto_out_aw_ready = nco_mux_1_auto_register_in_aw_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_8_auto_out_w_ready = nco_mux_1_auto_register_in_w_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_8_auto_out_b_valid = nco_mux_1_auto_register_in_b_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_8_auto_out_b_bits_id = nco_mux_1_auto_register_in_b_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_8_auto_out_b_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_8_auto_out_ar_ready = nco_mux_1_auto_register_in_ar_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_8_auto_out_r_valid = nco_mux_1_auto_register_in_r_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_8_auto_out_r_bits_id = nco_mux_1_auto_register_in_r_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_8_auto_out_r_bits_data = nco_mux_1_auto_register_in_r_bits_data; // @[LazyModule.scala 167:31]
  assign axi4buf_8_auto_out_r_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_8_auto_out_r_bits_last = 1'h1; // @[LazyModule.scala 167:31]
  assign axi4buf_9_clock = clock;
  assign axi4buf_9_reset = reset;
  assign axi4buf_9_auto_in_aw_valid = bus_auto_out_9_aw_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_9_auto_in_aw_bits_id = bus_auto_out_9_aw_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_9_auto_in_aw_bits_addr = bus_auto_out_9_aw_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_9_auto_in_aw_bits_size = bus_auto_out_9_aw_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_9_auto_in_w_valid = bus_auto_out_9_w_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_9_auto_in_w_bits_data = bus_auto_out_9_w_bits_data; // @[LazyModule.scala 167:57]
  assign axi4buf_9_auto_in_w_bits_strb = bus_auto_out_9_w_bits_strb; // @[LazyModule.scala 167:57]
  assign axi4buf_9_auto_in_w_bits_last = bus_auto_out_9_w_bits_last; // @[LazyModule.scala 167:57]
  assign axi4buf_9_auto_in_b_ready = bus_auto_out_9_b_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_9_auto_in_ar_valid = bus_auto_out_9_ar_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_9_auto_in_ar_bits_id = bus_auto_out_9_ar_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_9_auto_in_ar_bits_addr = bus_auto_out_9_ar_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_9_auto_in_ar_bits_size = bus_auto_out_9_ar_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_9_auto_in_r_ready = bus_auto_out_9_r_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_9_auto_out_aw_ready = fft_auto_mem_in_aw_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_9_auto_out_w_ready = fft_auto_mem_in_w_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_9_auto_out_b_valid = fft_auto_mem_in_b_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_9_auto_out_b_bits_id = fft_auto_mem_in_b_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_9_auto_out_b_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_9_auto_out_ar_ready = fft_auto_mem_in_ar_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_9_auto_out_r_valid = fft_auto_mem_in_r_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_9_auto_out_r_bits_id = fft_auto_mem_in_r_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_9_auto_out_r_bits_data = fft_auto_mem_in_r_bits_data; // @[LazyModule.scala 167:31]
  assign axi4buf_9_auto_out_r_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_9_auto_out_r_bits_last = 1'h1; // @[LazyModule.scala 167:31]
  assign axi4buf_10_clock = clock;
  assign axi4buf_10_reset = reset;
  assign axi4buf_10_auto_in_aw_valid = bus_auto_out_10_aw_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_10_auto_in_aw_bits_id = bus_auto_out_10_aw_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_10_auto_in_aw_bits_addr = bus_auto_out_10_aw_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_10_auto_in_aw_bits_size = bus_auto_out_10_aw_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_10_auto_in_w_valid = bus_auto_out_10_w_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_10_auto_in_w_bits_data = bus_auto_out_10_w_bits_data; // @[LazyModule.scala 167:57]
  assign axi4buf_10_auto_in_w_bits_strb = bus_auto_out_10_w_bits_strb; // @[LazyModule.scala 167:57]
  assign axi4buf_10_auto_in_w_bits_last = bus_auto_out_10_w_bits_last; // @[LazyModule.scala 167:57]
  assign axi4buf_10_auto_in_b_ready = bus_auto_out_10_b_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_10_auto_in_ar_valid = bus_auto_out_10_ar_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_10_auto_in_ar_bits_id = bus_auto_out_10_ar_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_10_auto_in_ar_bits_addr = bus_auto_out_10_ar_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_10_auto_in_ar_bits_size = bus_auto_out_10_ar_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_10_auto_in_r_ready = bus_auto_out_10_r_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_10_auto_out_aw_ready = fft_split_auto_mem_in_aw_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_10_auto_out_w_ready = fft_split_auto_mem_in_w_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_10_auto_out_b_valid = fft_split_auto_mem_in_b_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_10_auto_out_b_bits_id = fft_split_auto_mem_in_b_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_10_auto_out_b_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_10_auto_out_ar_ready = fft_split_auto_mem_in_ar_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_10_auto_out_r_valid = fft_split_auto_mem_in_r_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_10_auto_out_r_bits_id = fft_split_auto_mem_in_r_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_10_auto_out_r_bits_data = fft_split_auto_mem_in_r_bits_data; // @[LazyModule.scala 167:31]
  assign axi4buf_10_auto_out_r_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_10_auto_out_r_bits_last = 1'h1; // @[LazyModule.scala 167:31]
  assign axi4buf_11_clock = clock;
  assign axi4buf_11_reset = reset;
  assign axi4buf_11_auto_in_aw_valid = bus_auto_out_11_aw_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_11_auto_in_aw_bits_id = bus_auto_out_11_aw_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_11_auto_in_aw_bits_addr = bus_auto_out_11_aw_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_11_auto_in_aw_bits_size = bus_auto_out_11_aw_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_11_auto_in_w_valid = bus_auto_out_11_w_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_11_auto_in_w_bits_data = bus_auto_out_11_w_bits_data; // @[LazyModule.scala 167:57]
  assign axi4buf_11_auto_in_w_bits_strb = bus_auto_out_11_w_bits_strb; // @[LazyModule.scala 167:57]
  assign axi4buf_11_auto_in_w_bits_last = bus_auto_out_11_w_bits_last; // @[LazyModule.scala 167:57]
  assign axi4buf_11_auto_in_b_ready = bus_auto_out_11_b_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_11_auto_in_ar_valid = bus_auto_out_11_ar_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_11_auto_in_ar_bits_id = bus_auto_out_11_ar_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_11_auto_in_ar_bits_addr = bus_auto_out_11_ar_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_11_auto_in_ar_bits_size = bus_auto_out_11_ar_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_11_auto_in_r_ready = bus_auto_out_11_r_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_11_auto_out_aw_ready = fft_mux_0_auto_register_in_aw_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_11_auto_out_w_ready = fft_mux_0_auto_register_in_w_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_11_auto_out_b_valid = fft_mux_0_auto_register_in_b_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_11_auto_out_b_bits_id = fft_mux_0_auto_register_in_b_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_11_auto_out_b_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_11_auto_out_ar_ready = fft_mux_0_auto_register_in_ar_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_11_auto_out_r_valid = fft_mux_0_auto_register_in_r_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_11_auto_out_r_bits_id = fft_mux_0_auto_register_in_r_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_11_auto_out_r_bits_data = fft_mux_0_auto_register_in_r_bits_data; // @[LazyModule.scala 167:31]
  assign axi4buf_11_auto_out_r_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_11_auto_out_r_bits_last = 1'h1; // @[LazyModule.scala 167:31]
  assign axi4buf_12_clock = clock;
  assign axi4buf_12_reset = reset;
  assign axi4buf_12_auto_in_aw_valid = bus_auto_out_12_aw_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_12_auto_in_aw_bits_id = bus_auto_out_12_aw_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_12_auto_in_aw_bits_addr = bus_auto_out_12_aw_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_12_auto_in_aw_bits_size = bus_auto_out_12_aw_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_12_auto_in_w_valid = bus_auto_out_12_w_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_12_auto_in_w_bits_data = bus_auto_out_12_w_bits_data; // @[LazyModule.scala 167:57]
  assign axi4buf_12_auto_in_w_bits_strb = bus_auto_out_12_w_bits_strb; // @[LazyModule.scala 167:57]
  assign axi4buf_12_auto_in_w_bits_last = bus_auto_out_12_w_bits_last; // @[LazyModule.scala 167:57]
  assign axi4buf_12_auto_in_b_ready = bus_auto_out_12_b_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_12_auto_in_ar_valid = bus_auto_out_12_ar_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_12_auto_in_ar_bits_id = bus_auto_out_12_ar_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_12_auto_in_ar_bits_addr = bus_auto_out_12_ar_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_12_auto_in_ar_bits_size = bus_auto_out_12_ar_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_12_auto_in_r_ready = bus_auto_out_12_r_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_12_auto_out_aw_ready = fft_mux_1_auto_register_in_aw_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_12_auto_out_w_ready = fft_mux_1_auto_register_in_w_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_12_auto_out_b_valid = fft_mux_1_auto_register_in_b_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_12_auto_out_b_bits_id = fft_mux_1_auto_register_in_b_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_12_auto_out_b_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_12_auto_out_ar_ready = fft_mux_1_auto_register_in_ar_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_12_auto_out_r_valid = fft_mux_1_auto_register_in_r_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_12_auto_out_r_bits_id = fft_mux_1_auto_register_in_r_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_12_auto_out_r_bits_data = fft_mux_1_auto_register_in_r_bits_data; // @[LazyModule.scala 167:31]
  assign axi4buf_12_auto_out_r_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_12_auto_out_r_bits_last = 1'h1; // @[LazyModule.scala 167:31]
  assign axi4buf_13_clock = clock;
  assign axi4buf_13_reset = reset;
  assign axi4buf_13_auto_in_aw_valid = bus_auto_out_13_aw_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_13_auto_in_aw_bits_id = bus_auto_out_13_aw_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_13_auto_in_aw_bits_addr = bus_auto_out_13_aw_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_13_auto_in_aw_bits_size = bus_auto_out_13_aw_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_13_auto_in_w_valid = bus_auto_out_13_w_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_13_auto_in_w_bits_data = bus_auto_out_13_w_bits_data; // @[LazyModule.scala 167:57]
  assign axi4buf_13_auto_in_w_bits_strb = bus_auto_out_13_w_bits_strb; // @[LazyModule.scala 167:57]
  assign axi4buf_13_auto_in_w_bits_last = bus_auto_out_13_w_bits_last; // @[LazyModule.scala 167:57]
  assign axi4buf_13_auto_in_b_ready = bus_auto_out_13_b_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_13_auto_in_ar_valid = bus_auto_out_13_ar_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_13_auto_in_ar_bits_id = bus_auto_out_13_ar_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_13_auto_in_ar_bits_addr = bus_auto_out_13_ar_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_13_auto_in_ar_bits_size = bus_auto_out_13_ar_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_13_auto_in_r_ready = bus_auto_out_13_r_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_13_auto_out_aw_ready = mag_auto_mem_in_aw_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_13_auto_out_w_ready = mag_auto_mem_in_w_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_13_auto_out_b_valid = mag_auto_mem_in_b_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_13_auto_out_b_bits_id = mag_auto_mem_in_b_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_13_auto_out_b_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_13_auto_out_ar_ready = mag_auto_mem_in_ar_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_13_auto_out_r_valid = mag_auto_mem_in_r_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_13_auto_out_r_bits_id = mag_auto_mem_in_r_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_13_auto_out_r_bits_data = mag_auto_mem_in_r_bits_data; // @[LazyModule.scala 167:31]
  assign axi4buf_13_auto_out_r_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_13_auto_out_r_bits_last = 1'h1; // @[LazyModule.scala 167:31]
  assign axi4buf_14_clock = clock;
  assign axi4buf_14_reset = reset;
  assign axi4buf_14_auto_in_aw_valid = bus_auto_out_14_aw_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_14_auto_in_aw_bits_id = bus_auto_out_14_aw_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_14_auto_in_aw_bits_addr = bus_auto_out_14_aw_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_14_auto_in_aw_bits_size = bus_auto_out_14_aw_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_14_auto_in_w_valid = bus_auto_out_14_w_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_14_auto_in_w_bits_data = bus_auto_out_14_w_bits_data; // @[LazyModule.scala 167:57]
  assign axi4buf_14_auto_in_w_bits_strb = bus_auto_out_14_w_bits_strb; // @[LazyModule.scala 167:57]
  assign axi4buf_14_auto_in_w_bits_last = bus_auto_out_14_w_bits_last; // @[LazyModule.scala 167:57]
  assign axi4buf_14_auto_in_b_ready = bus_auto_out_14_b_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_14_auto_in_ar_valid = bus_auto_out_14_ar_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_14_auto_in_ar_bits_id = bus_auto_out_14_ar_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_14_auto_in_ar_bits_addr = bus_auto_out_14_ar_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_14_auto_in_ar_bits_size = bus_auto_out_14_ar_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_14_auto_in_r_ready = bus_auto_out_14_r_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_14_auto_out_aw_ready = mag_split_auto_mem_in_aw_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_14_auto_out_w_ready = mag_split_auto_mem_in_w_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_14_auto_out_b_valid = mag_split_auto_mem_in_b_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_14_auto_out_b_bits_id = mag_split_auto_mem_in_b_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_14_auto_out_b_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_14_auto_out_ar_ready = mag_split_auto_mem_in_ar_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_14_auto_out_r_valid = mag_split_auto_mem_in_r_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_14_auto_out_r_bits_id = mag_split_auto_mem_in_r_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_14_auto_out_r_bits_data = mag_split_auto_mem_in_r_bits_data; // @[LazyModule.scala 167:31]
  assign axi4buf_14_auto_out_r_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_14_auto_out_r_bits_last = 1'h1; // @[LazyModule.scala 167:31]
  assign axi4buf_15_clock = clock;
  assign axi4buf_15_reset = reset;
  assign axi4buf_15_auto_in_aw_valid = bus_auto_out_15_aw_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_15_auto_in_aw_bits_id = bus_auto_out_15_aw_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_15_auto_in_aw_bits_addr = bus_auto_out_15_aw_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_15_auto_in_aw_bits_size = bus_auto_out_15_aw_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_15_auto_in_w_valid = bus_auto_out_15_w_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_15_auto_in_w_bits_data = bus_auto_out_15_w_bits_data; // @[LazyModule.scala 167:57]
  assign axi4buf_15_auto_in_w_bits_strb = bus_auto_out_15_w_bits_strb; // @[LazyModule.scala 167:57]
  assign axi4buf_15_auto_in_w_bits_last = bus_auto_out_15_w_bits_last; // @[LazyModule.scala 167:57]
  assign axi4buf_15_auto_in_b_ready = bus_auto_out_15_b_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_15_auto_in_ar_valid = bus_auto_out_15_ar_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_15_auto_in_ar_bits_id = bus_auto_out_15_ar_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_15_auto_in_ar_bits_addr = bus_auto_out_15_ar_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_15_auto_in_ar_bits_size = bus_auto_out_15_ar_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_15_auto_in_r_ready = bus_auto_out_15_r_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_15_auto_out_aw_ready = mag_mux_0_auto_register_in_aw_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_15_auto_out_w_ready = mag_mux_0_auto_register_in_w_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_15_auto_out_b_valid = mag_mux_0_auto_register_in_b_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_15_auto_out_b_bits_id = mag_mux_0_auto_register_in_b_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_15_auto_out_b_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_15_auto_out_ar_ready = mag_mux_0_auto_register_in_ar_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_15_auto_out_r_valid = mag_mux_0_auto_register_in_r_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_15_auto_out_r_bits_id = mag_mux_0_auto_register_in_r_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_15_auto_out_r_bits_data = mag_mux_0_auto_register_in_r_bits_data; // @[LazyModule.scala 167:31]
  assign axi4buf_15_auto_out_r_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_15_auto_out_r_bits_last = 1'h1; // @[LazyModule.scala 167:31]
  assign axi4buf_16_clock = clock;
  assign axi4buf_16_reset = reset;
  assign axi4buf_16_auto_in_aw_valid = bus_auto_out_16_aw_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_16_auto_in_aw_bits_id = bus_auto_out_16_aw_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_16_auto_in_aw_bits_addr = bus_auto_out_16_aw_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_16_auto_in_aw_bits_size = bus_auto_out_16_aw_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_16_auto_in_w_valid = bus_auto_out_16_w_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_16_auto_in_w_bits_data = bus_auto_out_16_w_bits_data; // @[LazyModule.scala 167:57]
  assign axi4buf_16_auto_in_w_bits_strb = bus_auto_out_16_w_bits_strb; // @[LazyModule.scala 167:57]
  assign axi4buf_16_auto_in_w_bits_last = bus_auto_out_16_w_bits_last; // @[LazyModule.scala 167:57]
  assign axi4buf_16_auto_in_b_ready = bus_auto_out_16_b_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_16_auto_in_ar_valid = bus_auto_out_16_ar_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_16_auto_in_ar_bits_id = bus_auto_out_16_ar_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_16_auto_in_ar_bits_addr = bus_auto_out_16_ar_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_16_auto_in_ar_bits_size = bus_auto_out_16_ar_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_16_auto_in_r_ready = bus_auto_out_16_r_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_16_auto_out_aw_ready = mag_mux_1_auto_register_in_aw_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_16_auto_out_w_ready = mag_mux_1_auto_register_in_w_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_16_auto_out_b_valid = mag_mux_1_auto_register_in_b_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_16_auto_out_b_bits_id = mag_mux_1_auto_register_in_b_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_16_auto_out_b_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_16_auto_out_ar_ready = mag_mux_1_auto_register_in_ar_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_16_auto_out_r_valid = mag_mux_1_auto_register_in_r_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_16_auto_out_r_bits_id = mag_mux_1_auto_register_in_r_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_16_auto_out_r_bits_data = mag_mux_1_auto_register_in_r_bits_data; // @[LazyModule.scala 167:31]
  assign axi4buf_16_auto_out_r_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_16_auto_out_r_bits_last = 1'h1; // @[LazyModule.scala 167:31]
  assign axi4buf_17_clock = clock;
  assign axi4buf_17_reset = reset;
  assign axi4buf_17_auto_in_aw_valid = bus_auto_out_17_aw_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_17_auto_in_aw_bits_id = bus_auto_out_17_aw_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_17_auto_in_aw_bits_addr = bus_auto_out_17_aw_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_17_auto_in_aw_bits_size = bus_auto_out_17_aw_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_17_auto_in_w_valid = bus_auto_out_17_w_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_17_auto_in_w_bits_data = bus_auto_out_17_w_bits_data; // @[LazyModule.scala 167:57]
  assign axi4buf_17_auto_in_w_bits_strb = bus_auto_out_17_w_bits_strb; // @[LazyModule.scala 167:57]
  assign axi4buf_17_auto_in_w_bits_last = bus_auto_out_17_w_bits_last; // @[LazyModule.scala 167:57]
  assign axi4buf_17_auto_in_b_ready = bus_auto_out_17_b_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_17_auto_in_ar_valid = bus_auto_out_17_ar_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_17_auto_in_ar_bits_id = bus_auto_out_17_ar_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_17_auto_in_ar_bits_addr = bus_auto_out_17_ar_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_17_auto_in_ar_bits_size = bus_auto_out_17_ar_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_17_auto_in_r_ready = bus_auto_out_17_r_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_17_auto_out_aw_ready = out_mux_auto_register_in_aw_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_17_auto_out_w_ready = out_mux_auto_register_in_w_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_17_auto_out_b_valid = out_mux_auto_register_in_b_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_17_auto_out_b_bits_id = out_mux_auto_register_in_b_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_17_auto_out_b_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_17_auto_out_ar_ready = out_mux_auto_register_in_ar_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_17_auto_out_r_valid = out_mux_auto_register_in_r_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_17_auto_out_r_bits_id = out_mux_auto_register_in_r_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_17_auto_out_r_bits_data = out_mux_auto_register_in_r_bits_data; // @[LazyModule.scala 167:31]
  assign axi4buf_17_auto_out_r_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_17_auto_out_r_bits_last = 1'h1; // @[LazyModule.scala 167:31]
  assign axi4buf_18_clock = clock;
  assign axi4buf_18_reset = reset;
  assign axi4buf_18_auto_in_aw_valid = bus_auto_out_18_aw_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_18_auto_in_aw_bits_id = bus_auto_out_18_aw_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_18_auto_in_aw_bits_addr = bus_auto_out_18_aw_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_18_auto_in_aw_bits_size = bus_auto_out_18_aw_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_18_auto_in_w_valid = bus_auto_out_18_w_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_18_auto_in_w_bits_data = bus_auto_out_18_w_bits_data; // @[LazyModule.scala 167:57]
  assign axi4buf_18_auto_in_w_bits_strb = bus_auto_out_18_w_bits_strb; // @[LazyModule.scala 167:57]
  assign axi4buf_18_auto_in_w_bits_last = bus_auto_out_18_w_bits_last; // @[LazyModule.scala 167:57]
  assign axi4buf_18_auto_in_b_ready = bus_auto_out_18_b_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_18_auto_in_ar_valid = bus_auto_out_18_ar_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_18_auto_in_ar_bits_id = bus_auto_out_18_ar_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_18_auto_in_ar_bits_addr = bus_auto_out_18_ar_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_18_auto_in_ar_bits_size = bus_auto_out_18_ar_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_18_auto_in_r_ready = bus_auto_out_18_r_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_18_auto_out_aw_ready = out_split_auto_mem_in_aw_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_18_auto_out_w_ready = out_split_auto_mem_in_w_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_18_auto_out_b_valid = out_split_auto_mem_in_b_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_18_auto_out_b_bits_id = out_split_auto_mem_in_b_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_18_auto_out_b_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_18_auto_out_ar_ready = out_split_auto_mem_in_ar_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_18_auto_out_r_valid = out_split_auto_mem_in_r_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_18_auto_out_r_bits_id = out_split_auto_mem_in_r_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_18_auto_out_r_bits_data = out_split_auto_mem_in_r_bits_data; // @[LazyModule.scala 167:31]
  assign axi4buf_18_auto_out_r_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_18_auto_out_r_bits_last = 1'h1; // @[LazyModule.scala 167:31]
  assign axi4buf_19_clock = clock;
  assign axi4buf_19_reset = reset;
  assign axi4buf_19_auto_in_aw_valid = bus_auto_out_19_aw_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_19_auto_in_aw_bits_id = bus_auto_out_19_aw_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_19_auto_in_aw_bits_addr = bus_auto_out_19_aw_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_19_auto_in_aw_bits_size = bus_auto_out_19_aw_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_19_auto_in_w_valid = bus_auto_out_19_w_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_19_auto_in_w_bits_data = bus_auto_out_19_w_bits_data; // @[LazyModule.scala 167:57]
  assign axi4buf_19_auto_in_w_bits_strb = bus_auto_out_19_w_bits_strb; // @[LazyModule.scala 167:57]
  assign axi4buf_19_auto_in_w_bits_last = bus_auto_out_19_w_bits_last; // @[LazyModule.scala 167:57]
  assign axi4buf_19_auto_in_b_ready = bus_auto_out_19_b_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_19_auto_in_ar_valid = bus_auto_out_19_ar_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_19_auto_in_ar_bits_id = bus_auto_out_19_ar_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_19_auto_in_ar_bits_addr = bus_auto_out_19_ar_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_19_auto_in_ar_bits_size = bus_auto_out_19_ar_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_19_auto_in_r_ready = bus_auto_out_19_r_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_19_auto_out_aw_ready = uart_auto_mem_in_aw_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_19_auto_out_w_ready = uart_auto_mem_in_w_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_19_auto_out_b_valid = uart_auto_mem_in_b_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_19_auto_out_b_bits_id = uart_auto_mem_in_b_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_19_auto_out_b_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_19_auto_out_ar_ready = uart_auto_mem_in_ar_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_19_auto_out_r_valid = uart_auto_mem_in_r_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_19_auto_out_r_bits_id = uart_auto_mem_in_r_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_19_auto_out_r_bits_data = uart_auto_mem_in_r_bits_data; // @[LazyModule.scala 167:31]
  assign axi4buf_19_auto_out_r_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_19_auto_out_r_bits_last = 1'h1; // @[LazyModule.scala 167:31]
  assign axi4buf_20_clock = clock;
  assign axi4buf_20_reset = reset;
  assign axi4buf_20_auto_in_aw_valid = bus_auto_out_20_aw_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_20_auto_in_aw_bits_id = bus_auto_out_20_aw_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_20_auto_in_aw_bits_addr = bus_auto_out_20_aw_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_20_auto_in_aw_bits_size = bus_auto_out_20_aw_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_20_auto_in_w_valid = bus_auto_out_20_w_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_20_auto_in_w_bits_data = bus_auto_out_20_w_bits_data; // @[LazyModule.scala 167:57]
  assign axi4buf_20_auto_in_w_bits_strb = bus_auto_out_20_w_bits_strb; // @[LazyModule.scala 167:57]
  assign axi4buf_20_auto_in_w_bits_last = bus_auto_out_20_w_bits_last; // @[LazyModule.scala 167:57]
  assign axi4buf_20_auto_in_b_ready = bus_auto_out_20_b_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_20_auto_in_ar_valid = bus_auto_out_20_ar_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_20_auto_in_ar_bits_id = bus_auto_out_20_ar_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_20_auto_in_ar_bits_addr = bus_auto_out_20_ar_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_20_auto_in_ar_bits_size = bus_auto_out_20_ar_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_20_auto_in_r_ready = bus_auto_out_20_r_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_20_auto_out_aw_ready = uRx_split_auto_mem_in_aw_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_20_auto_out_w_ready = uRx_split_auto_mem_in_w_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_20_auto_out_b_valid = uRx_split_auto_mem_in_b_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_20_auto_out_b_bits_id = uRx_split_auto_mem_in_b_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_20_auto_out_b_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_20_auto_out_ar_ready = uRx_split_auto_mem_in_ar_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_20_auto_out_r_valid = uRx_split_auto_mem_in_r_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_20_auto_out_r_bits_id = uRx_split_auto_mem_in_r_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_20_auto_out_r_bits_data = uRx_split_auto_mem_in_r_bits_data; // @[LazyModule.scala 167:31]
  assign axi4buf_20_auto_out_r_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_20_auto_out_r_bits_last = 1'h1; // @[LazyModule.scala 167:31]
  assign buffer_clock = clock;
  assign buffer_reset = reset;
  assign buffer_auto_in_valid = nco_mux_0_auto_stream_out_0_valid; // @[LazyModule.scala 167:57]
  assign buffer_auto_in_bits_data = nco_mux_0_auto_stream_out_0_bits_data; // @[LazyModule.scala 167:57]
  assign buffer_auto_in_bits_last = nco_mux_0_auto_stream_out_0_bits_last; // @[LazyModule.scala 167:57]
  assign buffer_auto_out_ready = fft_auto_stream_in_ready; // @[LazyModule.scala 167:31]
  assign buffer_1_clock = clock;
  assign buffer_1_reset = reset;
  assign buffer_1_auto_in_valid = fft_mux_0_auto_stream_out_0_valid; // @[LazyModule.scala 167:57]
  assign buffer_1_auto_in_bits_data = fft_mux_0_auto_stream_out_0_bits_data; // @[LazyModule.scala 167:57]
  assign buffer_1_auto_in_bits_last = fft_mux_0_auto_stream_out_0_bits_last; // @[LazyModule.scala 167:57]
  assign buffer_1_auto_out_ready = mag_auto_stream_in_ready; // @[LazyModule.scala 167:31]
  assign buffer_2_clock = clock;
  assign buffer_2_reset = reset;
  assign buffer_2_auto_in_valid = mag_mux_0_auto_stream_out_0_valid; // @[LazyModule.scala 167:57]
  assign buffer_2_auto_in_bits_data = mag_mux_0_auto_stream_out_0_bits_data; // @[LazyModule.scala 167:57]
  assign buffer_2_auto_in_bits_last = mag_mux_0_auto_stream_out_0_bits_last; // @[LazyModule.scala 167:57]
  assign buffer_2_auto_out_ready = acc_auto_accumulator_slave_in_ready; // @[LazyModule.scala 167:31]
  assign buffer_3_clock = clock;
  assign buffer_3_reset = reset;
  assign buffer_3_auto_in_valid = mag_mux_1_auto_stream_out_1_valid; // @[LazyModule.scala 167:57]
  assign buffer_3_auto_in_bits_data = mag_mux_1_auto_stream_out_1_bits_data; // @[LazyModule.scala 167:57]
  assign buffer_3_auto_in_bits_last = mag_mux_1_auto_stream_out_1_bits_last; // @[LazyModule.scala 167:57]
  assign buffer_3_auto_out_ready = out_mux_auto_stream_in_1_ready; // @[LazyModule.scala 167:31]
  assign buffer_4_clock = clock;
  assign buffer_4_reset = reset;
  assign buffer_4_auto_in_valid = fft_mux_1_auto_stream_out_1_valid; // @[LazyModule.scala 167:57]
  assign buffer_4_auto_in_bits_data = fft_mux_1_auto_stream_out_1_bits_data; // @[LazyModule.scala 167:57]
  assign buffer_4_auto_in_bits_last = fft_mux_1_auto_stream_out_1_bits_last; // @[LazyModule.scala 167:57]
  assign buffer_4_auto_out_ready = out_mux_auto_stream_in_2_ready; // @[LazyModule.scala 167:31]
  assign buffer_5_clock = clock;
  assign buffer_5_reset = reset;
  assign buffer_5_auto_in_valid = nco_mux_1_auto_stream_out_1_valid; // @[LazyModule.scala 167:57]
  assign buffer_5_auto_in_bits_data = nco_mux_1_auto_stream_out_1_bits_data; // @[LazyModule.scala 167:57]
  assign buffer_5_auto_in_bits_last = nco_mux_1_auto_stream_out_1_bits_last; // @[LazyModule.scala 167:57]
  assign buffer_5_auto_out_ready = out_mux_auto_stream_in_3_ready; // @[LazyModule.scala 167:31]
  assign buffer_6_clock = clock;
  assign buffer_6_reset = reset;
  assign buffer_6_auto_in_valid = plfg_mux_1_auto_stream_out_1_valid; // @[LazyModule.scala 167:57]
  assign buffer_6_auto_in_bits_data = plfg_mux_1_auto_stream_out_1_bits_data; // @[LazyModule.scala 167:57]
  assign buffer_6_auto_in_bits_last = plfg_mux_1_auto_stream_out_1_bits_last; // @[LazyModule.scala 167:57]
  assign buffer_6_auto_out_ready = out_mux_auto_stream_in_4_ready; // @[LazyModule.scala 167:31]
  assign buffer_7_clock = clock;
  assign buffer_7_reset = reset;
  assign buffer_7_auto_in_valid = in_split_auto_stream_out_4_valid; // @[LazyModule.scala 167:57]
  assign buffer_7_auto_in_bits_data = in_split_auto_stream_out_4_bits_data; // @[LazyModule.scala 167:57]
  assign buffer_7_auto_in_bits_last = in_split_auto_stream_out_4_bits_last; // @[LazyModule.scala 167:57]
  assign buffer_7_auto_out_ready = out_mux_auto_stream_in_5_ready; // @[LazyModule.scala 167:31]
  assign buffer_8_clock = clock;
  assign buffer_8_reset = reset;
  assign buffer_8_auto_in_valid = uRx_split_auto_stream_out_4_valid; // @[LazyModule.scala 167:57]
  assign buffer_8_auto_in_bits_data = uRx_split_auto_stream_out_4_bits_data; // @[LazyModule.scala 167:57]
  assign buffer_8_auto_in_bits_last = uRx_split_auto_stream_out_4_bits_last; // @[LazyModule.scala 167:57]
  assign buffer_8_auto_out_ready = out_mux_auto_stream_in_6_ready; // @[LazyModule.scala 167:31]
  assign buffer_9_clock = clock;
  assign buffer_9_reset = reset;
  assign buffer_9_auto_in_valid = out_mux_auto_stream_out_0_valid; // @[LazyModule.scala 167:57]
  assign buffer_9_auto_in_bits_data = out_mux_auto_stream_out_0_bits_data; // @[LazyModule.scala 167:57]
  assign buffer_9_auto_in_bits_last = out_mux_auto_stream_out_0_bits_last; // @[LazyModule.scala 167:57]
  assign buffer_9_auto_out_ready = out_queue_auto_in_in_ready; // @[LazyModule.scala 167:31]
  assign converter_auto_in_aw_valid = ioMem_0_aw_valid; // @[LazyModule.scala 167:57]
  assign converter_auto_in_aw_bits_id = ioMem_0_aw_bits_id; // @[LazyModule.scala 167:57]
  assign converter_auto_in_aw_bits_addr = ioMem_0_aw_bits_addr; // @[LazyModule.scala 167:57]
  assign converter_auto_in_aw_bits_size = ioMem_0_aw_bits_size; // @[LazyModule.scala 167:57]
  assign converter_auto_in_w_valid = ioMem_0_w_valid; // @[LazyModule.scala 167:57]
  assign converter_auto_in_w_bits_data = ioMem_0_w_bits_data; // @[LazyModule.scala 167:57]
  assign converter_auto_in_w_bits_strb = ioMem_0_w_bits_strb; // @[LazyModule.scala 167:57]
  assign converter_auto_in_w_bits_last = ioMem_0_w_bits_last; // @[LazyModule.scala 167:57]
  assign converter_auto_in_b_ready = ioMem_0_b_ready; // @[LazyModule.scala 167:57]
  assign converter_auto_in_ar_valid = ioMem_0_ar_valid; // @[LazyModule.scala 167:57]
  assign converter_auto_in_ar_bits_id = ioMem_0_ar_bits_id; // @[LazyModule.scala 167:57]
  assign converter_auto_in_ar_bits_addr = ioMem_0_ar_bits_addr; // @[LazyModule.scala 167:57]
  assign converter_auto_in_ar_bits_size = ioMem_0_ar_bits_size; // @[LazyModule.scala 167:57]
  assign converter_auto_in_r_ready = ioMem_0_r_ready; // @[LazyModule.scala 167:57]
  assign converter_auto_out_aw_ready = bus_auto_in_aw_ready; // @[LazyModule.scala 167:31]
  assign converter_auto_out_w_ready = bus_auto_in_w_ready; // @[LazyModule.scala 167:31]
  assign converter_auto_out_b_valid = bus_auto_in_b_valid; // @[LazyModule.scala 167:31]
  assign converter_auto_out_b_bits_resp = bus_auto_in_b_bits_resp; // @[LazyModule.scala 167:31]
  assign converter_auto_out_ar_ready = bus_auto_in_ar_ready; // @[LazyModule.scala 167:31]
  assign converter_auto_out_r_valid = bus_auto_in_r_valid; // @[LazyModule.scala 167:31]
  assign converter_auto_out_r_bits_data = bus_auto_in_r_bits_data; // @[LazyModule.scala 167:31]
  assign converter_auto_out_r_bits_resp = bus_auto_in_r_bits_resp; // @[LazyModule.scala 167:31]
  assign converter_auto_out_r_bits_last = bus_auto_in_r_bits_last; // @[LazyModule.scala 167:31]
  assign converter_1_auto_in_valid = widthAdapter_2_auto_out_valid; // @[LazyModule.scala 167:57]
  assign converter_1_auto_in_bits_data = widthAdapter_2_auto_out_bits_data; // @[LazyModule.scala 167:57]
  assign converter_1_auto_in_bits_last = widthAdapter_2_auto_out_bits_last; // @[LazyModule.scala 167:57]
  assign converter_1_auto_out_ready = outStream_0_ready; // @[LazyModule.scala 167:31]
  assign converter_2_auto_in_valid = inStream_0_valid; // @[LazyModule.scala 167:57]
  assign converter_2_auto_in_bits_data = inStream_0_bits_data; // @[LazyModule.scala 167:57]
  assign converter_2_auto_in_bits_last = inStream_0_bits_last; // @[LazyModule.scala 167:57]
  assign converter_2_auto_out_ready = in_queue_auto_in_in_ready; // @[LazyModule.scala 167:31]
endmodule
