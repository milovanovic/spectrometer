module AXI4StreamWidthAdapater_4_to_1(
  input         clock,
  input         reset,
  output        auto_in_ready,
  input         auto_in_valid,
  input  [7:0]  auto_in_bits_data,
  input         auto_in_bits_last,
  input         auto_out_ready,
  output        auto_out_valid,
  output [31:0] auto_out_bits_data,
  output        auto_out_bits_last
);
  reg [7:0] _T; // @[AXI4StreamWidthAdapter.scala 101:37]
  reg [31:0] _RAND_0;
  reg [7:0] _T_1; // @[AXI4StreamWidthAdapter.scala 101:37]
  reg [31:0] _RAND_1;
  reg [7:0] _T_2; // @[AXI4StreamWidthAdapter.scala 101:37]
  reg [31:0] _RAND_2;
  reg [1:0] _T_3; // @[AXI4StreamWidthAdapter.scala 102:22]
  reg [31:0] _RAND_3;
  wire  _T_4 = auto_in_valid & auto_out_ready; // @[AXI4StreamWidthAdapter.scala 103:14]
  wire  _T_5 = _T_3 == 2'h3; // @[AXI4StreamWidthAdapter.scala 103:38]
  wire [2:0] _T_6 = _T_3 + 2'h1; // @[AXI4StreamWidthAdapter.scala 103:60]
  wire [2:0] _T_7 = _T_5 ? 3'h0 : _T_6; // @[AXI4StreamWidthAdapter.scala 103:33]
  wire [2:0] _GEN_0 = _T_4 ? _T_7 : {{1'd0}, _T_3}; // @[AXI4StreamWidthAdapter.scala 103:21]
  wire  _T_9 = _T_3 == 2'h0; // @[AXI4StreamWidthAdapter.scala 106:29]
  wire  _T_10 = _T_4 & _T_9; // @[AXI4StreamWidthAdapter.scala 106:22]
  wire  _T_12 = _T_3 == 2'h1; // @[AXI4StreamWidthAdapter.scala 106:29]
  wire  _T_13 = _T_4 & _T_12; // @[AXI4StreamWidthAdapter.scala 106:22]
  wire  _T_15 = _T_3 == 2'h2; // @[AXI4StreamWidthAdapter.scala 106:29]
  wire  _T_16 = _T_4 & _T_15; // @[AXI4StreamWidthAdapter.scala 106:22]
  wire [23:0] _T_18 = {auto_in_bits_data,_T_2,_T_1}; // @[Cat.scala 29:58]
  wire  ov0 = _T_5 & auto_in_valid; // @[AXI4StreamWidthAdapter.scala 112:32]
  reg  _T_20; // @[AXI4StreamWidthAdapter.scala 101:37]
  reg [31:0] _RAND_4;
  reg  _T_21; // @[AXI4StreamWidthAdapter.scala 101:37]
  reg [31:0] _RAND_5;
  reg  _T_22; // @[AXI4StreamWidthAdapter.scala 101:37]
  reg [31:0] _RAND_6;
  reg [1:0] _T_23; // @[AXI4StreamWidthAdapter.scala 102:22]
  reg [31:0] _RAND_7;
  wire  _T_25 = _T_23 == 2'h3; // @[AXI4StreamWidthAdapter.scala 103:38]
  wire [2:0] _T_26 = _T_23 + 2'h1; // @[AXI4StreamWidthAdapter.scala 103:60]
  wire [2:0] _T_27 = _T_25 ? 3'h0 : _T_26; // @[AXI4StreamWidthAdapter.scala 103:33]
  wire [2:0] _GEN_4 = _T_4 ? _T_27 : {{1'd0}, _T_23}; // @[AXI4StreamWidthAdapter.scala 103:21]
  wire  _T_29 = _T_23 == 2'h0; // @[AXI4StreamWidthAdapter.scala 106:29]
  wire  _T_30 = _T_4 & _T_29; // @[AXI4StreamWidthAdapter.scala 106:22]
  wire  _T_32 = _T_23 == 2'h1; // @[AXI4StreamWidthAdapter.scala 106:29]
  wire  _T_33 = _T_4 & _T_32; // @[AXI4StreamWidthAdapter.scala 106:22]
  wire  _T_35 = _T_23 == 2'h2; // @[AXI4StreamWidthAdapter.scala 106:29]
  wire  _T_36 = _T_4 & _T_35; // @[AXI4StreamWidthAdapter.scala 106:22]
  wire [3:0] _T_39 = {auto_in_bits_last,_T_22,_T_21,_T_20}; // @[Cat.scala 29:58]
  wire  ov1 = _T_25 & auto_in_valid; // @[AXI4StreamWidthAdapter.scala 112:32]
  reg [1:0] _T_44; // @[AXI4StreamWidthAdapter.scala 102:22]
  reg [31:0] _RAND_8;
  wire  _T_46 = _T_44 == 2'h3; // @[AXI4StreamWidthAdapter.scala 103:38]
  wire [2:0] _T_47 = _T_44 + 2'h1; // @[AXI4StreamWidthAdapter.scala 103:60]
  wire [2:0] _T_48 = _T_46 ? 3'h0 : _T_47; // @[AXI4StreamWidthAdapter.scala 103:33]
  wire [2:0] _GEN_8 = _T_4 ? _T_48 : {{1'd0}, _T_44}; // @[AXI4StreamWidthAdapter.scala 103:21]
  wire  ov2 = _T_46 & auto_in_valid; // @[AXI4StreamWidthAdapter.scala 112:32]
  reg [1:0] _T_64; // @[AXI4StreamWidthAdapter.scala 102:22]
  reg [31:0] _RAND_9;
  wire  _T_66 = _T_64 == 2'h3; // @[AXI4StreamWidthAdapter.scala 103:38]
  wire [2:0] _T_67 = _T_64 + 2'h1; // @[AXI4StreamWidthAdapter.scala 103:60]
  wire [2:0] _T_68 = _T_66 ? 3'h0 : _T_67; // @[AXI4StreamWidthAdapter.scala 103:33]
  wire [2:0] _GEN_12 = _T_4 ? _T_68 : {{1'd0}, _T_64}; // @[AXI4StreamWidthAdapter.scala 103:21]
  wire  ov3 = _T_66 & auto_in_valid; // @[AXI4StreamWidthAdapter.scala 112:32]
  reg [1:0] _T_84; // @[AXI4StreamWidthAdapter.scala 102:22]
  reg [31:0] _RAND_10;
  wire  _T_86 = _T_84 == 2'h3; // @[AXI4StreamWidthAdapter.scala 103:38]
  wire [2:0] _T_87 = _T_84 + 2'h1; // @[AXI4StreamWidthAdapter.scala 103:60]
  wire [2:0] _T_88 = _T_86 ? 3'h0 : _T_87; // @[AXI4StreamWidthAdapter.scala 103:33]
  wire [2:0] _GEN_16 = _T_4 ? _T_88 : {{1'd0}, _T_84}; // @[AXI4StreamWidthAdapter.scala 103:21]
  wire  ov4 = _T_86 & auto_in_valid; // @[AXI4StreamWidthAdapter.scala 112:32]
  wire  _T_101 = ov0 == ov1; // @[AXI4StreamWidthAdapter.scala 42:16]
  wire  _T_103 = _T_101 | reset; // @[AXI4StreamWidthAdapter.scala 42:11]
  wire  _T_104 = ~_T_103; // @[AXI4StreamWidthAdapter.scala 42:11]
  wire  _T_105 = ov0 == ov2; // @[AXI4StreamWidthAdapter.scala 43:16]
  wire  _T_107 = _T_105 | reset; // @[AXI4StreamWidthAdapter.scala 43:11]
  wire  _T_108 = ~_T_107; // @[AXI4StreamWidthAdapter.scala 43:11]
  wire  _T_109 = ov0 == ov3; // @[AXI4StreamWidthAdapter.scala 44:16]
  wire  _T_111 = _T_109 | reset; // @[AXI4StreamWidthAdapter.scala 44:11]
  wire  _T_112 = ~_T_111; // @[AXI4StreamWidthAdapter.scala 44:11]
  wire  _T_113 = ov0 == ov4; // @[AXI4StreamWidthAdapter.scala 45:16]
  wire  _T_115 = _T_113 | reset; // @[AXI4StreamWidthAdapter.scala 45:11]
  wire  _T_116 = ~_T_115; // @[AXI4StreamWidthAdapter.scala 45:11]
  assign auto_in_ready = auto_out_ready; // @[LazyModule.scala 173:31]
  assign auto_out_valid = _T_5 & auto_in_valid; // @[LazyModule.scala 173:49]
  assign auto_out_bits_data = {_T_18,_T}; // @[LazyModule.scala 173:49]
  assign auto_out_bits_last = _T_39 != 4'h0; // @[LazyModule.scala 173:49]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T = _RAND_0[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1 = _RAND_1[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_2 = _RAND_2[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_3 = _RAND_3[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_20 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_21 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_22 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_23 = _RAND_7[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_44 = _RAND_8[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_64 = _RAND_9[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_84 = _RAND_10[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (_T_10) begin
      _T <= auto_in_bits_data;
    end
    if (_T_13) begin
      _T_1 <= auto_in_bits_data;
    end
    if (_T_16) begin
      _T_2 <= auto_in_bits_data;
    end
    if (reset) begin
      _T_3 <= 2'h0;
    end else begin
      _T_3 <= _GEN_0[1:0];
    end
    if (_T_30) begin
      _T_20 <= auto_in_bits_last;
    end
    if (_T_33) begin
      _T_21 <= auto_in_bits_last;
    end
    if (_T_36) begin
      _T_22 <= auto_in_bits_last;
    end
    if (reset) begin
      _T_23 <= 2'h0;
    end else begin
      _T_23 <= _GEN_4[1:0];
    end
    if (reset) begin
      _T_44 <= 2'h0;
    end else begin
      _T_44 <= _GEN_8[1:0];
    end
    if (reset) begin
      _T_64 <= 2'h0;
    end else begin
      _T_64 <= _GEN_12[1:0];
    end
    if (reset) begin
      _T_84 <= 2'h0;
    end else begin
      _T_84 <= _GEN_16[1:0];
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_104) begin
          $fwrite(32'h80000002,"Assertion failed\n    at AXI4StreamWidthAdapter.scala:42 assert(ov0 === ov1)\n"); // @[AXI4StreamWidthAdapter.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_104) begin
          $fatal; // @[AXI4StreamWidthAdapter.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_108) begin
          $fwrite(32'h80000002,"Assertion failed\n    at AXI4StreamWidthAdapter.scala:43 assert(ov0 === ov2)\n"); // @[AXI4StreamWidthAdapter.scala 43:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_108) begin
          $fatal; // @[AXI4StreamWidthAdapter.scala 43:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_112) begin
          $fwrite(32'h80000002,"Assertion failed\n    at AXI4StreamWidthAdapter.scala:44 assert(ov0 === ov3)\n"); // @[AXI4StreamWidthAdapter.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_112) begin
          $fatal; // @[AXI4StreamWidthAdapter.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_116) begin
          $fwrite(32'h80000002,"Assertion failed\n    at AXI4StreamWidthAdapter.scala:45 assert(ov0 === ov4)\n"); // @[AXI4StreamWidthAdapter.scala 45:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_116) begin
          $fatal; // @[AXI4StreamWidthAdapter.scala 45:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module Queue(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input         io_enq_bits_read,
  input  [31:0] io_enq_bits_data,
  input         io_enq_bits_extra,
  input         io_deq_ready,
  output        io_deq_valid,
  output        io_deq_bits_read,
  output [31:0] io_deq_bits_data,
  output        io_deq_bits_extra
);
  reg  _T_read [0:1]; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_0;
  wire  _T_read__T_18_data; // @[Decoupled.scala 218:24]
  wire  _T_read__T_18_addr; // @[Decoupled.scala 218:24]
  wire  _T_read__T_10_data; // @[Decoupled.scala 218:24]
  wire  _T_read__T_10_addr; // @[Decoupled.scala 218:24]
  wire  _T_read__T_10_mask; // @[Decoupled.scala 218:24]
  wire  _T_read__T_10_en; // @[Decoupled.scala 218:24]
  reg [31:0] _T_data [0:1]; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_1;
  wire [31:0] _T_data__T_18_data; // @[Decoupled.scala 218:24]
  wire  _T_data__T_18_addr; // @[Decoupled.scala 218:24]
  wire [31:0] _T_data__T_10_data; // @[Decoupled.scala 218:24]
  wire  _T_data__T_10_addr; // @[Decoupled.scala 218:24]
  wire  _T_data__T_10_mask; // @[Decoupled.scala 218:24]
  wire  _T_data__T_10_en; // @[Decoupled.scala 218:24]
  reg  _T_extra [0:1]; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_2;
  wire  _T_extra__T_18_data; // @[Decoupled.scala 218:24]
  wire  _T_extra__T_18_addr; // @[Decoupled.scala 218:24]
  wire  _T_extra__T_10_data; // @[Decoupled.scala 218:24]
  wire  _T_extra__T_10_addr; // @[Decoupled.scala 218:24]
  wire  _T_extra__T_10_mask; // @[Decoupled.scala 218:24]
  wire  _T_extra__T_10_en; // @[Decoupled.scala 218:24]
  reg  value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_3;
  reg  value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_4;
  reg  _T_1; // @[Decoupled.scala 221:35]
  reg [31:0] _RAND_5;
  wire  _T_2 = value == value_1; // @[Decoupled.scala 223:41]
  wire  _T_3 = ~_T_1; // @[Decoupled.scala 224:36]
  wire  _T_4 = _T_2 & _T_3; // @[Decoupled.scala 224:33]
  wire  _T_5 = _T_2 & _T_1; // @[Decoupled.scala 225:32]
  wire  _T_6 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  _T_8 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire  _T_12 = value + 1'h1; // @[Counter.scala 39:22]
  wire  _T_14 = value_1 + 1'h1; // @[Counter.scala 39:22]
  wire  _T_15 = _T_6 != _T_8; // @[Decoupled.scala 236:16]
  assign _T_read__T_18_addr = value_1;
  assign _T_read__T_18_data = _T_read[_T_read__T_18_addr]; // @[Decoupled.scala 218:24]
  assign _T_read__T_10_data = io_enq_bits_read;
  assign _T_read__T_10_addr = value;
  assign _T_read__T_10_mask = 1'h1;
  assign _T_read__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_data__T_18_addr = value_1;
  assign _T_data__T_18_data = _T_data[_T_data__T_18_addr]; // @[Decoupled.scala 218:24]
  assign _T_data__T_10_data = io_enq_bits_data;
  assign _T_data__T_10_addr = value;
  assign _T_data__T_10_mask = 1'h1;
  assign _T_data__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_extra__T_18_addr = value_1;
  assign _T_extra__T_18_data = _T_extra[_T_extra__T_18_addr]; // @[Decoupled.scala 218:24]
  assign _T_extra__T_10_data = io_enq_bits_extra;
  assign _T_extra__T_10_addr = value;
  assign _T_extra__T_10_mask = 1'h1;
  assign _T_extra__T_10_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~_T_5; // @[Decoupled.scala 241:16]
  assign io_deq_valid = ~_T_4; // @[Decoupled.scala 240:16]
  assign io_deq_bits_read = _T_read__T_18_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_data = _T_data__T_18_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_extra = _T_extra__T_18_data; // @[Decoupled.scala 242:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_read[initvar] = _RAND_0[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_data[initvar] = _RAND_1[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_extra[initvar] = _RAND_2[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  value = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  value_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_1 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T_read__T_10_en & _T_read__T_10_mask) begin
      _T_read[_T_read__T_10_addr] <= _T_read__T_10_data; // @[Decoupled.scala 218:24]
    end
    if(_T_data__T_10_en & _T_data__T_10_mask) begin
      _T_data[_T_data__T_10_addr] <= _T_data__T_10_data; // @[Decoupled.scala 218:24]
    end
    if(_T_extra__T_10_en & _T_extra__T_10_mask) begin
      _T_extra[_T_extra__T_10_addr] <= _T_extra__T_10_data; // @[Decoupled.scala 218:24]
    end
    if (reset) begin
      value <= 1'h0;
    end else if (_T_6) begin
      value <= _T_12;
    end
    if (reset) begin
      value_1 <= 1'h0;
    end else if (_T_8) begin
      value_1 <= _T_14;
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else if (_T_15) begin
      _T_1 <= _T_6;
    end
  end
endmodule
module AXI4Splitter(
  input         clock,
  input         reset,
  output        auto_mem_in_aw_ready,
  input         auto_mem_in_aw_valid,
  input         auto_mem_in_aw_bits_id,
  input  [29:0] auto_mem_in_aw_bits_addr,
  output        auto_mem_in_w_ready,
  input         auto_mem_in_w_valid,
  input  [31:0] auto_mem_in_w_bits_data,
  input  [3:0]  auto_mem_in_w_bits_strb,
  input         auto_mem_in_b_ready,
  output        auto_mem_in_b_valid,
  output        auto_mem_in_b_bits_id,
  output        auto_mem_in_ar_ready,
  input         auto_mem_in_ar_valid,
  input         auto_mem_in_ar_bits_id,
  input  [29:0] auto_mem_in_ar_bits_addr,
  input  [2:0]  auto_mem_in_ar_bits_size,
  input         auto_mem_in_r_ready,
  output        auto_mem_in_r_valid,
  output        auto_mem_in_r_bits_id,
  output [31:0] auto_mem_in_r_bits_data,
  output        auto_stream_in_ready,
  input         auto_stream_in_valid,
  input  [31:0] auto_stream_in_bits_data,
  input         auto_stream_in_bits_last,
  input         auto_stream_out_4_ready,
  output        auto_stream_out_4_valid,
  output [31:0] auto_stream_out_4_bits_data,
  output        auto_stream_out_4_bits_last,
  input         auto_stream_out_3_ready,
  output        auto_stream_out_3_valid,
  output [31:0] auto_stream_out_3_bits_data,
  output        auto_stream_out_3_bits_last,
  input         auto_stream_out_2_ready,
  output        auto_stream_out_2_valid,
  output [31:0] auto_stream_out_2_bits_data,
  output        auto_stream_out_2_bits_last,
  input         auto_stream_out_1_ready,
  output        auto_stream_out_1_valid,
  output [31:0] auto_stream_out_1_bits_data,
  output        auto_stream_out_1_bits_last,
  input         auto_stream_out_0_ready,
  output        auto_stream_out_0_valid,
  output [31:0] auto_stream_out_0_bits_data,
  output        auto_stream_out_0_bits_last
);
  wire  Queue_clock; // @[Decoupled.scala 296:21]
  wire  Queue_reset; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_bits_read; // @[Decoupled.scala 296:21]
  wire [31:0] Queue_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_bits_extra; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_bits_read; // @[Decoupled.scala 296:21]
  wire [31:0] Queue_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_bits_extra; // @[Decoupled.scala 296:21]
  reg [31:0] ctrlReg; // @[Splitter.scala 27:26]
  reg [31:0] _RAND_0;
  reg [31:0] maskReg; // @[Splitter.scala 28:26]
  reg [31:0] _RAND_1;
  wire  _T_7 = auto_mem_in_aw_valid & auto_mem_in_w_valid; // @[RegisterRouter.scala 40:39]
  wire  _T_8 = auto_mem_in_ar_valid | _T_7; // @[RegisterRouter.scala 40:26]
  wire  _T_9 = ~auto_mem_in_ar_valid; // @[RegisterRouter.scala 42:29]
  wire  _T_52_ready = Queue_io_enq_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 299:17]
  wire [29:0] _T_16 = auto_mem_in_ar_valid ? auto_mem_in_ar_bits_addr : auto_mem_in_aw_bits_addr; // @[RegisterRouter.scala 48:19]
  wire [1:0] _T_56 = _T_16[3:2] & 2'h2; // @[RegisterRouter.scala 59:16]
  wire  _T_58 = _T_56 == 2'h0; // @[RegisterRouter.scala 59:16]
  wire  _T_10 = _T_52_ready & _T_9; // @[RegisterRouter.scala 42:26]
  wire [1:0] _T_19 = 2'h1 << auto_mem_in_ar_bits_size[0]; // @[OneHot.scala 65:12]
  wire [1:0] _T_21 = _T_19 | 2'h1; // @[Misc.scala 200:81]
  wire  _T_22 = auto_mem_in_ar_bits_size >= 3'h2; // @[Misc.scala 204:21]
  wire  _T_25 = ~auto_mem_in_ar_bits_addr[1]; // @[Misc.scala 209:20]
  wire  _T_27 = _T_21[1] & _T_25; // @[Misc.scala 213:38]
  wire  _T_28 = _T_22 | _T_27; // @[Misc.scala 213:29]
  wire  _T_30 = _T_21[1] & auto_mem_in_ar_bits_addr[1]; // @[Misc.scala 213:38]
  wire  _T_31 = _T_22 | _T_30; // @[Misc.scala 213:29]
  wire  _T_34 = ~auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 209:20]
  wire  _T_35 = _T_25 & _T_34; // @[Misc.scala 212:27]
  wire  _T_36 = _T_21[0] & _T_35; // @[Misc.scala 213:38]
  wire  _T_37 = _T_28 | _T_36; // @[Misc.scala 213:29]
  wire  _T_38 = _T_25 & auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  wire  _T_39 = _T_21[0] & _T_38; // @[Misc.scala 213:38]
  wire  _T_40 = _T_28 | _T_39; // @[Misc.scala 213:29]
  wire  _T_41 = auto_mem_in_ar_bits_addr[1] & _T_34; // @[Misc.scala 212:27]
  wire  _T_42 = _T_21[0] & _T_41; // @[Misc.scala 213:38]
  wire  _T_43 = _T_31 | _T_42; // @[Misc.scala 213:29]
  wire  _T_44 = auto_mem_in_ar_bits_addr[1] & auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  wire  _T_45 = _T_21[0] & _T_44; // @[Misc.scala 213:38]
  wire  _T_46 = _T_31 | _T_45; // @[Misc.scala 213:29]
  wire [3:0] _T_49 = {_T_46,_T_43,_T_40,_T_37}; // @[Cat.scala 29:58]
  wire [3:0] _T_51 = auto_mem_in_ar_valid ? _T_49 : auto_mem_in_w_bits_strb; // @[RegisterRouter.scala 54:25]
  wire [7:0] _T_70 = _T_51[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_72 = _T_51[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_74 = _T_51[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_76 = _T_51[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_79 = {_T_76,_T_74,_T_72,_T_70}; // @[Cat.scala 29:58]
  wire  _T_98 = _T_79 == 32'hffffffff; // @[RegisterRouter.scala 59:16]
  wire  _T_151 = _T_8 & _T_52_ready; // @[RegisterRouter.scala 59:16]
  wire [1:0] _T_145 = 2'h1 << _T_16[2]; // @[OneHot.scala 58:35]
  wire  _T_168 = _T_151 & _T_9; // @[RegisterRouter.scala 59:16]
  wire  _T_175 = _T_168 & _T_145[1]; // @[RegisterRouter.scala 59:16]
  wire  _T_176 = _T_175 & _T_58; // @[RegisterRouter.scala 59:16]
  wire  _T_105 = _T_176 & _T_98; // @[RegisterRouter.scala 59:16]
  wire  _T_170 = _T_168 & _T_145[0]; // @[RegisterRouter.scala 59:16]
  wire  _T_171 = _T_170 & _T_58; // @[RegisterRouter.scala 59:16]
  wire  _T_128 = _T_171 & _T_98; // @[RegisterRouter.scala 59:16]
  wire  _GEN_11 = _T_16[2] ? _T_58 : _T_58; // @[MuxLiteral.scala 48:10]
  wire [31:0] _GEN_13 = _T_16[2] ? maskReg : ctrlReg; // @[MuxLiteral.scala 48:10]
  wire  _T_226_bits_read = Queue_io_deq_bits_read; // @[Decoupled.scala 317:19 Decoupled.scala 318:14]
  wire  _T_226_valid = Queue_io_deq_valid; // @[Decoupled.scala 317:19 Decoupled.scala 319:15]
  wire  _T_229 = ~_T_226_bits_read; // @[RegisterRouter.scala 65:29]
  wire  _T_232 = auto_stream_out_0_ready | auto_stream_out_1_ready; // @[Splitter.scala 45:34]
  wire  _T_233 = _T_232 | auto_stream_out_2_ready; // @[Splitter.scala 45:34]
  wire  _T_234 = _T_233 | auto_stream_out_3_ready; // @[Splitter.scala 45:34]
  wire  readyOR = _T_234 | auto_stream_out_4_ready; // @[Splitter.scala 45:34]
  wire  _T_235 = auto_stream_out_0_ready & auto_stream_out_1_ready; // @[Splitter.scala 46:34]
  wire  _T_236 = _T_235 & auto_stream_out_2_ready; // @[Splitter.scala 46:34]
  wire  _T_237 = _T_236 & auto_stream_out_3_ready; // @[Splitter.scala 46:34]
  wire  readyAND = _T_237 & auto_stream_out_4_ready; // @[Splitter.scala 46:34]
  wire  _T_238 = ctrlReg == 32'h0; // @[Splitter.scala 49:19]
  wire  _T_239 = ctrlReg == 32'h1; // @[Splitter.scala 52:24]
  wire  _GEN_14 = _T_239 & readyOR; // @[Splitter.scala 52:33]
  wire  _T_242 = ~maskReg[0]; // @[Splitter.scala 62:34]
  wire  _T_246 = ~maskReg[1]; // @[Splitter.scala 62:34]
  wire  _T_250 = ~maskReg[2]; // @[Splitter.scala 62:34]
  wire  _T_254 = ~maskReg[3]; // @[Splitter.scala 62:34]
  wire  _T_258 = ~maskReg[4]; // @[Splitter.scala 62:34]
  Queue Queue ( // @[Decoupled.scala 296:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_read(Queue_io_enq_bits_read),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_extra(Queue_io_enq_bits_extra),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_read(Queue_io_deq_bits_read),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_extra(Queue_io_deq_bits_extra)
  );
  assign auto_mem_in_aw_ready = _T_10 & auto_mem_in_w_valid; // @[LazyModule.scala 173:31]
  assign auto_mem_in_w_ready = _T_10 & auto_mem_in_aw_valid; // @[LazyModule.scala 173:31]
  assign auto_mem_in_b_valid = _T_226_valid & _T_229; // @[LazyModule.scala 173:31]
  assign auto_mem_in_b_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_mem_in_ar_ready = Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_valid = _T_226_valid & _T_226_bits_read; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 173:31]
  assign auto_stream_in_ready = _T_238 ? readyAND : _GEN_14; // @[LazyModule.scala 173:31]
  assign auto_stream_out_4_valid = auto_stream_in_valid & _T_258; // @[LazyModule.scala 173:49]
  assign auto_stream_out_4_bits_data = auto_stream_in_bits_data; // @[LazyModule.scala 173:49]
  assign auto_stream_out_4_bits_last = auto_stream_in_bits_last; // @[LazyModule.scala 173:49]
  assign auto_stream_out_3_valid = auto_stream_in_valid & _T_254; // @[LazyModule.scala 173:49]
  assign auto_stream_out_3_bits_data = auto_stream_in_bits_data; // @[LazyModule.scala 173:49]
  assign auto_stream_out_3_bits_last = auto_stream_in_bits_last; // @[LazyModule.scala 173:49]
  assign auto_stream_out_2_valid = auto_stream_in_valid & _T_250; // @[LazyModule.scala 173:49]
  assign auto_stream_out_2_bits_data = auto_stream_in_bits_data; // @[LazyModule.scala 173:49]
  assign auto_stream_out_2_bits_last = auto_stream_in_bits_last; // @[LazyModule.scala 173:49]
  assign auto_stream_out_1_valid = auto_stream_in_valid & _T_246; // @[LazyModule.scala 173:49]
  assign auto_stream_out_1_bits_data = auto_stream_in_bits_data; // @[LazyModule.scala 173:49]
  assign auto_stream_out_1_bits_last = auto_stream_in_bits_last; // @[LazyModule.scala 173:49]
  assign auto_stream_out_0_valid = auto_stream_in_valid & _T_242; // @[LazyModule.scala 173:49]
  assign auto_stream_out_0_bits_data = auto_stream_in_bits_data; // @[LazyModule.scala 173:49]
  assign auto_stream_out_0_bits_last = auto_stream_in_bits_last; // @[LazyModule.scala 173:49]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_mem_in_ar_valid | _T_7; // @[Decoupled.scala 297:22]
  assign Queue_io_enq_bits_read = auto_mem_in_ar_valid; // @[Decoupled.scala 298:21]
  assign Queue_io_enq_bits_data = _GEN_11 ? _GEN_13 : 32'h0; // @[Decoupled.scala 298:21]
  assign Queue_io_enq_bits_extra = auto_mem_in_ar_valid ? auto_mem_in_ar_bits_id : auto_mem_in_aw_bits_id; // @[Decoupled.scala 298:21]
  assign Queue_io_deq_ready = _T_226_bits_read ? auto_mem_in_r_ready : auto_mem_in_b_ready; // @[Decoupled.scala 320:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ctrlReg = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  maskReg = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      ctrlReg <= 32'h0;
    end else if (_T_128) begin
      ctrlReg <= auto_mem_in_w_bits_data;
    end
    if (reset) begin
      maskReg <= 32'h0;
    end else if (_T_105) begin
      maskReg <= auto_mem_in_w_bits_data;
    end
  end
endmodule
module Queue_1(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input  [7:0] io_enq_bits_data,
  input        io_enq_bits_last,
  input        io_deq_ready,
  output       io_deq_valid,
  output [7:0] io_deq_bits_data,
  output       io_deq_bits_last
);
  reg [7:0] _T_data [0:0]; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_0;
  wire [7:0] _T_data__T_14_data; // @[Decoupled.scala 218:24]
  wire  _T_data__T_14_addr; // @[Decoupled.scala 218:24]
  wire [7:0] _T_data__T_10_data; // @[Decoupled.scala 218:24]
  wire  _T_data__T_10_addr; // @[Decoupled.scala 218:24]
  wire  _T_data__T_10_mask; // @[Decoupled.scala 218:24]
  wire  _T_data__T_10_en; // @[Decoupled.scala 218:24]
  reg  _T_last [0:0]; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_1;
  wire  _T_last__T_14_data; // @[Decoupled.scala 218:24]
  wire  _T_last__T_14_addr; // @[Decoupled.scala 218:24]
  wire  _T_last__T_10_data; // @[Decoupled.scala 218:24]
  wire  _T_last__T_10_addr; // @[Decoupled.scala 218:24]
  wire  _T_last__T_10_mask; // @[Decoupled.scala 218:24]
  wire  _T_last__T_10_en; // @[Decoupled.scala 218:24]
  reg  _T_1; // @[Decoupled.scala 221:35]
  reg [31:0] _RAND_2;
  wire  _T_3 = ~_T_1; // @[Decoupled.scala 224:36]
  wire  _T_6 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  _T_8 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_13 = io_deq_ready ? 1'h0 : _T_6; // @[Decoupled.scala 249:27]
  wire  _GEN_22 = _T_3 ? _GEN_13 : _T_6; // @[Decoupled.scala 246:18]
  wire  _GEN_21 = _T_3 ? 1'h0 : _T_8; // @[Decoupled.scala 246:18]
  wire  _T_11 = _GEN_22 != _GEN_21; // @[Decoupled.scala 236:16]
  wire  _T_12 = ~_T_3; // @[Decoupled.scala 240:19]
  assign _T_data__T_14_addr = 1'h0;
  assign _T_data__T_14_data = _T_data[_T_data__T_14_addr]; // @[Decoupled.scala 218:24]
  assign _T_data__T_10_data = io_enq_bits_data;
  assign _T_data__T_10_addr = 1'h0;
  assign _T_data__T_10_mask = 1'h1;
  assign _T_data__T_10_en = _T_3 ? _GEN_13 : _T_6;
  assign _T_last__T_14_addr = 1'h0;
  assign _T_last__T_14_data = _T_last[_T_last__T_14_addr]; // @[Decoupled.scala 218:24]
  assign _T_last__T_10_data = io_enq_bits_last;
  assign _T_last__T_10_addr = 1'h0;
  assign _T_last__T_10_mask = 1'h1;
  assign _T_last__T_10_en = _T_3 ? _GEN_13 : _T_6;
  assign io_enq_ready = io_deq_ready | _T_3; // @[Decoupled.scala 241:16 Decoupled.scala 254:40]
  assign io_deq_valid = io_enq_valid | _T_12; // @[Decoupled.scala 240:16 Decoupled.scala 245:40]
  assign io_deq_bits_data = _T_3 ? io_enq_bits_data : _T_data__T_14_data; // @[Decoupled.scala 242:15 Decoupled.scala 247:19]
  assign io_deq_bits_last = _T_3 ? io_enq_bits_last : _T_last__T_14_data; // @[Decoupled.scala 242:15 Decoupled.scala 247:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_data[initvar] = _RAND_0[7:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_last[initvar] = _RAND_1[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_1 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T_data__T_10_en & _T_data__T_10_mask) begin
      _T_data[_T_data__T_10_addr] <= _T_data__T_10_data; // @[Decoupled.scala 218:24]
    end
    if(_T_last__T_10_en & _T_last__T_10_mask) begin
      _T_last[_T_last__T_10_addr] <= _T_last__T_10_data; // @[Decoupled.scala 218:24]
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else if (_T_11) begin
      if (_T_3) begin
        if (io_deq_ready) begin
          _T_1 <= 1'h0;
        end else begin
          _T_1 <= _T_6;
        end
      end else begin
        _T_1 <= _T_6;
      end
    end
  end
endmodule
module StreamBuffer(
  input        clock,
  input        reset,
  input        auto_out_out_ready,
  output       auto_out_out_valid,
  output [7:0] auto_out_out_bits_data,
  output       auto_out_out_bits_last,
  output       auto_in_in_ready,
  input        auto_in_in_valid,
  input  [7:0] auto_in_in_bits_data,
  input        auto_in_in_bits_last
);
  wire  Queue_clock; // @[Decoupled.scala 296:21]
  wire  Queue_reset; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [7:0] Queue_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_bits_last; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [7:0] Queue_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_bits_last; // @[Decoupled.scala 296:21]
  Queue_1 Queue ( // @[Decoupled.scala 296:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_last(Queue_io_enq_bits_last),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_last(Queue_io_deq_bits_last)
  );
  assign auto_out_out_valid = Queue_io_deq_valid; // @[LazyModule.scala 173:49]
  assign auto_out_out_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_out_bits_last = Queue_io_deq_bits_last; // @[LazyModule.scala 173:49]
  assign auto_in_in_ready = Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_in_in_valid; // @[Decoupled.scala 297:22]
  assign Queue_io_enq_bits_data = auto_in_in_bits_data; // @[Decoupled.scala 298:21]
  assign Queue_io_enq_bits_last = auto_in_in_bits_last; // @[Decoupled.scala 298:21]
  assign Queue_io_deq_ready = auto_out_out_ready; // @[Decoupled.scala 320:15]
endmodule
module QueueCompatibility(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input  [1:0] io_enq_bits,
  input        io_deq_ready,
  output       io_deq_valid,
  output [1:0] io_deq_bits
);
  reg [1:0] _T [0:1]; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_0;
  wire [1:0] _T__T_18_data; // @[Decoupled.scala 218:24]
  wire  _T__T_18_addr; // @[Decoupled.scala 218:24]
  wire [1:0] _T__T_10_data; // @[Decoupled.scala 218:24]
  wire  _T__T_10_addr; // @[Decoupled.scala 218:24]
  wire  _T__T_10_mask; // @[Decoupled.scala 218:24]
  wire  _T__T_10_en; // @[Decoupled.scala 218:24]
  reg  value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_1;
  reg  value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_2;
  reg  _T_1; // @[Decoupled.scala 221:35]
  reg [31:0] _RAND_3;
  wire  _T_2 = value == value_1; // @[Decoupled.scala 223:41]
  wire  _T_3 = ~_T_1; // @[Decoupled.scala 224:36]
  wire  _T_4 = _T_2 & _T_3; // @[Decoupled.scala 224:33]
  wire  _T_5 = _T_2 & _T_1; // @[Decoupled.scala 225:32]
  wire  _T_6 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  _T_8 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire  _T_12 = value + 1'h1; // @[Counter.scala 39:22]
  wire  _GEN_9 = io_deq_ready ? 1'h0 : _T_6; // @[Decoupled.scala 249:27]
  wire  _GEN_12 = _T_4 ? _GEN_9 : _T_6; // @[Decoupled.scala 246:18]
  wire  _T_14 = value_1 + 1'h1; // @[Counter.scala 39:22]
  wire  _GEN_11 = _T_4 ? 1'h0 : _T_8; // @[Decoupled.scala 246:18]
  wire  _T_15 = _GEN_12 != _GEN_11; // @[Decoupled.scala 236:16]
  wire  _T_16 = ~_T_4; // @[Decoupled.scala 240:19]
  assign _T__T_18_addr = value_1;
  assign _T__T_18_data = _T[_T__T_18_addr]; // @[Decoupled.scala 218:24]
  assign _T__T_10_data = io_enq_bits;
  assign _T__T_10_addr = value;
  assign _T__T_10_mask = 1'h1;
  assign _T__T_10_en = _T_4 ? _GEN_9 : _T_6;
  assign io_enq_ready = ~_T_5; // @[Decoupled.scala 241:16]
  assign io_deq_valid = io_enq_valid | _T_16; // @[Decoupled.scala 240:16 Decoupled.scala 245:40]
  assign io_deq_bits = _T_4 ? io_enq_bits : _T__T_18_data; // @[Decoupled.scala 242:15 Decoupled.scala 247:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T[initvar] = _RAND_0[1:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  value = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  value_1 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_1 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T__T_10_en & _T__T_10_mask) begin
      _T[_T__T_10_addr] <= _T__T_10_data; // @[Decoupled.scala 218:24]
    end
    if (reset) begin
      value <= 1'h0;
    end else if (_GEN_12) begin
      value <= _T_12;
    end
    if (reset) begin
      value_1 <= 1'h0;
    end else if (_GEN_11) begin
      value_1 <= _T_14;
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else if (_T_15) begin
      if (_T_4) begin
        if (io_deq_ready) begin
          _T_1 <= 1'h0;
        end else begin
          _T_1 <= _T_6;
        end
      end else begin
        _T_1 <= _T_6;
      end
    end
  end
endmodule
module AXI4Xbar(
  input         clock,
  input         reset,
  output        auto_in_aw_ready,
  input         auto_in_aw_valid,
  input         auto_in_aw_bits_id,
  input  [29:0] auto_in_aw_bits_addr,
  output        auto_in_w_ready,
  input         auto_in_w_valid,
  input  [31:0] auto_in_w_bits_data,
  input  [3:0]  auto_in_w_bits_strb,
  input         auto_in_w_bits_last,
  input         auto_in_b_ready,
  output        auto_in_b_valid,
  output [1:0]  auto_in_b_bits_resp,
  output        auto_in_ar_ready,
  input         auto_in_ar_valid,
  input         auto_in_ar_bits_id,
  input  [29:0] auto_in_ar_bits_addr,
  input  [2:0]  auto_in_ar_bits_size,
  input         auto_in_r_ready,
  output        auto_in_r_valid,
  output [31:0] auto_in_r_bits_data,
  output [1:0]  auto_in_r_bits_resp,
  output        auto_in_r_bits_last,
  input         auto_out_1_aw_ready,
  output        auto_out_1_aw_valid,
  output        auto_out_1_aw_bits_id,
  output [29:0] auto_out_1_aw_bits_addr,
  input         auto_out_1_w_ready,
  output        auto_out_1_w_valid,
  output [31:0] auto_out_1_w_bits_data,
  output [3:0]  auto_out_1_w_bits_strb,
  output        auto_out_1_b_ready,
  input         auto_out_1_b_valid,
  input         auto_out_1_b_bits_id,
  input         auto_out_1_ar_ready,
  output        auto_out_1_ar_valid,
  output        auto_out_1_ar_bits_id,
  output [29:0] auto_out_1_ar_bits_addr,
  output [2:0]  auto_out_1_ar_bits_size,
  output        auto_out_1_r_ready,
  input         auto_out_1_r_valid,
  input         auto_out_1_r_bits_id,
  input  [31:0] auto_out_1_r_bits_data,
  input         auto_out_0_aw_ready,
  output        auto_out_0_aw_valid,
  output [29:0] auto_out_0_aw_bits_addr,
  input         auto_out_0_w_ready,
  output        auto_out_0_w_valid,
  output [31:0] auto_out_0_w_bits_data,
  output        auto_out_0_b_ready,
  input         auto_out_0_b_valid
);
  wire  awIn_0_clock; // @[Xbar.scala 55:47]
  wire  awIn_0_reset; // @[Xbar.scala 55:47]
  wire  awIn_0_io_enq_ready; // @[Xbar.scala 55:47]
  wire  awIn_0_io_enq_valid; // @[Xbar.scala 55:47]
  wire [1:0] awIn_0_io_enq_bits; // @[Xbar.scala 55:47]
  wire  awIn_0_io_deq_ready; // @[Xbar.scala 55:47]
  wire  awIn_0_io_deq_valid; // @[Xbar.scala 55:47]
  wire [1:0] awIn_0_io_deq_bits; // @[Xbar.scala 55:47]
  wire [30:0] _T_1 = {1'b0,$signed(auto_in_ar_bits_addr)}; // @[Parameters.scala 137:49]
  wire [30:0] _T_3 = $signed(_T_1) & 31'sh2000; // @[Parameters.scala 137:52]
  wire  requestARIO_0_0 = $signed(_T_3) == 31'sh0; // @[Parameters.scala 137:67]
  wire [29:0] _T_5 = auto_in_ar_bits_addr ^ 30'h2000; // @[Parameters.scala 137:31]
  wire [30:0] _T_6 = {1'b0,$signed(_T_5)}; // @[Parameters.scala 137:49]
  wire [30:0] _T_8 = $signed(_T_6) & 31'sh2000; // @[Parameters.scala 137:52]
  wire  requestARIO_0_1 = $signed(_T_8) == 31'sh0; // @[Parameters.scala 137:67]
  wire [30:0] _T_11 = {1'b0,$signed(auto_in_aw_bits_addr)}; // @[Parameters.scala 137:49]
  wire [30:0] _T_13 = $signed(_T_11) & 31'sh2000; // @[Parameters.scala 137:52]
  wire  requestAWIO_0_0 = $signed(_T_13) == 31'sh0; // @[Parameters.scala 137:67]
  wire [29:0] _T_15 = auto_in_aw_bits_addr ^ 30'h2000; // @[Parameters.scala 137:31]
  wire [30:0] _T_16 = {1'b0,$signed(_T_15)}; // @[Parameters.scala 137:49]
  wire [30:0] _T_18 = $signed(_T_16) & 31'sh2000; // @[Parameters.scala 137:52]
  wire  requestAWIO_0_1 = $signed(_T_18) == 31'sh0; // @[Parameters.scala 137:67]
  wire  requestROI_1_0 = ~auto_out_1_r_bits_id; // @[Parameters.scala 47:9]
  wire  requestBOI_1_0 = ~auto_out_1_b_bits_id; // @[Parameters.scala 47:9]
  wire [1:0] _T_20 = {requestAWIO_0_1,requestAWIO_0_0}; // @[Xbar.scala 64:75]
  wire  requestWIO_0_0 = awIn_0_io_deq_bits[0]; // @[Xbar.scala 65:73]
  wire  requestWIO_0_1 = awIn_0_io_deq_bits[1]; // @[Xbar.scala 65:73]
  wire [1:0] _T_27 = {requestARIO_0_1,requestARIO_0_0}; // @[Xbar.scala 93:45]
  wire  in_0_ar_ready = requestARIO_0_1 & auto_out_1_ar_ready; // @[Mux.scala 27:72]
  reg [2:0] _T_36; // @[Xbar.scala 104:34]
  reg [31:0] _RAND_0;
  wire  _T_55 = _T_36 == 3'h0; // @[Xbar.scala 112:22]
  reg  _T_37; // @[Xbar.scala 105:29]
  reg [31:0] _RAND_1;
  wire  _T_54 = _T_37 == _T_27[1]; // @[Xbar.scala 111:75]
  wire  _T_56 = _T_55 | _T_54; // @[Xbar.scala 112:34]
  wire  _T_57 = _T_36 != 3'h7; // @[Xbar.scala 112:80]
  wire  _T_59 = _T_56 & _T_57; // @[Xbar.scala 112:48]
  wire  io_in_0_ar_ready = in_0_ar_ready & _T_59; // @[Xbar.scala 130:45]
  wire  _T_31 = io_in_0_ar_ready & auto_in_ar_valid; // @[Decoupled.scala 40:37]
  reg  _T_222; // @[Xbar.scala 242:23]
  reg [31:0] _RAND_2;
  wire  _T_129 = auto_out_1_r_valid & requestROI_1_0; // @[Xbar.scala 222:40]
  reg  _T_278_1; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_3;
  wire  _T_285 = _T_278_1 & _T_129; // @[Mux.scala 27:72]
  wire  in_0_r_valid = _T_222 ? _T_129 : _T_285; // @[Xbar.scala 278:22]
  wire  _T_33 = auto_in_r_ready & in_0_r_valid; // @[Decoupled.scala 40:37]
  wire [1:0] _T_224 = {_T_129,1'h0}; // @[Cat.scala 29:58]
  reg [1:0] _T_231; // @[Arbiter.scala 20:23]
  reg [31:0] _RAND_4;
  wire [1:0] _T_232 = ~_T_231; // @[Arbiter.scala 21:30]
  wire [1:0] _T_233 = _T_224 & _T_232; // @[Arbiter.scala 21:28]
  wire [3:0] _T_234 = {_T_233,_T_129,1'h0}; // @[Cat.scala 29:58]
  wire [3:0] _GEN_18 = {{1'd0}, _T_234[3:1]}; // @[package.scala 208:43]
  wire [3:0] _T_236 = _T_234 | _GEN_18; // @[package.scala 208:43]
  wire [3:0] _T_239 = {_T_231, 2'h0}; // @[Arbiter.scala 22:66]
  wire [3:0] _GEN_19 = {{1'd0}, _T_236[3:1]}; // @[Arbiter.scala 22:58]
  wire [3:0] _T_240 = _GEN_19 | _T_239; // @[Arbiter.scala 22:58]
  wire [1:0] _T_243 = _T_240[3:2] & _T_240[1:0]; // @[Arbiter.scala 23:39]
  wire [1:0] _T_244 = ~_T_243; // @[Arbiter.scala 23:18]
  wire  _T_257 = _T_244[1] & _T_129; // @[Xbar.scala 250:63]
  wire  _T_279_1 = _T_222 ? _T_257 : _T_278_1; // @[Xbar.scala 262:23]
  wire [35:0] _T_295 = {auto_out_1_r_bits_id,auto_out_1_r_bits_data,3'h1}; // @[Mux.scala 27:72]
  wire [35:0] _T_296 = _T_279_1 ? _T_295 : 36'h0; // @[Mux.scala 27:72]
  wire  in_0_r_bits_last = _T_296[0]; // @[Mux.scala 27:72]
  wire  _T_35 = _T_33 & in_0_r_bits_last; // @[Xbar.scala 120:45]
  wire [2:0] _GEN_20 = {{2'd0}, _T_31}; // @[Xbar.scala 106:30]
  wire [2:0] _T_39 = _T_36 + _GEN_20; // @[Xbar.scala 106:30]
  wire [2:0] _GEN_21 = {{2'd0}, _T_35}; // @[Xbar.scala 106:48]
  wire [2:0] _T_41 = _T_39 - _GEN_21; // @[Xbar.scala 106:48]
  wire  _T_42 = ~_T_35; // @[Xbar.scala 107:23]
  wire  _T_43 = _T_36 != 3'h0; // @[Xbar.scala 107:43]
  wire  _T_44 = _T_42 | _T_43; // @[Xbar.scala 107:34]
  wire  _T_46 = _T_44 | reset; // @[Xbar.scala 107:22]
  wire  _T_47 = ~_T_46; // @[Xbar.scala 107:22]
  wire  _T_48 = ~_T_31; // @[Xbar.scala 108:23]
  wire  _T_50 = _T_48 | _T_57; // @[Xbar.scala 108:34]
  wire  _T_52 = _T_50 | reset; // @[Xbar.scala 108:22]
  wire  _T_53 = ~_T_52; // @[Xbar.scala 108:22]
  wire  _T_115 = requestAWIO_0_0 & auto_out_0_aw_ready; // @[Mux.scala 27:72]
  wire  _T_116 = requestAWIO_0_1 & auto_out_1_aw_ready; // @[Mux.scala 27:72]
  wire  in_0_aw_ready = _T_115 | _T_116; // @[Mux.scala 27:72]
  reg  _T_90; // @[Xbar.scala 137:30]
  reg [31:0] _RAND_5;
  wire  _T_94 = _T_90 | awIn_0_io_enq_ready; // @[Xbar.scala 139:57]
  wire  _T_95 = in_0_aw_ready & _T_94; // @[Xbar.scala 139:45]
  reg [2:0] _T_64; // @[Xbar.scala 104:34]
  reg [31:0] _RAND_6;
  wire  _T_83 = _T_64 == 3'h0; // @[Xbar.scala 112:22]
  reg  _T_65; // @[Xbar.scala 105:29]
  reg [31:0] _RAND_7;
  wire  _T_82 = _T_65 == _T_20[1]; // @[Xbar.scala 111:75]
  wire  _T_84 = _T_83 | _T_82; // @[Xbar.scala 112:34]
  wire  _T_85 = _T_64 != 3'h7; // @[Xbar.scala 112:80]
  wire  _T_87 = _T_84 & _T_85; // @[Xbar.scala 112:48]
  wire  io_in_0_aw_ready = _T_95 & _T_87; // @[Xbar.scala 139:82]
  wire  _T_60 = io_in_0_aw_ready & auto_in_aw_valid; // @[Decoupled.scala 40:37]
  reg  _T_304; // @[Xbar.scala 242:23]
  reg [31:0] _RAND_8;
  wire  _T_133 = auto_out_1_b_valid & requestBOI_1_0; // @[Xbar.scala 222:40]
  wire  _T_305 = auto_out_0_b_valid | _T_133; // @[Xbar.scala 246:36]
  reg  _T_360_0; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_9;
  wire  _T_366 = _T_360_0 & auto_out_0_b_valid; // @[Mux.scala 27:72]
  reg  _T_360_1; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_10;
  wire  _T_367 = _T_360_1 & _T_133; // @[Mux.scala 27:72]
  wire  _T_368 = _T_366 | _T_367; // @[Mux.scala 27:72]
  wire  in_0_b_valid = _T_304 ? _T_305 : _T_368; // @[Xbar.scala 278:22]
  wire  _T_62 = auto_in_b_ready & in_0_b_valid; // @[Decoupled.scala 40:37]
  wire [2:0] _GEN_22 = {{2'd0}, _T_60}; // @[Xbar.scala 106:30]
  wire [2:0] _T_67 = _T_64 + _GEN_22; // @[Xbar.scala 106:30]
  wire [2:0] _GEN_23 = {{2'd0}, _T_62}; // @[Xbar.scala 106:48]
  wire [2:0] _T_69 = _T_67 - _GEN_23; // @[Xbar.scala 106:48]
  wire  _T_70 = ~_T_62; // @[Xbar.scala 107:23]
  wire  _T_71 = _T_64 != 3'h0; // @[Xbar.scala 107:43]
  wire  _T_72 = _T_70 | _T_71; // @[Xbar.scala 107:34]
  wire  _T_74 = _T_72 | reset; // @[Xbar.scala 107:22]
  wire  _T_75 = ~_T_74; // @[Xbar.scala 107:22]
  wire  _T_76 = ~_T_60; // @[Xbar.scala 108:23]
  wire  _T_78 = _T_76 | _T_85; // @[Xbar.scala 108:34]
  wire  _T_80 = _T_78 | reset; // @[Xbar.scala 108:22]
  wire  _T_81 = ~_T_80; // @[Xbar.scala 108:22]
  wire  in_0_ar_valid = auto_in_ar_valid & _T_59; // @[Xbar.scala 129:45]
  wire  _T_92 = auto_in_aw_valid & _T_94; // @[Xbar.scala 138:45]
  wire  in_0_aw_valid = _T_92 & _T_87; // @[Xbar.scala 138:82]
  wire  _T_97 = ~_T_90; // @[Xbar.scala 140:54]
  wire  _T_99 = awIn_0_io_enq_ready & awIn_0_io_enq_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_2 = _T_99 | _T_90; // @[Xbar.scala 141:38]
  wire  _T_100 = in_0_aw_ready & in_0_aw_valid; // @[Decoupled.scala 40:37]
  wire  in_0_w_valid = auto_in_w_valid & awIn_0_io_deq_valid; // @[Xbar.scala 145:43]
  wire  _T_122 = requestWIO_0_0 & auto_out_0_w_ready; // @[Mux.scala 27:72]
  wire  _T_123 = requestWIO_0_1 & auto_out_1_w_ready; // @[Mux.scala 27:72]
  wire  in_0_w_ready = _T_122 | _T_123; // @[Mux.scala 27:72]
  wire  _T_103 = auto_in_w_valid & auto_in_w_bits_last; // @[Xbar.scala 147:50]
  wire  out_0_ar_valid = in_0_ar_valid & requestARIO_0_0; // @[Xbar.scala 222:40]
  wire  out_1_ar_valid = in_0_ar_valid & requestARIO_0_1; // @[Xbar.scala 222:40]
  wire  out_0_aw_valid = in_0_aw_valid & requestAWIO_0_0; // @[Xbar.scala 222:40]
  wire  out_1_aw_valid = in_0_aw_valid & requestAWIO_0_1; // @[Xbar.scala 222:40]
  wire  _T_140 = ~out_0_aw_valid; // @[Xbar.scala 256:60]
  wire  _T_146 = _T_140 | out_0_aw_valid; // @[Xbar.scala 258:23]
  wire  _T_148 = _T_146 | reset; // @[Xbar.scala 258:12]
  wire  _T_149 = ~_T_148; // @[Xbar.scala 258:12]
  wire  _T_161 = ~out_0_ar_valid; // @[Xbar.scala 256:60]
  wire  _T_167 = _T_161 | out_0_ar_valid; // @[Xbar.scala 258:23]
  wire  _T_169 = _T_167 | reset; // @[Xbar.scala 258:12]
  wire  _T_170 = ~_T_169; // @[Xbar.scala 258:12]
  wire  _T_184 = ~out_1_aw_valid; // @[Xbar.scala 256:60]
  wire  _T_190 = _T_184 | out_1_aw_valid; // @[Xbar.scala 258:23]
  wire  _T_192 = _T_190 | reset; // @[Xbar.scala 258:12]
  wire  _T_193 = ~_T_192; // @[Xbar.scala 258:12]
  wire  _T_205 = ~out_1_ar_valid; // @[Xbar.scala 256:60]
  wire  _T_211 = _T_205 | out_1_ar_valid; // @[Xbar.scala 258:23]
  wire  _T_213 = _T_211 | reset; // @[Xbar.scala 258:12]
  wire  _T_214 = ~_T_213; // @[Xbar.scala 258:12]
  wire  _T_245 = _T_224 != 2'h0; // @[Arbiter.scala 24:27]
  wire  _T_246 = _T_222 & _T_245; // @[Arbiter.scala 24:18]
  wire [1:0] _T_247 = _T_244 & _T_224; // @[Arbiter.scala 25:29]
  wire [2:0] _T_248 = {_T_247, 1'h0}; // @[package.scala 199:48]
  wire [1:0] _T_250 = _T_247 | _T_248[1:0]; // @[package.scala 199:43]
  wire  _T_271 = ~_T_129; // @[Xbar.scala 258:13]
  wire  _T_273 = _T_271 | _T_257; // @[Xbar.scala 258:23]
  wire  _T_275 = _T_273 | reset; // @[Xbar.scala 258:12]
  wire  _T_276 = ~_T_275; // @[Xbar.scala 258:12]
  wire  _GEN_13 = _T_129 ? 1'h0 : _T_222; // @[Xbar.scala 266:21]
  wire  _GEN_14 = _T_33 | _GEN_13; // @[Xbar.scala 267:24]
  wire  _T_281_1 = _T_222 ? _T_244[1] : _T_278_1; // @[Xbar.scala 270:24]
  wire [1:0] _T_306 = {_T_133,auto_out_0_b_valid}; // @[Cat.scala 29:58]
  reg [1:0] _T_313; // @[Arbiter.scala 20:23]
  reg [31:0] _RAND_11;
  wire [1:0] _T_314 = ~_T_313; // @[Arbiter.scala 21:30]
  wire [1:0] _T_315 = _T_306 & _T_314; // @[Arbiter.scala 21:28]
  wire [3:0] _T_316 = {_T_315,_T_133,auto_out_0_b_valid}; // @[Cat.scala 29:58]
  wire [3:0] _GEN_24 = {{1'd0}, _T_316[3:1]}; // @[package.scala 208:43]
  wire [3:0] _T_318 = _T_316 | _GEN_24; // @[package.scala 208:43]
  wire [3:0] _T_321 = {_T_313, 2'h0}; // @[Arbiter.scala 22:66]
  wire [3:0] _GEN_25 = {{1'd0}, _T_318[3:1]}; // @[Arbiter.scala 22:58]
  wire [3:0] _T_322 = _GEN_25 | _T_321; // @[Arbiter.scala 22:58]
  wire [1:0] _T_325 = _T_322[3:2] & _T_322[1:0]; // @[Arbiter.scala 23:39]
  wire [1:0] _T_326 = ~_T_325; // @[Arbiter.scala 23:18]
  wire  _T_327 = _T_306 != 2'h0; // @[Arbiter.scala 24:27]
  wire  _T_328 = _T_304 & _T_327; // @[Arbiter.scala 24:18]
  wire [1:0] _T_329 = _T_326 & _T_306; // @[Arbiter.scala 25:29]
  wire [2:0] _T_330 = {_T_329, 1'h0}; // @[package.scala 199:48]
  wire [1:0] _T_332 = _T_329 | _T_330[1:0]; // @[package.scala 199:43]
  wire  _T_338 = _T_326[0] & auto_out_0_b_valid; // @[Xbar.scala 250:63]
  wire  _T_339 = _T_326[1] & _T_133; // @[Xbar.scala 250:63]
  wire  _T_342 = _T_338 | _T_339; // @[Xbar.scala 255:50]
  wire  _T_344 = ~_T_338; // @[Xbar.scala 256:60]
  wire  _T_347 = ~_T_339; // @[Xbar.scala 256:60]
  wire  _T_348 = _T_344 | _T_347; // @[Xbar.scala 256:57]
  wire  _T_351 = _T_348 | reset; // @[Xbar.scala 256:11]
  wire  _T_352 = ~_T_351; // @[Xbar.scala 256:11]
  wire  _T_353 = ~_T_305; // @[Xbar.scala 258:13]
  wire  _T_355 = _T_353 | _T_342; // @[Xbar.scala 258:23]
  wire  _T_357 = _T_355 | reset; // @[Xbar.scala 258:12]
  wire  _T_358 = ~_T_357; // @[Xbar.scala 258:12]
  wire  _T_361_1 = _T_304 ? _T_339 : _T_360_1; // @[Xbar.scala 262:23]
  wire  _GEN_16 = _T_305 ? 1'h0 : _T_304; // @[Xbar.scala 266:21]
  wire  _GEN_17 = _T_62 | _GEN_16; // @[Xbar.scala 267:24]
  wire  _T_363_0 = _T_304 ? _T_326[0] : _T_360_0; // @[Xbar.scala 270:24]
  wire  _T_363_1 = _T_304 ? _T_326[1] : _T_360_1; // @[Xbar.scala 270:24]
  wire [2:0] _T_373 = {auto_out_1_b_bits_id,2'h0}; // @[Mux.scala 27:72]
  wire [2:0] _T_374 = _T_361_1 ? _T_373 : 3'h0; // @[Mux.scala 27:72]
  QueueCompatibility awIn_0 ( // @[Xbar.scala 55:47]
    .clock(awIn_0_clock),
    .reset(awIn_0_reset),
    .io_enq_ready(awIn_0_io_enq_ready),
    .io_enq_valid(awIn_0_io_enq_valid),
    .io_enq_bits(awIn_0_io_enq_bits),
    .io_deq_ready(awIn_0_io_deq_ready),
    .io_deq_valid(awIn_0_io_deq_valid),
    .io_deq_bits(awIn_0_io_deq_bits)
  );
  assign auto_in_aw_ready = _T_95 & _T_87; // @[LazyModule.scala 173:31]
  assign auto_in_w_ready = in_0_w_ready & awIn_0_io_deq_valid; // @[LazyModule.scala 173:31]
  assign auto_in_b_valid = _T_304 ? _T_305 : _T_368; // @[LazyModule.scala 173:31]
  assign auto_in_b_bits_resp = _T_374[1:0]; // @[LazyModule.scala 173:31]
  assign auto_in_ar_ready = in_0_ar_ready & _T_59; // @[LazyModule.scala 173:31]
  assign auto_in_r_valid = _T_222 ? _T_129 : _T_285; // @[LazyModule.scala 173:31]
  assign auto_in_r_bits_data = _T_296[34:3]; // @[LazyModule.scala 173:31]
  assign auto_in_r_bits_resp = _T_296[2:1]; // @[LazyModule.scala 173:31]
  assign auto_in_r_bits_last = _T_296[0]; // @[LazyModule.scala 173:31]
  assign auto_out_1_aw_valid = in_0_aw_valid & requestAWIO_0_1; // @[LazyModule.scala 173:49]
  assign auto_out_1_aw_bits_id = auto_in_aw_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_1_aw_bits_addr = auto_in_aw_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_1_w_valid = in_0_w_valid & requestWIO_0_1; // @[LazyModule.scala 173:49]
  assign auto_out_1_w_bits_data = auto_in_w_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_1_w_bits_strb = auto_in_w_bits_strb; // @[LazyModule.scala 173:49]
  assign auto_out_1_b_ready = auto_in_b_ready & _T_363_1; // @[LazyModule.scala 173:49]
  assign auto_out_1_ar_valid = in_0_ar_valid & requestARIO_0_1; // @[LazyModule.scala 173:49]
  assign auto_out_1_ar_bits_id = auto_in_ar_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_1_ar_bits_addr = auto_in_ar_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_1_ar_bits_size = auto_in_ar_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_1_r_ready = auto_in_r_ready & _T_281_1; // @[LazyModule.scala 173:49]
  assign auto_out_0_aw_valid = in_0_aw_valid & requestAWIO_0_0; // @[LazyModule.scala 173:49]
  assign auto_out_0_aw_bits_addr = auto_in_aw_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_0_w_valid = in_0_w_valid & requestWIO_0_0; // @[LazyModule.scala 173:49]
  assign auto_out_0_w_bits_data = auto_in_w_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_0_b_ready = auto_in_b_ready & _T_363_0; // @[LazyModule.scala 173:49]
  assign awIn_0_clock = clock;
  assign awIn_0_reset = reset;
  assign awIn_0_io_enq_valid = auto_in_aw_valid & _T_97; // @[Xbar.scala 140:30]
  assign awIn_0_io_enq_bits = {requestAWIO_0_1,requestAWIO_0_0}; // @[Xbar.scala 64:57]
  assign awIn_0_io_deq_ready = _T_103 & in_0_w_ready; // @[Xbar.scala 147:30]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_36 = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_37 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_222 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_278_1 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_231 = _RAND_4[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_90 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_64 = _RAND_6[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_65 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_304 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_360_0 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_360_1 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_313 = _RAND_11[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      _T_36 <= 3'h0;
    end else begin
      _T_36 <= _T_41;
    end
    if (_T_31) begin
      _T_37 <= _T_27[1];
    end
    _T_222 <= reset | _GEN_14;
    if (reset) begin
      _T_278_1 <= 1'h0;
    end else if (_T_222) begin
      _T_278_1 <= _T_257;
    end
    if (reset) begin
      _T_231 <= 2'h3;
    end else if (_T_246) begin
      _T_231 <= _T_250;
    end
    if (reset) begin
      _T_90 <= 1'h0;
    end else if (_T_100) begin
      _T_90 <= 1'h0;
    end else begin
      _T_90 <= _GEN_2;
    end
    if (reset) begin
      _T_64 <= 3'h0;
    end else begin
      _T_64 <= _T_69;
    end
    if (_T_60) begin
      _T_65 <= _T_20[1];
    end
    _T_304 <= reset | _GEN_17;
    if (reset) begin
      _T_360_0 <= 1'h0;
    end else if (_T_304) begin
      _T_360_0 <= _T_338;
    end
    if (reset) begin
      _T_360_1 <= 1'h0;
    end else if (_T_304) begin
      _T_360_1 <= _T_339;
    end
    if (reset) begin
      _T_313 <= 2'h3;
    end else if (_T_328) begin
      _T_313 <= _T_332;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_47) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:107 assert (!resp_fire || count =/= UInt(0))\n"); // @[Xbar.scala 107:22]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_47) begin
          $fatal; // @[Xbar.scala 107:22]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_53) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:108 assert (!req_fire  || count =/= UInt(flight))\n"); // @[Xbar.scala 108:22]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_53) begin
          $fatal; // @[Xbar.scala 108:22]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_75) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:107 assert (!resp_fire || count =/= UInt(0))\n"); // @[Xbar.scala 107:22]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_75) begin
          $fatal; // @[Xbar.scala 107:22]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_81) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:108 assert (!req_fire  || count =/= UInt(flight))\n"); // @[Xbar.scala 108:22]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_81) begin
          $fatal; // @[Xbar.scala 108:22]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_149) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_149) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_170) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_170) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_193) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_193) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_214) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_214) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_276) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_276) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_352) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:256 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n"); // @[Xbar.scala 256:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_352) begin
          $fatal; // @[Xbar.scala 256:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_358) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_358) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module PLFGDspBlockMem(
  input         clock,
  input         reset,
  output        auto_mem_in_aw_ready,
  input         auto_mem_in_aw_valid,
  input         auto_mem_in_aw_bits_id,
  input  [29:0] auto_mem_in_aw_bits_addr,
  output        auto_mem_in_w_ready,
  input         auto_mem_in_w_valid,
  input  [31:0] auto_mem_in_w_bits_data,
  input  [3:0]  auto_mem_in_w_bits_strb,
  input         auto_mem_in_w_bits_last,
  input         auto_mem_in_b_ready,
  output        auto_mem_in_b_valid,
  output [1:0]  auto_mem_in_b_bits_resp,
  output        auto_mem_in_ar_ready,
  input         auto_mem_in_ar_valid,
  input         auto_mem_in_ar_bits_id,
  input  [29:0] auto_mem_in_ar_bits_addr,
  input  [2:0]  auto_mem_in_ar_bits_size,
  input         auto_mem_in_r_ready,
  output        auto_mem_in_r_valid,
  output [31:0] auto_mem_in_r_bits_data,
  output [1:0]  auto_mem_in_r_bits_resp,
  output        auto_mem_in_r_bits_last,
  input         auto_stream_out_ready,
  output        auto_stream_out_valid,
  output [31:0] auto_stream_out_bits_data,
  output        auto_stream_out_bits_last
);
  wire  axi4xbar_clock; // @[Xbar.scala 211:30]
  wire  axi4xbar_reset; // @[Xbar.scala 211:30]
  wire  axi4xbar_auto_in_aw_ready; // @[Xbar.scala 211:30]
  wire  axi4xbar_auto_in_aw_valid; // @[Xbar.scala 211:30]
  wire  axi4xbar_auto_in_aw_bits_id; // @[Xbar.scala 211:30]
  wire [29:0] axi4xbar_auto_in_aw_bits_addr; // @[Xbar.scala 211:30]
  wire  axi4xbar_auto_in_w_ready; // @[Xbar.scala 211:30]
  wire  axi4xbar_auto_in_w_valid; // @[Xbar.scala 211:30]
  wire [31:0] axi4xbar_auto_in_w_bits_data; // @[Xbar.scala 211:30]
  wire [3:0] axi4xbar_auto_in_w_bits_strb; // @[Xbar.scala 211:30]
  wire  axi4xbar_auto_in_w_bits_last; // @[Xbar.scala 211:30]
  wire  axi4xbar_auto_in_b_ready; // @[Xbar.scala 211:30]
  wire  axi4xbar_auto_in_b_valid; // @[Xbar.scala 211:30]
  wire [1:0] axi4xbar_auto_in_b_bits_resp; // @[Xbar.scala 211:30]
  wire  axi4xbar_auto_in_ar_ready; // @[Xbar.scala 211:30]
  wire  axi4xbar_auto_in_ar_valid; // @[Xbar.scala 211:30]
  wire  axi4xbar_auto_in_ar_bits_id; // @[Xbar.scala 211:30]
  wire [29:0] axi4xbar_auto_in_ar_bits_addr; // @[Xbar.scala 211:30]
  wire [2:0] axi4xbar_auto_in_ar_bits_size; // @[Xbar.scala 211:30]
  wire  axi4xbar_auto_in_r_ready; // @[Xbar.scala 211:30]
  wire  axi4xbar_auto_in_r_valid; // @[Xbar.scala 211:30]
  wire [31:0] axi4xbar_auto_in_r_bits_data; // @[Xbar.scala 211:30]
  wire [1:0] axi4xbar_auto_in_r_bits_resp; // @[Xbar.scala 211:30]
  wire  axi4xbar_auto_in_r_bits_last; // @[Xbar.scala 211:30]
  wire  axi4xbar_auto_out_1_aw_ready; // @[Xbar.scala 211:30]
  wire  axi4xbar_auto_out_1_aw_valid; // @[Xbar.scala 211:30]
  wire  axi4xbar_auto_out_1_aw_bits_id; // @[Xbar.scala 211:30]
  wire [29:0] axi4xbar_auto_out_1_aw_bits_addr; // @[Xbar.scala 211:30]
  wire  axi4xbar_auto_out_1_w_ready; // @[Xbar.scala 211:30]
  wire  axi4xbar_auto_out_1_w_valid; // @[Xbar.scala 211:30]
  wire [31:0] axi4xbar_auto_out_1_w_bits_data; // @[Xbar.scala 211:30]
  wire [3:0] axi4xbar_auto_out_1_w_bits_strb; // @[Xbar.scala 211:30]
  wire  axi4xbar_auto_out_1_b_ready; // @[Xbar.scala 211:30]
  wire  axi4xbar_auto_out_1_b_valid; // @[Xbar.scala 211:30]
  wire  axi4xbar_auto_out_1_b_bits_id; // @[Xbar.scala 211:30]
  wire  axi4xbar_auto_out_1_ar_ready; // @[Xbar.scala 211:30]
  wire  axi4xbar_auto_out_1_ar_valid; // @[Xbar.scala 211:30]
  wire  axi4xbar_auto_out_1_ar_bits_id; // @[Xbar.scala 211:30]
  wire [29:0] axi4xbar_auto_out_1_ar_bits_addr; // @[Xbar.scala 211:30]
  wire [2:0] axi4xbar_auto_out_1_ar_bits_size; // @[Xbar.scala 211:30]
  wire  axi4xbar_auto_out_1_r_ready; // @[Xbar.scala 211:30]
  wire  axi4xbar_auto_out_1_r_valid; // @[Xbar.scala 211:30]
  wire  axi4xbar_auto_out_1_r_bits_id; // @[Xbar.scala 211:30]
  wire [31:0] axi4xbar_auto_out_1_r_bits_data; // @[Xbar.scala 211:30]
  wire  axi4xbar_auto_out_0_aw_ready; // @[Xbar.scala 211:30]
  wire  axi4xbar_auto_out_0_aw_valid; // @[Xbar.scala 211:30]
  wire [29:0] axi4xbar_auto_out_0_aw_bits_addr; // @[Xbar.scala 211:30]
  wire  axi4xbar_auto_out_0_w_ready; // @[Xbar.scala 211:30]
  wire  axi4xbar_auto_out_0_w_valid; // @[Xbar.scala 211:30]
  wire [31:0] axi4xbar_auto_out_0_w_bits_data; // @[Xbar.scala 211:30]
  wire  axi4xbar_auto_out_0_b_ready; // @[Xbar.scala 211:30]
  wire  axi4xbar_auto_out_0_b_valid; // @[Xbar.scala 211:30]
  reg [25:0] configParamsMem1 [0:15]; // @[PLFGDspBlockMem.scala 110:39]
  reg [31:0] _RAND_0;
  wire [25:0] configParamsMem1__T_64_data; // @[PLFGDspBlockMem.scala 110:39]
  wire [3:0] configParamsMem1__T_64_addr; // @[PLFGDspBlockMem.scala 110:39]
  wire [25:0] configParamsMem1__T_14_data; // @[PLFGDspBlockMem.scala 110:39]
  wire [3:0] configParamsMem1__T_14_addr; // @[PLFGDspBlockMem.scala 110:39]
  wire  configParamsMem1__T_14_mask; // @[PLFGDspBlockMem.scala 110:39]
  wire  configParamsMem1__T_14_en; // @[PLFGDspBlockMem.scala 110:39]
  reg  configParamsMem1__T_64_en_pipe_0;
  reg [31:0] _RAND_1;
  reg [3:0] configParamsMem1__T_64_addr_pipe_0;
  reg [31:0] _RAND_2;
  wire  Queue_clock; // @[Decoupled.scala 296:21]
  wire  Queue_reset; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_bits_read; // @[Decoupled.scala 296:21]
  wire [31:0] Queue_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_bits_extra; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_bits_read; // @[Decoupled.scala 296:21]
  wire [31:0] Queue_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_bits_extra; // @[Decoupled.scala 296:21]
  reg  w_full1; // @[PLFGDspBlockMem.scala 114:26]
  reg [31:0] _RAND_3;
  wire [29:0] ramIn1_aw_bits_addr = axi4xbar_auto_out_0_aw_bits_addr; // @[Nodes.scala 370:76 LazyModule.scala 167:31]
  wire  _T_5 = ~w_full1; // @[PLFGDspBlockMem.scala 119:62]
  wire  ramIn1_b_ready = axi4xbar_auto_out_0_b_ready; // @[Nodes.scala 370:76 LazyModule.scala 167:31]
  wire  _T_6 = ramIn1_b_ready | _T_5; // @[PLFGDspBlockMem.scala 119:59]
  wire  ramIn1_w_valid = axi4xbar_auto_out_0_w_valid; // @[Nodes.scala 370:76 LazyModule.scala 167:31]
  wire  ramIn1_aw_ready = ramIn1_w_valid & _T_6; // @[PLFGDspBlockMem.scala 119:40]
  wire  ramIn1_aw_valid = axi4xbar_auto_out_0_aw_valid; // @[Nodes.scala 370:76 LazyModule.scala 167:31]
  wire  _T_11 = ramIn1_b_ready & w_full1; // @[Decoupled.scala 40:37]
  wire  _GEN_0 = _T_11 ? 1'h0 : w_full1; // @[PLFGDspBlockMem.scala 121:29]
  wire  _T_12 = ramIn1_aw_ready & ramIn1_aw_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_1 = _T_12 | _GEN_0; // @[PLFGDspBlockMem.scala 122:29]
  wire [31:0] ramIn1_w_bits_data = axi4xbar_auto_out_0_w_bits_data; // @[Nodes.scala 370:76 LazyModule.scala 167:31]
  reg  enable; // @[PLFGDspBlockMem.scala 130:25]
  reg [31:0] _RAND_4;
  reg  reset_bit; // @[PLFGDspBlockMem.scala 131:28]
  reg [31:0] _RAND_5;
  reg [1:0] frameNum; // @[PLFGDspBlockMem.scala 132:27]
  reg [31:0] _RAND_6;
  reg [15:0] startingPoint; // @[PLFGDspBlockMem.scala 133:32]
  reg [31:0] _RAND_7;
  reg [7:0] interframeNumOfSamples; // @[PLFGDspBlockMem.scala 134:41]
  reg [31:0] _RAND_8;
  reg [2:0] differentChirpsNum; // @[PLFGDspBlockMem.scala 135:37]
  reg [31:0] _RAND_9;
  reg [15:0] currentVal; // @[PLFGDspBlockMem.scala 138:29]
  reg [31:0] _RAND_10;
  reg [7:0] samplesCounter; // @[PLFGDspBlockMem.scala 139:33]
  reg [31:0] _RAND_11;
  reg [1:0] segmentCounter; // @[PLFGDspBlockMem.scala 140:33]
  reg [31:0] _RAND_12;
  reg [1:0] frameCounter; // @[PLFGDspBlockMem.scala 141:31]
  reg [31:0] _RAND_13;
  reg [5:0] framePauseCounter; // @[PLFGDspBlockMem.scala 142:36]
  reg [31:0] _RAND_14;
  reg  end_; // @[PLFGDspBlockMem.scala 143:22]
  reg [31:0] _RAND_15;
  reg [7:0] samplesCounter2; // @[PLFGDspBlockMem.scala 145:34]
  reg [31:0] _RAND_16;
  reg [1:0] segmentCounter2; // @[PLFGDspBlockMem.scala 146:34]
  reg [31:0] _RAND_17;
  reg [1:0] frameCounter2; // @[PLFGDspBlockMem.scala 147:32]
  reg [31:0] _RAND_18;
  reg  end2; // @[PLFGDspBlockMem.scala 149:23]
  reg [31:0] _RAND_19;
  reg [2:0] repeatedChirpsCounter; // @[PLFGDspBlockMem.scala 151:40]
  reg [31:0] _RAND_20;
  reg [2:0] differentChirpsCounter; // @[PLFGDspBlockMem.scala 152:41]
  reg [31:0] _RAND_21;
  reg [2:0] _T_19; // @[PLFGDspBlockMem.scala 154:49]
  reg [31:0] _RAND_22;
  reg [2:0] repeatedChirpsCounter2; // @[PLFGDspBlockMem.scala 154:41]
  reg [31:0] _RAND_23;
  reg [2:0] _T_20; // @[PLFGDspBlockMem.scala 155:50]
  reg [31:0] _RAND_24;
  reg [2:0] differentChirpsCounter2; // @[PLFGDspBlockMem.scala 155:42]
  reg [31:0] _RAND_25;
  reg [1:0] segmentNums_0; // @[PLFGDspBlockMem.scala 158:30]
  reg [31:0] _RAND_26;
  reg [1:0] segmentNums_1; // @[PLFGDspBlockMem.scala 158:30]
  reg [31:0] _RAND_27;
  reg [1:0] segmentNums_2; // @[PLFGDspBlockMem.scala 158:30]
  reg [31:0] _RAND_28;
  reg [1:0] segmentNums_3; // @[PLFGDspBlockMem.scala 158:30]
  reg [31:0] _RAND_29;
  reg [2:0] repeatedChirpNums_0; // @[PLFGDspBlockMem.scala 159:36]
  reg [31:0] _RAND_30;
  reg [2:0] repeatedChirpNums_1; // @[PLFGDspBlockMem.scala 159:36]
  reg [31:0] _RAND_31;
  reg [2:0] repeatedChirpNums_2; // @[PLFGDspBlockMem.scala 159:36]
  reg [31:0] _RAND_32;
  reg [2:0] repeatedChirpNums_3; // @[PLFGDspBlockMem.scala 159:36]
  reg [31:0] _RAND_33;
  reg [2:0] repeatedChirpNums_4; // @[PLFGDspBlockMem.scala 159:36]
  reg [31:0] _RAND_34;
  reg [2:0] repeatedChirpNums_5; // @[PLFGDspBlockMem.scala 159:36]
  reg [31:0] _RAND_35;
  reg [2:0] repeatedChirpNums_6; // @[PLFGDspBlockMem.scala 159:36]
  reg [31:0] _RAND_36;
  reg [2:0] repeatedChirpNums_7; // @[PLFGDspBlockMem.scala 159:36]
  reg [31:0] _RAND_37;
  reg [1:0] chirpOrdinalNums_0; // @[PLFGDspBlockMem.scala 160:35]
  reg [31:0] _RAND_38;
  reg [1:0] chirpOrdinalNums_1; // @[PLFGDspBlockMem.scala 160:35]
  reg [31:0] _RAND_39;
  reg [1:0] chirpOrdinalNums_2; // @[PLFGDspBlockMem.scala 160:35]
  reg [31:0] _RAND_40;
  reg [1:0] chirpOrdinalNums_3; // @[PLFGDspBlockMem.scala 160:35]
  reg [31:0] _RAND_41;
  reg [1:0] chirpOrdinalNums_4; // @[PLFGDspBlockMem.scala 160:35]
  reg [31:0] _RAND_42;
  reg [1:0] chirpOrdinalNums_5; // @[PLFGDspBlockMem.scala 160:35]
  reg [31:0] _RAND_43;
  reg [1:0] chirpOrdinalNums_6; // @[PLFGDspBlockMem.scala 160:35]
  reg [31:0] _RAND_44;
  reg [1:0] chirpOrdinalNums_7; // @[PLFGDspBlockMem.scala 160:35]
  reg [31:0] _RAND_45;
  wire [25:0] dataFromMem = configParamsMem1__T_64_data; // @[PLFGDspBlockMem.scala 162:27 PLFGDspBlockMem.scala 163:17]
  wire  _T_66 = dataFromMem[23:16] > 8'h1; // @[UIntTypeClass.scala 54:47]
  wire [7:0] _T_70 = dataFromMem[23:16] + 8'h1; // @[UIntTypeClass.scala 18:40]
  wire [7:0] numsOfSamples = _T_66 ? dataFromMem[23:16] : _T_70; // @[PLFGDspBlockMem.scala 172:28]
  wire  slopeSigns = dataFromMem[24]; // @[PLFGDspBlockMem.scala 174:33]
  wire  segmentResets = dataFromMem[25]; // @[PLFGDspBlockMem.scala 175:36]
  wire  _T_2_aw_valid = axi4xbar_auto_out_1_aw_valid; // @[Nodes.scala 370:76 LazyModule.scala 167:31]
  wire  _T_2_w_valid = axi4xbar_auto_out_1_w_valid; // @[Nodes.scala 370:76 LazyModule.scala 167:31]
  wire  _T_72 = _T_2_aw_valid & _T_2_w_valid; // @[RegisterRouter.scala 40:39]
  wire  _T_2_ar_valid = axi4xbar_auto_out_1_ar_valid; // @[Nodes.scala 370:76 LazyModule.scala 167:31]
  wire  _T_73 = _T_2_ar_valid | _T_72; // @[RegisterRouter.scala 40:26]
  wire  _T_74 = ~_T_2_ar_valid; // @[RegisterRouter.scala 42:29]
  wire  _T_117_ready = Queue_io_enq_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 299:17]
  wire [29:0] _T_2_ar_bits_addr = axi4xbar_auto_out_1_ar_bits_addr; // @[Nodes.scala 370:76 LazyModule.scala 167:31]
  wire [29:0] _T_2_aw_bits_addr = axi4xbar_auto_out_1_aw_bits_addr; // @[Nodes.scala 370:76 LazyModule.scala 167:31]
  wire [29:0] _T_81 = _T_2_ar_valid ? _T_2_ar_bits_addr : _T_2_aw_bits_addr; // @[RegisterRouter.scala 48:19]
  wire [4:0] _T_825 = {_T_81[6],_T_81[5],_T_81[4],_T_81[3],_T_81[2]}; // @[Cat.scala 29:58]
  wire [5:0] _T_121 = _T_81[7:2] & 6'h20; // @[RegisterRouter.scala 59:16]
  wire  _T_131 = _T_121 == 6'h0; // @[RegisterRouter.scala 59:16]
  wire  _T_75 = _T_117_ready & _T_74; // @[RegisterRouter.scala 42:26]
  wire  _T_2_ar_bits_id = axi4xbar_auto_out_1_ar_bits_id; // @[Nodes.scala 370:76 LazyModule.scala 167:31]
  wire  _T_2_aw_bits_id = axi4xbar_auto_out_1_aw_bits_id; // @[Nodes.scala 370:76 LazyModule.scala 167:31]
  wire [2:0] _T_2_ar_bits_size = axi4xbar_auto_out_1_ar_bits_size; // @[Nodes.scala 370:76 LazyModule.scala 167:31]
  wire [1:0] _T_84 = 2'h1 << _T_2_ar_bits_size[0]; // @[OneHot.scala 65:12]
  wire [1:0] _T_86 = _T_84 | 2'h1; // @[Misc.scala 200:81]
  wire  _T_87 = _T_2_ar_bits_size >= 3'h2; // @[Misc.scala 204:21]
  wire  _T_90 = ~_T_2_ar_bits_addr[1]; // @[Misc.scala 209:20]
  wire  _T_92 = _T_86[1] & _T_90; // @[Misc.scala 213:38]
  wire  _T_93 = _T_87 | _T_92; // @[Misc.scala 213:29]
  wire  _T_95 = _T_86[1] & _T_2_ar_bits_addr[1]; // @[Misc.scala 213:38]
  wire  _T_96 = _T_87 | _T_95; // @[Misc.scala 213:29]
  wire  _T_99 = ~_T_2_ar_bits_addr[0]; // @[Misc.scala 209:20]
  wire  _T_100 = _T_90 & _T_99; // @[Misc.scala 212:27]
  wire  _T_101 = _T_86[0] & _T_100; // @[Misc.scala 213:38]
  wire  _T_102 = _T_93 | _T_101; // @[Misc.scala 213:29]
  wire  _T_103 = _T_90 & _T_2_ar_bits_addr[0]; // @[Misc.scala 212:27]
  wire  _T_104 = _T_86[0] & _T_103; // @[Misc.scala 213:38]
  wire  _T_105 = _T_93 | _T_104; // @[Misc.scala 213:29]
  wire  _T_106 = _T_2_ar_bits_addr[1] & _T_99; // @[Misc.scala 212:27]
  wire  _T_107 = _T_86[0] & _T_106; // @[Misc.scala 213:38]
  wire  _T_108 = _T_96 | _T_107; // @[Misc.scala 213:29]
  wire  _T_109 = _T_2_ar_bits_addr[1] & _T_2_ar_bits_addr[0]; // @[Misc.scala 212:27]
  wire  _T_110 = _T_86[0] & _T_109; // @[Misc.scala 213:38]
  wire  _T_111 = _T_96 | _T_110; // @[Misc.scala 213:29]
  wire [3:0] _T_114 = {_T_111,_T_108,_T_105,_T_102}; // @[Cat.scala 29:58]
  wire [3:0] _T_2_w_bits_strb = axi4xbar_auto_out_1_w_bits_strb; // @[Nodes.scala 370:76 LazyModule.scala 167:31]
  wire [3:0] _T_116 = _T_2_ar_valid ? _T_114 : _T_2_w_bits_strb; // @[RegisterRouter.scala 54:25]
  wire [7:0] _T_183 = _T_116[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_185 = _T_116[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_187 = _T_116[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_189 = _T_116[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_192 = {_T_189,_T_187,_T_185,_T_183}; // @[Cat.scala 29:58]
  wire  _T_892 = _T_73 & _T_117_ready; // @[RegisterRouter.scala 59:16]
  wire [31:0] _T_826 = 32'h1 << _T_825; // @[OneHot.scala 58:35]
  wire  _T_1059 = _T_892 & _T_74; // @[RegisterRouter.scala 59:16]
  wire  _T_1061 = _T_1059 & _T_826[0]; // @[RegisterRouter.scala 59:16]
  wire  _T_1062 = _T_1061 & _T_131; // @[RegisterRouter.scala 59:16]
  wire  _T_218 = _T_1062 & _T_192[0]; // @[RegisterRouter.scala 59:16]
  wire [31:0] _T_2_w_bits_data = axi4xbar_auto_out_1_w_bits_data; // @[Nodes.scala 370:76 LazyModule.scala 167:31]
  wire  _T_234 = _T_192[15:0] == 16'hffff; // @[RegisterRouter.scala 59:16]
  wire  _T_1086 = _T_1059 & _T_826[5]; // @[RegisterRouter.scala 59:16]
  wire  _T_1087 = _T_1086 & _T_131; // @[RegisterRouter.scala 59:16]
  wire  _T_241 = _T_1087 & _T_234; // @[RegisterRouter.scala 59:16]
  wire  _T_257 = _T_192[2:0] == 3'h7; // @[RegisterRouter.scala 59:16]
  wire  _T_1111 = _T_1059 & _T_826[10]; // @[RegisterRouter.scala 59:16]
  wire  _T_1112 = _T_1111 & _T_131; // @[RegisterRouter.scala 59:16]
  wire  _T_264 = _T_1112 & _T_257; // @[RegisterRouter.scala 59:16]
  wire  _T_280 = _T_192[1:0] == 2'h3; // @[RegisterRouter.scala 59:16]
  wire  _T_1181 = _T_1059 & _T_826[24]; // @[RegisterRouter.scala 59:16]
  wire  _T_1182 = _T_1181 & _T_131; // @[RegisterRouter.scala 59:16]
  wire  _T_287 = _T_1182 & _T_280; // @[RegisterRouter.scala 59:16]
  wire  _T_1186 = _T_1059 & _T_826[25]; // @[RegisterRouter.scala 59:16]
  wire  _T_1187 = _T_1186 & _T_131; // @[RegisterRouter.scala 59:16]
  wire  _T_310 = _T_1187 & _T_280; // @[RegisterRouter.scala 59:16]
  wire  _T_1131 = _T_1059 & _T_826[14]; // @[RegisterRouter.scala 59:16]
  wire  _T_1132 = _T_1131 & _T_131; // @[RegisterRouter.scala 59:16]
  wire  _T_333 = _T_1132 & _T_257; // @[RegisterRouter.scala 59:16]
  wire  _T_1161 = _T_1059 & _T_826[20]; // @[RegisterRouter.scala 59:16]
  wire  _T_1162 = _T_1161 & _T_131; // @[RegisterRouter.scala 59:16]
  wire  _T_356 = _T_1162 & _T_280; // @[RegisterRouter.scala 59:16]
  wire  _T_1066 = _T_1059 & _T_826[1]; // @[RegisterRouter.scala 59:16]
  wire  _T_1067 = _T_1066 & _T_131; // @[RegisterRouter.scala 59:16]
  wire  _T_379 = _T_1067 & _T_192[0]; // @[RegisterRouter.scala 59:16]
  wire  _T_1091 = _T_1059 & _T_826[6]; // @[RegisterRouter.scala 59:16]
  wire  _T_1092 = _T_1091 & _T_131; // @[RegisterRouter.scala 59:16]
  wire  _T_402 = _T_1092 & _T_280; // @[RegisterRouter.scala 59:16]
  wire  _T_1166 = _T_1059 & _T_826[21]; // @[RegisterRouter.scala 59:16]
  wire  _T_1167 = _T_1166 & _T_131; // @[RegisterRouter.scala 59:16]
  wire  _T_425 = _T_1167 & _T_280; // @[RegisterRouter.scala 59:16]
  wire  _T_1106 = _T_1059 & _T_826[9]; // @[RegisterRouter.scala 59:16]
  wire  _T_1107 = _T_1106 & _T_131; // @[RegisterRouter.scala 59:16]
  wire  _T_448 = _T_1107 & _T_280; // @[RegisterRouter.scala 59:16]
  wire  _T_1126 = _T_1059 & _T_826[13]; // @[RegisterRouter.scala 59:16]
  wire  _T_1127 = _T_1126 & _T_131; // @[RegisterRouter.scala 59:16]
  wire  _T_471 = _T_1127 & _T_257; // @[RegisterRouter.scala 59:16]
  wire  _T_1071 = _T_1059 & _T_826[2]; // @[RegisterRouter.scala 59:16]
  wire  _T_1072 = _T_1071 & _T_131; // @[RegisterRouter.scala 59:16]
  wire  _T_494 = _T_1072 & _T_280; // @[RegisterRouter.scala 59:16]
  wire  _T_1146 = _T_1059 & _T_826[17]; // @[RegisterRouter.scala 59:16]
  wire  _T_1147 = _T_1146 & _T_131; // @[RegisterRouter.scala 59:16]
  wire  _T_517 = _T_1147 & _T_257; // @[RegisterRouter.scala 59:16]
  wire  _T_1171 = _T_1059 & _T_826[22]; // @[RegisterRouter.scala 59:16]
  wire  _T_1172 = _T_1171 & _T_131; // @[RegisterRouter.scala 59:16]
  wire  _T_540 = _T_1172 & _T_280; // @[RegisterRouter.scala 59:16]
  wire  _T_1121 = _T_1059 & _T_826[12]; // @[RegisterRouter.scala 59:16]
  wire  _T_1122 = _T_1121 & _T_131; // @[RegisterRouter.scala 59:16]
  wire  _T_563 = _T_1122 & _T_257; // @[RegisterRouter.scala 59:16]
  wire  _T_1096 = _T_1059 & _T_826[7]; // @[RegisterRouter.scala 59:16]
  wire  _T_1097 = _T_1096 & _T_131; // @[RegisterRouter.scala 59:16]
  wire  _T_586 = _T_1097 & _T_280; // @[RegisterRouter.scala 59:16]
  wire  _T_602 = _T_192[9:0] == 10'h3ff; // @[RegisterRouter.scala 59:16]
  wire  _T_1076 = _T_1059 & _T_826[3]; // @[RegisterRouter.scala 59:16]
  wire  _T_1077 = _T_1076 & _T_131; // @[RegisterRouter.scala 59:16]
  wire  _T_609 = _T_1077 & _T_602; // @[RegisterRouter.scala 59:16]
  wire [9:0] _GEN_24 = _T_609 ? _T_2_w_bits_data[9:0] : {{2'd0}, interframeNumOfSamples}; // @[RegField.scala 134:88]
  wire [9:0] _T_620 = {{2'd0}, interframeNumOfSamples}; // @[RegisterRouter.scala 59:16]
  wire  _T_1151 = _T_1059 & _T_826[18]; // @[RegisterRouter.scala 59:16]
  wire  _T_1152 = _T_1151 & _T_131; // @[RegisterRouter.scala 59:16]
  wire  _T_632 = _T_1152 & _T_280; // @[RegisterRouter.scala 59:16]
  wire  _T_1141 = _T_1059 & _T_826[16]; // @[RegisterRouter.scala 59:16]
  wire  _T_1142 = _T_1141 & _T_131; // @[RegisterRouter.scala 59:16]
  wire  _T_655 = _T_1142 & _T_257; // @[RegisterRouter.scala 59:16]
  wire  _T_1116 = _T_1059 & _T_826[11]; // @[RegisterRouter.scala 59:16]
  wire  _T_1117 = _T_1116 & _T_131; // @[RegisterRouter.scala 59:16]
  wire  _T_678 = _T_1117 & _T_257; // @[RegisterRouter.scala 59:16]
  wire  _T_1176 = _T_1059 & _T_826[23]; // @[RegisterRouter.scala 59:16]
  wire  _T_1177 = _T_1176 & _T_131; // @[RegisterRouter.scala 59:16]
  wire  _T_701 = _T_1177 & _T_280; // @[RegisterRouter.scala 59:16]
  wire  _T_1101 = _T_1059 & _T_826[8]; // @[RegisterRouter.scala 59:16]
  wire  _T_1102 = _T_1101 & _T_131; // @[RegisterRouter.scala 59:16]
  wire  _T_724 = _T_1102 & _T_280; // @[RegisterRouter.scala 59:16]
  wire  _T_1156 = _T_1059 & _T_826[19]; // @[RegisterRouter.scala 59:16]
  wire  _T_1157 = _T_1156 & _T_131; // @[RegisterRouter.scala 59:16]
  wire  _T_747 = _T_1157 & _T_280; // @[RegisterRouter.scala 59:16]
  wire  _T_1081 = _T_1059 & _T_826[4]; // @[RegisterRouter.scala 59:16]
  wire  _T_1082 = _T_1081 & _T_131; // @[RegisterRouter.scala 59:16]
  wire  _T_770 = _T_1082 & _T_257; // @[RegisterRouter.scala 59:16]
  wire  _T_1136 = _T_1059 & _T_826[15]; // @[RegisterRouter.scala 59:16]
  wire  _T_1137 = _T_1136 & _T_131; // @[RegisterRouter.scala 59:16]
  wire  _T_793 = _T_1137 & _T_257; // @[RegisterRouter.scala 59:16]
  wire  _GEN_162 = 5'h1 == _T_825 ? _T_131 : _T_131; // @[MuxLiteral.scala 48:10]
  wire  _GEN_163 = 5'h2 == _T_825 ? _T_131 : _GEN_162; // @[MuxLiteral.scala 48:10]
  wire  _GEN_164 = 5'h3 == _T_825 ? _T_131 : _GEN_163; // @[MuxLiteral.scala 48:10]
  wire  _GEN_165 = 5'h4 == _T_825 ? _T_131 : _GEN_164; // @[MuxLiteral.scala 48:10]
  wire  _GEN_166 = 5'h5 == _T_825 ? _T_131 : _GEN_165; // @[MuxLiteral.scala 48:10]
  wire  _GEN_167 = 5'h6 == _T_825 ? _T_131 : _GEN_166; // @[MuxLiteral.scala 48:10]
  wire  _GEN_168 = 5'h7 == _T_825 ? _T_131 : _GEN_167; // @[MuxLiteral.scala 48:10]
  wire  _GEN_169 = 5'h8 == _T_825 ? _T_131 : _GEN_168; // @[MuxLiteral.scala 48:10]
  wire  _GEN_170 = 5'h9 == _T_825 ? _T_131 : _GEN_169; // @[MuxLiteral.scala 48:10]
  wire  _GEN_171 = 5'ha == _T_825 ? _T_131 : _GEN_170; // @[MuxLiteral.scala 48:10]
  wire  _GEN_172 = 5'hb == _T_825 ? _T_131 : _GEN_171; // @[MuxLiteral.scala 48:10]
  wire  _GEN_173 = 5'hc == _T_825 ? _T_131 : _GEN_172; // @[MuxLiteral.scala 48:10]
  wire  _GEN_174 = 5'hd == _T_825 ? _T_131 : _GEN_173; // @[MuxLiteral.scala 48:10]
  wire  _GEN_175 = 5'he == _T_825 ? _T_131 : _GEN_174; // @[MuxLiteral.scala 48:10]
  wire  _GEN_176 = 5'hf == _T_825 ? _T_131 : _GEN_175; // @[MuxLiteral.scala 48:10]
  wire  _GEN_177 = 5'h10 == _T_825 ? _T_131 : _GEN_176; // @[MuxLiteral.scala 48:10]
  wire  _GEN_178 = 5'h11 == _T_825 ? _T_131 : _GEN_177; // @[MuxLiteral.scala 48:10]
  wire  _GEN_179 = 5'h12 == _T_825 ? _T_131 : _GEN_178; // @[MuxLiteral.scala 48:10]
  wire  _GEN_180 = 5'h13 == _T_825 ? _T_131 : _GEN_179; // @[MuxLiteral.scala 48:10]
  wire  _GEN_181 = 5'h14 == _T_825 ? _T_131 : _GEN_180; // @[MuxLiteral.scala 48:10]
  wire  _GEN_182 = 5'h15 == _T_825 ? _T_131 : _GEN_181; // @[MuxLiteral.scala 48:10]
  wire  _GEN_183 = 5'h16 == _T_825 ? _T_131 : _GEN_182; // @[MuxLiteral.scala 48:10]
  wire  _GEN_184 = 5'h17 == _T_825 ? _T_131 : _GEN_183; // @[MuxLiteral.scala 48:10]
  wire  _GEN_185 = 5'h18 == _T_825 ? _T_131 : _GEN_184; // @[MuxLiteral.scala 48:10]
  wire  _GEN_186 = 5'h19 == _T_825 ? _T_131 : _GEN_185; // @[MuxLiteral.scala 48:10]
  wire  _GEN_351 = 5'h1a == _T_825; // @[MuxLiteral.scala 48:10]
  wire  _GEN_187 = _GEN_351 | _GEN_186; // @[MuxLiteral.scala 48:10]
  wire  _GEN_352 = 5'h1b == _T_825; // @[MuxLiteral.scala 48:10]
  wire  _GEN_188 = _GEN_352 | _GEN_187; // @[MuxLiteral.scala 48:10]
  wire  _GEN_353 = 5'h1c == _T_825; // @[MuxLiteral.scala 48:10]
  wire  _GEN_189 = _GEN_353 | _GEN_188; // @[MuxLiteral.scala 48:10]
  wire  _GEN_354 = 5'h1d == _T_825; // @[MuxLiteral.scala 48:10]
  wire  _GEN_190 = _GEN_354 | _GEN_189; // @[MuxLiteral.scala 48:10]
  wire  _GEN_355 = 5'h1e == _T_825; // @[MuxLiteral.scala 48:10]
  wire  _GEN_191 = _GEN_355 | _GEN_190; // @[MuxLiteral.scala 48:10]
  wire  _GEN_356 = 5'h1f == _T_825; // @[MuxLiteral.scala 48:10]
  wire  _GEN_192 = _GEN_356 | _GEN_191; // @[MuxLiteral.scala 48:10]
  wire [15:0] _T_1564_0 = {{15'd0}, enable}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [15:0] _T_1564_1 = {{15'd0}, reset_bit}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [15:0] _GEN_194 = 5'h1 == _T_825 ? _T_1564_1 : _T_1564_0; // @[MuxLiteral.scala 48:10]
  wire [15:0] _T_1564_2 = {{14'd0}, frameNum}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [15:0] _GEN_195 = 5'h2 == _T_825 ? _T_1564_2 : _GEN_194; // @[MuxLiteral.scala 48:10]
  wire [15:0] _T_1564_3 = {{6'd0}, _T_620}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [15:0] _GEN_196 = 5'h3 == _T_825 ? _T_1564_3 : _GEN_195; // @[MuxLiteral.scala 48:10]
  wire [15:0] _T_1564_4 = {{13'd0}, differentChirpsNum}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [15:0] _GEN_197 = 5'h4 == _T_825 ? _T_1564_4 : _GEN_196; // @[MuxLiteral.scala 48:10]
  wire [15:0] _GEN_198 = 5'h5 == _T_825 ? startingPoint : _GEN_197; // @[MuxLiteral.scala 48:10]
  wire [15:0] _T_1564_6 = {{14'd0}, segmentNums_0}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [15:0] _GEN_199 = 5'h6 == _T_825 ? _T_1564_6 : _GEN_198; // @[MuxLiteral.scala 48:10]
  wire [15:0] _T_1564_7 = {{14'd0}, segmentNums_1}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [15:0] _GEN_200 = 5'h7 == _T_825 ? _T_1564_7 : _GEN_199; // @[MuxLiteral.scala 48:10]
  wire [15:0] _T_1564_8 = {{14'd0}, segmentNums_2}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [15:0] _GEN_201 = 5'h8 == _T_825 ? _T_1564_8 : _GEN_200; // @[MuxLiteral.scala 48:10]
  wire [15:0] _T_1564_9 = {{14'd0}, segmentNums_3}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [15:0] _GEN_202 = 5'h9 == _T_825 ? _T_1564_9 : _GEN_201; // @[MuxLiteral.scala 48:10]
  wire [15:0] _T_1564_10 = {{13'd0}, repeatedChirpNums_0}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [15:0] _GEN_203 = 5'ha == _T_825 ? _T_1564_10 : _GEN_202; // @[MuxLiteral.scala 48:10]
  wire [15:0] _T_1564_11 = {{13'd0}, repeatedChirpNums_1}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [15:0] _GEN_204 = 5'hb == _T_825 ? _T_1564_11 : _GEN_203; // @[MuxLiteral.scala 48:10]
  wire [15:0] _T_1564_12 = {{13'd0}, repeatedChirpNums_2}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [15:0] _GEN_205 = 5'hc == _T_825 ? _T_1564_12 : _GEN_204; // @[MuxLiteral.scala 48:10]
  wire [15:0] _T_1564_13 = {{13'd0}, repeatedChirpNums_3}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [15:0] _GEN_206 = 5'hd == _T_825 ? _T_1564_13 : _GEN_205; // @[MuxLiteral.scala 48:10]
  wire [15:0] _T_1564_14 = {{13'd0}, repeatedChirpNums_4}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [15:0] _GEN_207 = 5'he == _T_825 ? _T_1564_14 : _GEN_206; // @[MuxLiteral.scala 48:10]
  wire [15:0] _T_1564_15 = {{13'd0}, repeatedChirpNums_5}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [15:0] _GEN_208 = 5'hf == _T_825 ? _T_1564_15 : _GEN_207; // @[MuxLiteral.scala 48:10]
  wire [15:0] _T_1564_16 = {{13'd0}, repeatedChirpNums_6}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [15:0] _GEN_209 = 5'h10 == _T_825 ? _T_1564_16 : _GEN_208; // @[MuxLiteral.scala 48:10]
  wire [15:0] _T_1564_17 = {{13'd0}, repeatedChirpNums_7}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [15:0] _GEN_210 = 5'h11 == _T_825 ? _T_1564_17 : _GEN_209; // @[MuxLiteral.scala 48:10]
  wire [15:0] _T_1564_18 = {{14'd0}, chirpOrdinalNums_0}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [15:0] _GEN_211 = 5'h12 == _T_825 ? _T_1564_18 : _GEN_210; // @[MuxLiteral.scala 48:10]
  wire [15:0] _T_1564_19 = {{14'd0}, chirpOrdinalNums_1}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [15:0] _GEN_212 = 5'h13 == _T_825 ? _T_1564_19 : _GEN_211; // @[MuxLiteral.scala 48:10]
  wire [15:0] _T_1564_20 = {{14'd0}, chirpOrdinalNums_2}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [15:0] _GEN_213 = 5'h14 == _T_825 ? _T_1564_20 : _GEN_212; // @[MuxLiteral.scala 48:10]
  wire [15:0] _T_1564_21 = {{14'd0}, chirpOrdinalNums_3}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [15:0] _GEN_214 = 5'h15 == _T_825 ? _T_1564_21 : _GEN_213; // @[MuxLiteral.scala 48:10]
  wire [15:0] _T_1564_22 = {{14'd0}, chirpOrdinalNums_4}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [15:0] _GEN_215 = 5'h16 == _T_825 ? _T_1564_22 : _GEN_214; // @[MuxLiteral.scala 48:10]
  wire [15:0] _T_1564_23 = {{14'd0}, chirpOrdinalNums_5}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [15:0] _GEN_216 = 5'h17 == _T_825 ? _T_1564_23 : _GEN_215; // @[MuxLiteral.scala 48:10]
  wire [15:0] _T_1564_24 = {{14'd0}, chirpOrdinalNums_6}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [15:0] _GEN_217 = 5'h18 == _T_825 ? _T_1564_24 : _GEN_216; // @[MuxLiteral.scala 48:10]
  wire [15:0] _T_1564_25 = {{14'd0}, chirpOrdinalNums_7}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [15:0] _GEN_218 = 5'h19 == _T_825 ? _T_1564_25 : _GEN_217; // @[MuxLiteral.scala 48:10]
  wire [15:0] _GEN_219 = 5'h1a == _T_825 ? 16'h0 : _GEN_218; // @[MuxLiteral.scala 48:10]
  wire [15:0] _GEN_220 = 5'h1b == _T_825 ? 16'h0 : _GEN_219; // @[MuxLiteral.scala 48:10]
  wire [15:0] _GEN_221 = 5'h1c == _T_825 ? 16'h0 : _GEN_220; // @[MuxLiteral.scala 48:10]
  wire [15:0] _GEN_222 = 5'h1d == _T_825 ? 16'h0 : _GEN_221; // @[MuxLiteral.scala 48:10]
  wire [15:0] _GEN_223 = 5'h1e == _T_825 ? 16'h0 : _GEN_222; // @[MuxLiteral.scala 48:10]
  wire [15:0] _GEN_224 = 5'h1f == _T_825 ? 16'h0 : _GEN_223; // @[MuxLiteral.scala 48:10]
  wire [15:0] _T_1566 = _GEN_192 ? _GEN_224 : 16'h0; // @[RegisterRouter.scala 59:16]
  wire  _T_1567_bits_read = Queue_io_deq_bits_read; // @[Decoupled.scala 317:19 Decoupled.scala 318:14]
  wire  _T_2_r_ready = axi4xbar_auto_out_1_r_ready; // @[Nodes.scala 370:76 LazyModule.scala 167:31]
  wire  _T_2_b_ready = axi4xbar_auto_out_1_b_ready; // @[Nodes.scala 370:76 LazyModule.scala 167:31]
  wire  _T_1567_valid = Queue_io_deq_valid; // @[Decoupled.scala 317:19 Decoupled.scala 319:15]
  wire  _T_1570 = ~_T_1567_bits_read; // @[RegisterRouter.scala 65:29]
  reg  enable2; // @[PLFGDspBlockMem.scala 218:26]
  reg [31:0] _RAND_46;
  reg [1:0] chirpIndexOld; // @[PLFGDspBlockMem.scala 219:32]
  reg [31:0] _RAND_47;
  reg  started; // @[PLFGDspBlockMem.scala 220:26]
  reg [31:0] _RAND_48;
  wire [1:0] _GEN_226 = 3'h1 == differentChirpsCounter ? chirpOrdinalNums_1 : chirpOrdinalNums_0; // @[PLFGDspBlockMem.scala 238:18]
  wire [1:0] _GEN_227 = 3'h2 == differentChirpsCounter ? chirpOrdinalNums_2 : _GEN_226; // @[PLFGDspBlockMem.scala 238:18]
  wire [1:0] _GEN_228 = 3'h3 == differentChirpsCounter ? chirpOrdinalNums_3 : _GEN_227; // @[PLFGDspBlockMem.scala 238:18]
  wire [1:0] _GEN_229 = 3'h4 == differentChirpsCounter ? chirpOrdinalNums_4 : _GEN_228; // @[PLFGDspBlockMem.scala 238:18]
  wire [1:0] _GEN_230 = 3'h5 == differentChirpsCounter ? chirpOrdinalNums_5 : _GEN_229; // @[PLFGDspBlockMem.scala 238:18]
  wire [1:0] _GEN_231 = 3'h6 == differentChirpsCounter ? chirpOrdinalNums_6 : _GEN_230; // @[PLFGDspBlockMem.scala 238:18]
  wire [1:0] _GEN_232 = 3'h7 == differentChirpsCounter ? chirpOrdinalNums_7 : _GEN_231; // @[PLFGDspBlockMem.scala 238:18]
  wire  _T_1573 = enable & auto_stream_out_ready; // @[PLFGDspBlockMem.scala 239:19]
  wire  _T_1574 = ~end_; // @[PLFGDspBlockMem.scala 239:35]
  wire  _T_1575 = _T_1573 & _T_1574; // @[PLFGDspBlockMem.scala 239:32]
  wire [7:0] _T_1577 = samplesCounter + 8'h1; // @[PLFGDspBlockMem.scala 241:30]
  wire  _T_1578 = _T_1577 >= numsOfSamples; // @[PLFGDspBlockMem.scala 241:37]
  wire [1:0] _T_1580 = segmentCounter + 2'h1; // @[PLFGDspBlockMem.scala 242:32]
  wire [1:0] chirpIndex = reset_bit ? 2'h0 : _GEN_232; // @[PLFGDspBlockMem.scala 224:20]
  wire [1:0] _GEN_234 = 2'h1 == chirpIndex ? segmentNums_1 : segmentNums_0; // @[PLFGDspBlockMem.scala 242:39]
  wire [1:0] _GEN_235 = 2'h2 == chirpIndex ? segmentNums_2 : _GEN_234; // @[PLFGDspBlockMem.scala 242:39]
  wire [1:0] _GEN_236 = 2'h3 == chirpIndex ? segmentNums_3 : _GEN_235; // @[PLFGDspBlockMem.scala 242:39]
  wire  _T_1581 = _T_1580 >= _GEN_236; // @[PLFGDspBlockMem.scala 242:39]
  wire [2:0] _T_1583 = repeatedChirpsCounter + 3'h1; // @[PLFGDspBlockMem.scala 243:41]
  wire [2:0] _GEN_238 = 3'h1 == differentChirpsCounter ? repeatedChirpNums_1 : repeatedChirpNums_0; // @[PLFGDspBlockMem.scala 243:48]
  wire [2:0] _GEN_239 = 3'h2 == differentChirpsCounter ? repeatedChirpNums_2 : _GEN_238; // @[PLFGDspBlockMem.scala 243:48]
  wire [2:0] _GEN_240 = 3'h3 == differentChirpsCounter ? repeatedChirpNums_3 : _GEN_239; // @[PLFGDspBlockMem.scala 243:48]
  wire [2:0] _GEN_241 = 3'h4 == differentChirpsCounter ? repeatedChirpNums_4 : _GEN_240; // @[PLFGDspBlockMem.scala 243:48]
  wire [2:0] _GEN_242 = 3'h5 == differentChirpsCounter ? repeatedChirpNums_5 : _GEN_241; // @[PLFGDspBlockMem.scala 243:48]
  wire [2:0] _GEN_243 = 3'h6 == differentChirpsCounter ? repeatedChirpNums_6 : _GEN_242; // @[PLFGDspBlockMem.scala 243:48]
  wire [2:0] _GEN_244 = 3'h7 == differentChirpsCounter ? repeatedChirpNums_7 : _GEN_243; // @[PLFGDspBlockMem.scala 243:48]
  wire  _T_1584 = _T_1583 >= _GEN_244; // @[PLFGDspBlockMem.scala 243:48]
  wire [2:0] _T_1586 = differentChirpsCounter + 3'h1; // @[PLFGDspBlockMem.scala 244:44]
  wire  _T_1587 = _T_1586 >= differentChirpsNum; // @[PLFGDspBlockMem.scala 244:51]
  wire  _T_1590 = frameNum == 2'h0; // @[PLFGDspBlockMem.scala 245:31]
  wire [5:0] _T_1592 = framePauseCounter + 6'h1; // @[PLFGDspBlockMem.scala 247:43]
  wire [7:0] _GEN_357 = {{2'd0}, _T_1592}; // @[PLFGDspBlockMem.scala 247:50]
  wire  _T_1593 = _GEN_357 >= interframeNumOfSamples; // @[PLFGDspBlockMem.scala 247:50]
  wire [1:0] _T_1597 = frameCounter + 2'h1; // @[PLFGDspBlockMem.scala 258:38]
  wire  _T_1598 = _T_1597 >= frameNum; // @[PLFGDspBlockMem.scala 258:45]
  wire  _GEN_257 = _T_1598 | end_; // @[PLFGDspBlockMem.scala 258:57]
  wire  _T_1616 = enable2 & auto_stream_out_ready; // @[PLFGDspBlockMem.scala 298:20]
  wire  _T_1617 = ~end2; // @[PLFGDspBlockMem.scala 298:36]
  wire  _T_1618 = _T_1616 & _T_1617; // @[PLFGDspBlockMem.scala 298:33]
  wire [7:0] _T_1620 = samplesCounter2 + 8'h1; // @[PLFGDspBlockMem.scala 300:31]
  wire  _T_1621 = _T_1620 >= numsOfSamples; // @[PLFGDspBlockMem.scala 300:38]
  wire [1:0] _T_1623 = segmentCounter2 + 2'h1; // @[PLFGDspBlockMem.scala 301:34]
  wire [1:0] _GEN_318 = 2'h1 == chirpIndexOld ? segmentNums_1 : segmentNums_0; // @[PLFGDspBlockMem.scala 301:41]
  wire [1:0] _GEN_319 = 2'h2 == chirpIndexOld ? segmentNums_2 : _GEN_318; // @[PLFGDspBlockMem.scala 301:41]
  wire [1:0] _GEN_320 = 2'h3 == chirpIndexOld ? segmentNums_3 : _GEN_319; // @[PLFGDspBlockMem.scala 301:41]
  wire  _T_1626 = _T_1623 >= _GEN_320; // @[PLFGDspBlockMem.scala 301:41]
  wire [2:0] _T_1630 = repeatedChirpsCounter2 + 3'h1; // @[PLFGDspBlockMem.scala 303:42]
  wire  _T_1631 = _T_1630 >= _GEN_244; // @[PLFGDspBlockMem.scala 303:49]
  wire [2:0] _T_1633 = differentChirpsCounter2 + 3'h1; // @[PLFGDspBlockMem.scala 304:45]
  wire  _T_1634 = _T_1633 >= differentChirpsNum; // @[PLFGDspBlockMem.scala 304:52]
  wire  _T_1640 = frameCounter2 >= frameNum; // @[PLFGDspBlockMem.scala 309:38]
  wire  _GEN_321 = _T_1640 | end2; // @[PLFGDspBlockMem.scala 309:50]
  wire [15:0] _T_1652 = dataFromMem[15:0]; // @[PLFGDspBlockMem.scala 326:73]
  wire [15:0] _T_1655 = $signed(currentVal) + $signed(_T_1652); // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] _T_1660 = $signed(currentVal) - $signed(_T_1652); // @[FixedPointTypeClass.scala 30:68]
  wire  _T_1675 = ~started; // @[PLFGDspBlockMem.scala 337:14]
  wire  _GEN_336 = _T_1618 | started; // @[PLFGDspBlockMem.scala 298:42]
  wire [15:0] _GEN_342 = reset_bit ? startingPoint : currentVal; // @[PLFGDspBlockMem.scala 295:20]
  reg  _T_1679; // @[PLFGDspBlockMem.scala 345:39]
  reg [31:0] _RAND_49;
  wire  _T_1680 = ~_T_1679; // @[PLFGDspBlockMem.scala 345:31]
  wire  _T_1681 = enable2 & _T_1680; // @[PLFGDspBlockMem.scala 345:28]
  reg  lastOutReg; // @[PLFGDspBlockMem.scala 351:29]
  reg [31:0] _RAND_50;
  reg  _T_1682; // @[PLFGDspBlockMem.scala 352:25]
  reg [31:0] _RAND_51;
  wire  _T_1683 = ~_T_1682; // @[PLFGDspBlockMem.scala 352:17]
  wire  lastOut = end_ & _T_1683; // @[PLFGDspBlockMem.scala 352:14]
  reg  _T_1685; // @[PLFGDspBlockMem.scala 357:25]
  reg [31:0] _RAND_52;
  wire  _T_1686 = ~_T_1685; // @[PLFGDspBlockMem.scala 357:17]
  wire  _T_1687 = end_ & _T_1686; // @[PLFGDspBlockMem.scala 357:14]
  reg  _T_1688; // @[PLFGDspBlockMem.scala 359:36]
  reg [31:0] _RAND_53;
  wire  _T_1689 = auto_stream_out_ready & _T_1688; // @[PLFGDspBlockMem.scala 359:26]
  wire  _GEN_345 = _T_1689 ? 1'h0 : lastOutReg; // @[PLFGDspBlockMem.scala 359:42]
  wire  _GEN_346 = _T_1687 | _GEN_345; // @[PLFGDspBlockMem.scala 357:31]
  wire  _T_1691 = lastOut | lastOutReg; // @[PLFGDspBlockMem.scala 362:46]
  wire  _T_1693 = ~reset_bit; // @[PLFGDspBlockMem.scala 365:10]
  wire [2:0] _GEN_359 = {{1'd0}, chirpIndex}; // @[UIntTypeClass.scala 39:41]
  wire [4:0] _T_1694 = _GEN_359 * 3'h4; // @[UIntTypeClass.scala 39:41]
  wire [4:0] _GEN_360 = {{3'd0}, segmentCounter}; // @[PLFGDspBlockMem.scala 367:57]
  wire [4:0] _T_1696 = _T_1694 + _GEN_360; // @[PLFGDspBlockMem.scala 367:57]
  AXI4Xbar axi4xbar ( // @[Xbar.scala 211:30]
    .clock(axi4xbar_clock),
    .reset(axi4xbar_reset),
    .auto_in_aw_ready(axi4xbar_auto_in_aw_ready),
    .auto_in_aw_valid(axi4xbar_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4xbar_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4xbar_auto_in_aw_bits_addr),
    .auto_in_w_ready(axi4xbar_auto_in_w_ready),
    .auto_in_w_valid(axi4xbar_auto_in_w_valid),
    .auto_in_w_bits_data(axi4xbar_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi4xbar_auto_in_w_bits_strb),
    .auto_in_w_bits_last(axi4xbar_auto_in_w_bits_last),
    .auto_in_b_ready(axi4xbar_auto_in_b_ready),
    .auto_in_b_valid(axi4xbar_auto_in_b_valid),
    .auto_in_b_bits_resp(axi4xbar_auto_in_b_bits_resp),
    .auto_in_ar_ready(axi4xbar_auto_in_ar_ready),
    .auto_in_ar_valid(axi4xbar_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4xbar_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4xbar_auto_in_ar_bits_addr),
    .auto_in_ar_bits_size(axi4xbar_auto_in_ar_bits_size),
    .auto_in_r_ready(axi4xbar_auto_in_r_ready),
    .auto_in_r_valid(axi4xbar_auto_in_r_valid),
    .auto_in_r_bits_data(axi4xbar_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4xbar_auto_in_r_bits_resp),
    .auto_in_r_bits_last(axi4xbar_auto_in_r_bits_last),
    .auto_out_1_aw_ready(axi4xbar_auto_out_1_aw_ready),
    .auto_out_1_aw_valid(axi4xbar_auto_out_1_aw_valid),
    .auto_out_1_aw_bits_id(axi4xbar_auto_out_1_aw_bits_id),
    .auto_out_1_aw_bits_addr(axi4xbar_auto_out_1_aw_bits_addr),
    .auto_out_1_w_ready(axi4xbar_auto_out_1_w_ready),
    .auto_out_1_w_valid(axi4xbar_auto_out_1_w_valid),
    .auto_out_1_w_bits_data(axi4xbar_auto_out_1_w_bits_data),
    .auto_out_1_w_bits_strb(axi4xbar_auto_out_1_w_bits_strb),
    .auto_out_1_b_ready(axi4xbar_auto_out_1_b_ready),
    .auto_out_1_b_valid(axi4xbar_auto_out_1_b_valid),
    .auto_out_1_b_bits_id(axi4xbar_auto_out_1_b_bits_id),
    .auto_out_1_ar_ready(axi4xbar_auto_out_1_ar_ready),
    .auto_out_1_ar_valid(axi4xbar_auto_out_1_ar_valid),
    .auto_out_1_ar_bits_id(axi4xbar_auto_out_1_ar_bits_id),
    .auto_out_1_ar_bits_addr(axi4xbar_auto_out_1_ar_bits_addr),
    .auto_out_1_ar_bits_size(axi4xbar_auto_out_1_ar_bits_size),
    .auto_out_1_r_ready(axi4xbar_auto_out_1_r_ready),
    .auto_out_1_r_valid(axi4xbar_auto_out_1_r_valid),
    .auto_out_1_r_bits_id(axi4xbar_auto_out_1_r_bits_id),
    .auto_out_1_r_bits_data(axi4xbar_auto_out_1_r_bits_data),
    .auto_out_0_aw_ready(axi4xbar_auto_out_0_aw_ready),
    .auto_out_0_aw_valid(axi4xbar_auto_out_0_aw_valid),
    .auto_out_0_aw_bits_addr(axi4xbar_auto_out_0_aw_bits_addr),
    .auto_out_0_w_ready(axi4xbar_auto_out_0_w_ready),
    .auto_out_0_w_valid(axi4xbar_auto_out_0_w_valid),
    .auto_out_0_w_bits_data(axi4xbar_auto_out_0_w_bits_data),
    .auto_out_0_b_ready(axi4xbar_auto_out_0_b_ready),
    .auto_out_0_b_valid(axi4xbar_auto_out_0_b_valid)
  );
  Queue Queue ( // @[Decoupled.scala 296:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_read(Queue_io_enq_bits_read),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_extra(Queue_io_enq_bits_extra),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_read(Queue_io_deq_bits_read),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_extra(Queue_io_deq_bits_extra)
  );
  assign configParamsMem1__T_64_addr = configParamsMem1__T_64_addr_pipe_0;
  assign configParamsMem1__T_64_data = configParamsMem1[configParamsMem1__T_64_addr]; // @[PLFGDspBlockMem.scala 110:39]
  assign configParamsMem1__T_14_data = ramIn1_w_bits_data[25:0];
  assign configParamsMem1__T_14_addr = ramIn1_aw_bits_addr[5:2];
  assign configParamsMem1__T_14_mask = 1'h1;
  assign configParamsMem1__T_14_en = ramIn1_aw_ready & ramIn1_aw_valid;
  assign auto_mem_in_aw_ready = axi4xbar_auto_in_aw_ready; // @[LazyModule.scala 173:31]
  assign auto_mem_in_w_ready = axi4xbar_auto_in_w_ready; // @[LazyModule.scala 173:31]
  assign auto_mem_in_b_valid = axi4xbar_auto_in_b_valid; // @[LazyModule.scala 173:31]
  assign auto_mem_in_b_bits_resp = axi4xbar_auto_in_b_bits_resp; // @[LazyModule.scala 173:31]
  assign auto_mem_in_ar_ready = axi4xbar_auto_in_ar_ready; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_valid = axi4xbar_auto_in_r_valid; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_bits_data = axi4xbar_auto_in_r_bits_data; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_bits_resp = axi4xbar_auto_in_r_bits_resp; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_bits_last = axi4xbar_auto_in_r_bits_last; // @[LazyModule.scala 173:31]
  assign auto_stream_out_valid = auto_stream_out_ready ? _T_1681 : auto_stream_out_ready; // @[LazyModule.scala 173:49]
  assign auto_stream_out_bits_data = {{16'd0}, _GEN_342}; // @[LazyModule.scala 173:49]
  assign auto_stream_out_bits_last = auto_stream_out_ready & _T_1691; // @[LazyModule.scala 173:49]
  assign axi4xbar_clock = clock;
  assign axi4xbar_reset = reset;
  assign axi4xbar_auto_in_aw_valid = auto_mem_in_aw_valid; // @[LazyModule.scala 167:57]
  assign axi4xbar_auto_in_aw_bits_id = auto_mem_in_aw_bits_id; // @[LazyModule.scala 167:57]
  assign axi4xbar_auto_in_aw_bits_addr = auto_mem_in_aw_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4xbar_auto_in_w_valid = auto_mem_in_w_valid; // @[LazyModule.scala 167:57]
  assign axi4xbar_auto_in_w_bits_data = auto_mem_in_w_bits_data; // @[LazyModule.scala 167:57]
  assign axi4xbar_auto_in_w_bits_strb = auto_mem_in_w_bits_strb; // @[LazyModule.scala 167:57]
  assign axi4xbar_auto_in_w_bits_last = auto_mem_in_w_bits_last; // @[LazyModule.scala 167:57]
  assign axi4xbar_auto_in_b_ready = auto_mem_in_b_ready; // @[LazyModule.scala 167:57]
  assign axi4xbar_auto_in_ar_valid = auto_mem_in_ar_valid; // @[LazyModule.scala 167:57]
  assign axi4xbar_auto_in_ar_bits_id = auto_mem_in_ar_bits_id; // @[LazyModule.scala 167:57]
  assign axi4xbar_auto_in_ar_bits_addr = auto_mem_in_ar_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4xbar_auto_in_ar_bits_size = auto_mem_in_ar_bits_size; // @[LazyModule.scala 167:57]
  assign axi4xbar_auto_in_r_ready = auto_mem_in_r_ready; // @[LazyModule.scala 167:57]
  assign axi4xbar_auto_out_1_aw_ready = _T_75 & _T_2_w_valid; // @[LazyModule.scala 167:31]
  assign axi4xbar_auto_out_1_w_ready = _T_75 & _T_2_aw_valid; // @[LazyModule.scala 167:31]
  assign axi4xbar_auto_out_1_b_valid = _T_1567_valid & _T_1570; // @[LazyModule.scala 167:31]
  assign axi4xbar_auto_out_1_b_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 167:31]
  assign axi4xbar_auto_out_1_ar_ready = Queue_io_enq_ready; // @[LazyModule.scala 167:31]
  assign axi4xbar_auto_out_1_r_valid = _T_1567_valid & _T_1567_bits_read; // @[LazyModule.scala 167:31]
  assign axi4xbar_auto_out_1_r_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 167:31]
  assign axi4xbar_auto_out_1_r_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 167:31]
  assign axi4xbar_auto_out_0_aw_ready = ramIn1_w_valid & _T_6; // @[LazyModule.scala 167:31]
  assign axi4xbar_auto_out_0_w_ready = ramIn1_aw_valid & _T_6; // @[LazyModule.scala 167:31]
  assign axi4xbar_auto_out_0_b_valid = w_full1; // @[LazyModule.scala 167:31]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = _T_2_ar_valid | _T_72; // @[Decoupled.scala 297:22]
  assign Queue_io_enq_bits_read = axi4xbar_auto_out_1_ar_valid; // @[Decoupled.scala 298:21]
  assign Queue_io_enq_bits_data = {{16'd0}, _T_1566}; // @[Decoupled.scala 298:21]
  assign Queue_io_enq_bits_extra = _T_2_ar_valid ? _T_2_ar_bits_id : _T_2_aw_bits_id; // @[Decoupled.scala 298:21]
  assign Queue_io_deq_ready = _T_1567_bits_read ? _T_2_r_ready : _T_2_b_ready; // @[Decoupled.scala 320:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    configParamsMem1[initvar] = _RAND_0[25:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  configParamsMem1__T_64_en_pipe_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  configParamsMem1__T_64_addr_pipe_0 = _RAND_2[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  w_full1 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  enable = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  reset_bit = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  frameNum = _RAND_6[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  startingPoint = _RAND_7[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  interframeNumOfSamples = _RAND_8[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  differentChirpsNum = _RAND_9[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  currentVal = _RAND_10[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  samplesCounter = _RAND_11[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  segmentCounter = _RAND_12[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  frameCounter = _RAND_13[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  framePauseCounter = _RAND_14[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  end_ = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  samplesCounter2 = _RAND_16[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  segmentCounter2 = _RAND_17[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  frameCounter2 = _RAND_18[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  end2 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  repeatedChirpsCounter = _RAND_20[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  differentChirpsCounter = _RAND_21[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_19 = _RAND_22[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  repeatedChirpsCounter2 = _RAND_23[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_20 = _RAND_24[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  differentChirpsCounter2 = _RAND_25[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  segmentNums_0 = _RAND_26[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  segmentNums_1 = _RAND_27[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  segmentNums_2 = _RAND_28[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  segmentNums_3 = _RAND_29[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  repeatedChirpNums_0 = _RAND_30[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  repeatedChirpNums_1 = _RAND_31[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  repeatedChirpNums_2 = _RAND_32[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  repeatedChirpNums_3 = _RAND_33[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  repeatedChirpNums_4 = _RAND_34[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  repeatedChirpNums_5 = _RAND_35[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  repeatedChirpNums_6 = _RAND_36[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  repeatedChirpNums_7 = _RAND_37[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  chirpOrdinalNums_0 = _RAND_38[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  chirpOrdinalNums_1 = _RAND_39[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  chirpOrdinalNums_2 = _RAND_40[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  chirpOrdinalNums_3 = _RAND_41[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  chirpOrdinalNums_4 = _RAND_42[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  chirpOrdinalNums_5 = _RAND_43[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  chirpOrdinalNums_6 = _RAND_44[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  chirpOrdinalNums_7 = _RAND_45[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  enable2 = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  chirpIndexOld = _RAND_47[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  started = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  _T_1679 = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  lastOutReg = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  _T_1682 = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  _T_1685 = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  _T_1688 = _RAND_53[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(configParamsMem1__T_14_en & configParamsMem1__T_14_mask) begin
      configParamsMem1[configParamsMem1__T_14_addr] <= configParamsMem1__T_14_data; // @[PLFGDspBlockMem.scala 110:39]
    end
    configParamsMem1__T_64_en_pipe_0 <= 1'h1;
    if (_T_1693) begin
      if (enable) begin
        configParamsMem1__T_64_addr_pipe_0 <= _T_1696[3:0];
      end else begin
        configParamsMem1__T_64_addr_pipe_0 <= 4'h0;
      end
    end else begin
      configParamsMem1__T_64_addr_pipe_0 <= 4'h0;
    end
    if (reset) begin
      w_full1 <= 1'h0;
    end else begin
      w_full1 <= _GEN_1;
    end
    if (reset) begin
      enable <= 1'h0;
    end else if (_T_218) begin
      enable <= _T_2_w_bits_data[0];
    end
    if (reset) begin
      reset_bit <= 1'h0;
    end else if (_T_379) begin
      reset_bit <= _T_2_w_bits_data[0];
    end
    if (reset) begin
      frameNum <= 2'h1;
    end else if (_T_494) begin
      frameNum <= _T_2_w_bits_data[1:0];
    end
    if (reset) begin
      startingPoint <= 16'h0;
    end else if (_T_241) begin
      startingPoint <= _T_2_w_bits_data[15:0];
    end
    if (reset) begin
      interframeNumOfSamples <= 8'h0;
    end else begin
      interframeNumOfSamples <= _GEN_24[7:0];
    end
    if (reset) begin
      differentChirpsNum <= 3'h1;
    end else if (_T_770) begin
      differentChirpsNum <= _T_2_w_bits_data[2:0];
    end
    if (reset) begin
      currentVal <= startingPoint;
    end else if (reset_bit) begin
      currentVal <= startingPoint;
    end else if (_T_1618) begin
      if (_T_1621) begin
        if (_T_1626) begin
          if (_T_1631) begin
            if (_T_1634) begin
              if (_T_1590) begin
                currentVal <= startingPoint;
              end else if (_T_1640) begin
                currentVal <= startingPoint;
              end else begin
                currentVal <= startingPoint;
              end
            end else begin
              currentVal <= startingPoint;
            end
          end else begin
            currentVal <= startingPoint;
          end
        end else if (segmentResets) begin
          currentVal <= startingPoint;
        end else if (slopeSigns) begin
          currentVal <= _T_1655;
        end else begin
          currentVal <= _T_1660;
        end
      end else if (segmentResets) begin
        currentVal <= startingPoint;
      end else if (slopeSigns) begin
        currentVal <= _T_1655;
      end else begin
        currentVal <= _T_1660;
      end
    end else if (_T_1675) begin
      currentVal <= startingPoint;
    end
    if (reset) begin
      samplesCounter <= 8'h0;
    end else if (reset_bit) begin
      samplesCounter <= 8'h0;
    end else if (_T_1575) begin
      if (_T_1578) begin
        if (_T_1581) begin
          if (_T_1584) begin
            if (_T_1587) begin
              if (_T_1590) begin
                if (_T_1593) begin
                  samplesCounter <= 8'h0;
                end
              end else if (!(_T_1598)) begin
                if (_T_1593) begin
                  samplesCounter <= 8'h0;
                end
              end
            end else begin
              samplesCounter <= 8'h0;
            end
          end else begin
            samplesCounter <= 8'h0;
          end
        end else begin
          samplesCounter <= 8'h0;
        end
      end else begin
        samplesCounter <= _T_1577;
      end
    end
    if (reset) begin
      segmentCounter <= 2'h0;
    end else if (reset_bit) begin
      segmentCounter <= 2'h0;
    end else if (_T_1575) begin
      if (_T_1578) begin
        if (_T_1581) begin
          if (_T_1584) begin
            if (_T_1587) begin
              if (_T_1590) begin
                if (_T_1593) begin
                  segmentCounter <= 2'h0;
                end
              end else if (!(_T_1598)) begin
                if (_T_1593) begin
                  segmentCounter <= 2'h0;
                end
              end
            end else begin
              segmentCounter <= 2'h0;
            end
          end else begin
            segmentCounter <= 2'h0;
          end
        end else begin
          segmentCounter <= _T_1580;
        end
      end
    end
    if (reset) begin
      frameCounter <= 2'h0;
    end else if (reset_bit) begin
      frameCounter <= 2'h0;
    end else if (_T_1575) begin
      if (_T_1578) begin
        if (_T_1581) begin
          if (_T_1584) begin
            if (_T_1587) begin
              if (_T_1590) begin
                if (_T_1593) begin
                  frameCounter <= 2'h0;
                end
              end else if (!(_T_1598)) begin
                if (_T_1593) begin
                  frameCounter <= _T_1597;
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      framePauseCounter <= 6'h0;
    end else if (reset_bit) begin
      framePauseCounter <= 6'h0;
    end else if (_T_1575) begin
      if (_T_1578) begin
        if (_T_1581) begin
          if (_T_1584) begin
            if (_T_1587) begin
              if (_T_1590) begin
                if (_T_1593) begin
                  framePauseCounter <= 6'h0;
                end else begin
                  framePauseCounter <= _T_1592;
                end
              end else if (!(_T_1598)) begin
                if (_T_1593) begin
                  framePauseCounter <= 6'h0;
                end else begin
                  framePauseCounter <= _T_1592;
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      end_ <= 1'h0;
    end else if (!(reset_bit)) begin
      if (_T_1575) begin
        if (_T_1578) begin
          if (_T_1581) begin
            if (_T_1584) begin
              if (_T_1587) begin
                if (_T_1590) begin
                  end_ <= 1'h0;
                end else begin
                  end_ <= _GEN_257;
                end
              end
            end
          end
        end
      end
    end
    samplesCounter2 <= samplesCounter;
    segmentCounter2 <= segmentCounter;
    frameCounter2 <= frameCounter;
    if (reset) begin
      end2 <= 1'h0;
    end else if (!(reset_bit)) begin
      if (_T_1618) begin
        if (_T_1621) begin
          if (_T_1626) begin
            if (_T_1631) begin
              if (_T_1634) begin
                if (_T_1590) begin
                  end2 <= 1'h0;
                end else begin
                  end2 <= _GEN_321;
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      repeatedChirpsCounter <= 3'h0;
    end else if (reset_bit) begin
      repeatedChirpsCounter <= 3'h0;
    end else if (_T_1575) begin
      if (_T_1578) begin
        if (_T_1581) begin
          if (_T_1584) begin
            if (_T_1587) begin
              if (_T_1590) begin
                if (_T_1593) begin
                  repeatedChirpsCounter <= 3'h0;
                end
              end else if (!(_T_1598)) begin
                if (_T_1593) begin
                  repeatedChirpsCounter <= 3'h0;
                end
              end
            end else begin
              repeatedChirpsCounter <= 3'h0;
            end
          end else begin
            repeatedChirpsCounter <= _T_1583;
          end
        end
      end
    end
    if (reset) begin
      differentChirpsCounter <= 3'h0;
    end else if (reset_bit) begin
      differentChirpsCounter <= 3'h0;
    end else if (_T_1575) begin
      if (_T_1578) begin
        if (_T_1581) begin
          if (_T_1584) begin
            if (_T_1587) begin
              if (_T_1590) begin
                if (_T_1593) begin
                  differentChirpsCounter <= 3'h0;
                end
              end else if (!(_T_1598)) begin
                if (_T_1593) begin
                  differentChirpsCounter <= 3'h0;
                end
              end
            end else begin
              differentChirpsCounter <= _T_1586;
            end
          end
        end
      end
    end
    _T_19 <= repeatedChirpsCounter;
    repeatedChirpsCounter2 <= _T_19;
    _T_20 <= differentChirpsCounter;
    differentChirpsCounter2 <= _T_20;
    if (reset) begin
      segmentNums_0 <= 2'h0;
    end else if (_T_402) begin
      segmentNums_0 <= _T_2_w_bits_data[1:0];
    end
    if (reset) begin
      segmentNums_1 <= 2'h0;
    end else if (_T_586) begin
      segmentNums_1 <= _T_2_w_bits_data[1:0];
    end
    if (reset) begin
      segmentNums_2 <= 2'h0;
    end else if (_T_724) begin
      segmentNums_2 <= _T_2_w_bits_data[1:0];
    end
    if (reset) begin
      segmentNums_3 <= 2'h0;
    end else if (_T_448) begin
      segmentNums_3 <= _T_2_w_bits_data[1:0];
    end
    if (reset) begin
      repeatedChirpNums_0 <= 3'h0;
    end else if (_T_264) begin
      repeatedChirpNums_0 <= _T_2_w_bits_data[2:0];
    end
    if (reset) begin
      repeatedChirpNums_1 <= 3'h0;
    end else if (_T_678) begin
      repeatedChirpNums_1 <= _T_2_w_bits_data[2:0];
    end
    if (reset) begin
      repeatedChirpNums_2 <= 3'h0;
    end else if (_T_563) begin
      repeatedChirpNums_2 <= _T_2_w_bits_data[2:0];
    end
    if (reset) begin
      repeatedChirpNums_3 <= 3'h0;
    end else if (_T_471) begin
      repeatedChirpNums_3 <= _T_2_w_bits_data[2:0];
    end
    if (reset) begin
      repeatedChirpNums_4 <= 3'h0;
    end else if (_T_333) begin
      repeatedChirpNums_4 <= _T_2_w_bits_data[2:0];
    end
    if (reset) begin
      repeatedChirpNums_5 <= 3'h0;
    end else if (_T_793) begin
      repeatedChirpNums_5 <= _T_2_w_bits_data[2:0];
    end
    if (reset) begin
      repeatedChirpNums_6 <= 3'h0;
    end else if (_T_655) begin
      repeatedChirpNums_6 <= _T_2_w_bits_data[2:0];
    end
    if (reset) begin
      repeatedChirpNums_7 <= 3'h0;
    end else if (_T_517) begin
      repeatedChirpNums_7 <= _T_2_w_bits_data[2:0];
    end
    if (reset) begin
      chirpOrdinalNums_0 <= 2'h0;
    end else if (_T_632) begin
      chirpOrdinalNums_0 <= _T_2_w_bits_data[1:0];
    end
    if (reset) begin
      chirpOrdinalNums_1 <= 2'h0;
    end else if (_T_747) begin
      chirpOrdinalNums_1 <= _T_2_w_bits_data[1:0];
    end
    if (reset) begin
      chirpOrdinalNums_2 <= 2'h0;
    end else if (_T_356) begin
      chirpOrdinalNums_2 <= _T_2_w_bits_data[1:0];
    end
    if (reset) begin
      chirpOrdinalNums_3 <= 2'h0;
    end else if (_T_425) begin
      chirpOrdinalNums_3 <= _T_2_w_bits_data[1:0];
    end
    if (reset) begin
      chirpOrdinalNums_4 <= 2'h0;
    end else if (_T_540) begin
      chirpOrdinalNums_4 <= _T_2_w_bits_data[1:0];
    end
    if (reset) begin
      chirpOrdinalNums_5 <= 2'h0;
    end else if (_T_701) begin
      chirpOrdinalNums_5 <= _T_2_w_bits_data[1:0];
    end
    if (reset) begin
      chirpOrdinalNums_6 <= 2'h0;
    end else if (_T_287) begin
      chirpOrdinalNums_6 <= _T_2_w_bits_data[1:0];
    end
    if (reset) begin
      chirpOrdinalNums_7 <= 2'h0;
    end else if (_T_310) begin
      chirpOrdinalNums_7 <= _T_2_w_bits_data[1:0];
    end
    enable2 <= enable;
    if (reset_bit) begin
      chirpIndexOld <= 2'h0;
    end else if (3'h7 == differentChirpsCounter) begin
      chirpIndexOld <= chirpOrdinalNums_7;
    end else if (3'h6 == differentChirpsCounter) begin
      chirpIndexOld <= chirpOrdinalNums_6;
    end else if (3'h5 == differentChirpsCounter) begin
      chirpIndexOld <= chirpOrdinalNums_5;
    end else if (3'h4 == differentChirpsCounter) begin
      chirpIndexOld <= chirpOrdinalNums_4;
    end else if (3'h3 == differentChirpsCounter) begin
      chirpIndexOld <= chirpOrdinalNums_3;
    end else if (3'h2 == differentChirpsCounter) begin
      chirpIndexOld <= chirpOrdinalNums_2;
    end else if (3'h1 == differentChirpsCounter) begin
      chirpIndexOld <= chirpOrdinalNums_1;
    end else begin
      chirpIndexOld <= chirpOrdinalNums_0;
    end
    if (reset) begin
      started <= 1'h0;
    end else if (!(reset_bit)) begin
      started <= _GEN_336;
    end
    _T_1679 <= end_;
    if (reset) begin
      lastOutReg <= 1'h0;
    end else begin
      lastOutReg <= _GEN_346;
    end
    _T_1682 <= end_;
    _T_1685 <= end_;
    _T_1688 <= end_;
  end
endmodule
module AXI4Splitter_1(
  input         clock,
  input         reset,
  output        auto_mem_in_aw_ready,
  input         auto_mem_in_aw_valid,
  input         auto_mem_in_aw_bits_id,
  input  [29:0] auto_mem_in_aw_bits_addr,
  output        auto_mem_in_w_ready,
  input         auto_mem_in_w_valid,
  input  [31:0] auto_mem_in_w_bits_data,
  input  [3:0]  auto_mem_in_w_bits_strb,
  input         auto_mem_in_b_ready,
  output        auto_mem_in_b_valid,
  output        auto_mem_in_b_bits_id,
  output        auto_mem_in_ar_ready,
  input         auto_mem_in_ar_valid,
  input         auto_mem_in_ar_bits_id,
  input  [29:0] auto_mem_in_ar_bits_addr,
  input  [2:0]  auto_mem_in_ar_bits_size,
  input         auto_mem_in_r_ready,
  output        auto_mem_in_r_valid,
  output        auto_mem_in_r_bits_id,
  output [31:0] auto_mem_in_r_bits_data,
  output        auto_stream_in_ready,
  input         auto_stream_in_valid,
  input  [31:0] auto_stream_in_bits_data,
  input         auto_stream_in_bits_last,
  input         auto_stream_out_1_ready,
  output        auto_stream_out_1_valid,
  output [31:0] auto_stream_out_1_bits_data,
  output        auto_stream_out_1_bits_last,
  input         auto_stream_out_0_ready,
  output        auto_stream_out_0_valid,
  output [31:0] auto_stream_out_0_bits_data,
  output        auto_stream_out_0_bits_last
);
  wire  Queue_clock; // @[Decoupled.scala 296:21]
  wire  Queue_reset; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_bits_read; // @[Decoupled.scala 296:21]
  wire [31:0] Queue_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_bits_extra; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_bits_read; // @[Decoupled.scala 296:21]
  wire [31:0] Queue_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_bits_extra; // @[Decoupled.scala 296:21]
  reg [31:0] ctrlReg; // @[Splitter.scala 27:26]
  reg [31:0] _RAND_0;
  reg [31:0] maskReg; // @[Splitter.scala 28:26]
  reg [31:0] _RAND_1;
  wire  _T_4 = auto_mem_in_aw_valid & auto_mem_in_w_valid; // @[RegisterRouter.scala 40:39]
  wire  _T_5 = auto_mem_in_ar_valid | _T_4; // @[RegisterRouter.scala 40:26]
  wire  _T_6 = ~auto_mem_in_ar_valid; // @[RegisterRouter.scala 42:29]
  wire  _T_49_ready = Queue_io_enq_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 299:17]
  wire [29:0] _T_13 = auto_mem_in_ar_valid ? auto_mem_in_ar_bits_addr : auto_mem_in_aw_bits_addr; // @[RegisterRouter.scala 48:19]
  wire [1:0] _T_53 = _T_13[3:2] & 2'h2; // @[RegisterRouter.scala 59:16]
  wire  _T_55 = _T_53 == 2'h0; // @[RegisterRouter.scala 59:16]
  wire  _T_7 = _T_49_ready & _T_6; // @[RegisterRouter.scala 42:26]
  wire [1:0] _T_16 = 2'h1 << auto_mem_in_ar_bits_size[0]; // @[OneHot.scala 65:12]
  wire [1:0] _T_18 = _T_16 | 2'h1; // @[Misc.scala 200:81]
  wire  _T_19 = auto_mem_in_ar_bits_size >= 3'h2; // @[Misc.scala 204:21]
  wire  _T_22 = ~auto_mem_in_ar_bits_addr[1]; // @[Misc.scala 209:20]
  wire  _T_24 = _T_18[1] & _T_22; // @[Misc.scala 213:38]
  wire  _T_25 = _T_19 | _T_24; // @[Misc.scala 213:29]
  wire  _T_27 = _T_18[1] & auto_mem_in_ar_bits_addr[1]; // @[Misc.scala 213:38]
  wire  _T_28 = _T_19 | _T_27; // @[Misc.scala 213:29]
  wire  _T_31 = ~auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 209:20]
  wire  _T_32 = _T_22 & _T_31; // @[Misc.scala 212:27]
  wire  _T_33 = _T_18[0] & _T_32; // @[Misc.scala 213:38]
  wire  _T_34 = _T_25 | _T_33; // @[Misc.scala 213:29]
  wire  _T_35 = _T_22 & auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  wire  _T_36 = _T_18[0] & _T_35; // @[Misc.scala 213:38]
  wire  _T_37 = _T_25 | _T_36; // @[Misc.scala 213:29]
  wire  _T_38 = auto_mem_in_ar_bits_addr[1] & _T_31; // @[Misc.scala 212:27]
  wire  _T_39 = _T_18[0] & _T_38; // @[Misc.scala 213:38]
  wire  _T_40 = _T_28 | _T_39; // @[Misc.scala 213:29]
  wire  _T_41 = auto_mem_in_ar_bits_addr[1] & auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  wire  _T_42 = _T_18[0] & _T_41; // @[Misc.scala 213:38]
  wire  _T_43 = _T_28 | _T_42; // @[Misc.scala 213:29]
  wire [3:0] _T_46 = {_T_43,_T_40,_T_37,_T_34}; // @[Cat.scala 29:58]
  wire [3:0] _T_48 = auto_mem_in_ar_valid ? _T_46 : auto_mem_in_w_bits_strb; // @[RegisterRouter.scala 54:25]
  wire [7:0] _T_67 = _T_48[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_69 = _T_48[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_71 = _T_48[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_73 = _T_48[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_76 = {_T_73,_T_71,_T_69,_T_67}; // @[Cat.scala 29:58]
  wire  _T_95 = _T_76 == 32'hffffffff; // @[RegisterRouter.scala 59:16]
  wire  _T_148 = _T_5 & _T_49_ready; // @[RegisterRouter.scala 59:16]
  wire [1:0] _T_142 = 2'h1 << _T_13[2]; // @[OneHot.scala 58:35]
  wire  _T_165 = _T_148 & _T_6; // @[RegisterRouter.scala 59:16]
  wire  _T_172 = _T_165 & _T_142[1]; // @[RegisterRouter.scala 59:16]
  wire  _T_173 = _T_172 & _T_55; // @[RegisterRouter.scala 59:16]
  wire  _T_102 = _T_173 & _T_95; // @[RegisterRouter.scala 59:16]
  wire  _T_167 = _T_165 & _T_142[0]; // @[RegisterRouter.scala 59:16]
  wire  _T_168 = _T_167 & _T_55; // @[RegisterRouter.scala 59:16]
  wire  _T_125 = _T_168 & _T_95; // @[RegisterRouter.scala 59:16]
  wire  _GEN_11 = _T_13[2] ? _T_55 : _T_55; // @[MuxLiteral.scala 48:10]
  wire [31:0] _GEN_13 = _T_13[2] ? maskReg : ctrlReg; // @[MuxLiteral.scala 48:10]
  wire  _T_223_bits_read = Queue_io_deq_bits_read; // @[Decoupled.scala 317:19 Decoupled.scala 318:14]
  wire  _T_223_valid = Queue_io_deq_valid; // @[Decoupled.scala 317:19 Decoupled.scala 319:15]
  wire  _T_226 = ~_T_223_bits_read; // @[RegisterRouter.scala 65:29]
  wire  readyOR = auto_stream_out_0_ready | auto_stream_out_1_ready; // @[Splitter.scala 45:34]
  wire  readyAND = auto_stream_out_0_ready & auto_stream_out_1_ready; // @[Splitter.scala 46:34]
  wire  _T_229 = ctrlReg == 32'h0; // @[Splitter.scala 49:19]
  wire  _T_230 = ctrlReg == 32'h1; // @[Splitter.scala 52:24]
  wire  _GEN_14 = _T_230 & readyOR; // @[Splitter.scala 52:33]
  wire  _T_233 = ~maskReg[0]; // @[Splitter.scala 62:34]
  wire  _T_237 = ~maskReg[1]; // @[Splitter.scala 62:34]
  Queue Queue ( // @[Decoupled.scala 296:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_read(Queue_io_enq_bits_read),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_extra(Queue_io_enq_bits_extra),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_read(Queue_io_deq_bits_read),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_extra(Queue_io_deq_bits_extra)
  );
  assign auto_mem_in_aw_ready = _T_7 & auto_mem_in_w_valid; // @[LazyModule.scala 173:31]
  assign auto_mem_in_w_ready = _T_7 & auto_mem_in_aw_valid; // @[LazyModule.scala 173:31]
  assign auto_mem_in_b_valid = _T_223_valid & _T_226; // @[LazyModule.scala 173:31]
  assign auto_mem_in_b_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_mem_in_ar_ready = Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_valid = _T_223_valid & _T_223_bits_read; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 173:31]
  assign auto_stream_in_ready = _T_229 ? readyAND : _GEN_14; // @[LazyModule.scala 173:31]
  assign auto_stream_out_1_valid = auto_stream_in_valid & _T_237; // @[LazyModule.scala 173:49]
  assign auto_stream_out_1_bits_data = auto_stream_in_bits_data; // @[LazyModule.scala 173:49]
  assign auto_stream_out_1_bits_last = auto_stream_in_bits_last; // @[LazyModule.scala 173:49]
  assign auto_stream_out_0_valid = auto_stream_in_valid & _T_233; // @[LazyModule.scala 173:49]
  assign auto_stream_out_0_bits_data = auto_stream_in_bits_data; // @[LazyModule.scala 173:49]
  assign auto_stream_out_0_bits_last = auto_stream_in_bits_last; // @[LazyModule.scala 173:49]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_mem_in_ar_valid | _T_4; // @[Decoupled.scala 297:22]
  assign Queue_io_enq_bits_read = auto_mem_in_ar_valid; // @[Decoupled.scala 298:21]
  assign Queue_io_enq_bits_data = _GEN_11 ? _GEN_13 : 32'h0; // @[Decoupled.scala 298:21]
  assign Queue_io_enq_bits_extra = auto_mem_in_ar_valid ? auto_mem_in_ar_bits_id : auto_mem_in_aw_bits_id; // @[Decoupled.scala 298:21]
  assign Queue_io_deq_ready = _T_223_bits_read ? auto_mem_in_r_ready : auto_mem_in_b_ready; // @[Decoupled.scala 320:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ctrlReg = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  maskReg = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      ctrlReg <= 32'h0;
    end else if (_T_125) begin
      ctrlReg <= auto_mem_in_w_bits_data;
    end
    if (reset) begin
      maskReg <= 32'h0;
    end else if (_T_102) begin
      maskReg <= auto_mem_in_w_bits_data;
    end
  end
endmodule
module AXI4StreamMux(
  input         clock,
  input         reset,
  output        auto_register_in_aw_ready,
  input         auto_register_in_aw_valid,
  input         auto_register_in_aw_bits_id,
  input  [29:0] auto_register_in_aw_bits_addr,
  output        auto_register_in_w_ready,
  input         auto_register_in_w_valid,
  input  [31:0] auto_register_in_w_bits_data,
  input  [3:0]  auto_register_in_w_bits_strb,
  input         auto_register_in_b_ready,
  output        auto_register_in_b_valid,
  output        auto_register_in_b_bits_id,
  output        auto_register_in_ar_ready,
  input         auto_register_in_ar_valid,
  input         auto_register_in_ar_bits_id,
  input  [29:0] auto_register_in_ar_bits_addr,
  input  [2:0]  auto_register_in_ar_bits_size,
  input         auto_register_in_r_ready,
  output        auto_register_in_r_valid,
  output        auto_register_in_r_bits_id,
  output [31:0] auto_register_in_r_bits_data,
  output        auto_stream_in_2_ready,
  input         auto_stream_in_2_valid,
  input  [31:0] auto_stream_in_2_bits_data,
  input         auto_stream_in_2_bits_last,
  output        auto_stream_in_1_ready,
  input         auto_stream_in_1_valid,
  input  [31:0] auto_stream_in_1_bits_data,
  input         auto_stream_in_1_bits_last,
  output        auto_stream_in_0_ready,
  input         auto_stream_in_0_valid,
  input  [31:0] auto_stream_in_0_bits_data,
  input         auto_stream_in_0_bits_last,
  input         auto_stream_out_0_ready,
  output        auto_stream_out_0_valid,
  output [31:0] auto_stream_out_0_bits_data,
  output        auto_stream_out_0_bits_last
);
  wire  Queue_clock; // @[Decoupled.scala 296:21]
  wire  Queue_reset; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_bits_read; // @[Decoupled.scala 296:21]
  wire [31:0] Queue_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_bits_extra; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_bits_read; // @[Decoupled.scala 296:21]
  wire [31:0] Queue_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_bits_extra; // @[Decoupled.scala 296:21]
  reg [2:0] sels_0; // @[Mux.scala 32:23]
  reg [31:0] _RAND_0;
  reg [2:0] sels_1; // @[Mux.scala 32:23]
  reg [31:0] _RAND_1;
  wire  _T_3 = sels_0 == 3'h0; // @[Mux.scala 45:28]
  wire  _GEN_7 = _T_3 & auto_stream_in_0_valid; // @[Mux.scala 45:41]
  wire  _GEN_8 = _T_3 & auto_stream_out_0_ready; // @[Mux.scala 45:41]
  wire  _T_4 = sels_0 == 3'h1; // @[Mux.scala 45:28]
  wire  _GEN_12 = _T_4 ? auto_stream_in_1_bits_last : auto_stream_in_0_bits_last; // @[Mux.scala 45:41]
  wire [31:0] _GEN_15 = _T_4 ? auto_stream_in_1_bits_data : auto_stream_in_0_bits_data; // @[Mux.scala 45:41]
  wire  _GEN_16 = _T_4 ? auto_stream_in_1_valid : _GEN_7; // @[Mux.scala 45:41]
  wire  _GEN_17 = _T_4 & auto_stream_out_0_ready; // @[Mux.scala 45:41]
  wire  _T_5 = sels_0 == 3'h2; // @[Mux.scala 45:28]
  wire  _GEN_21 = _T_5 ? auto_stream_in_2_bits_last : _GEN_12; // @[Mux.scala 45:41]
  wire [31:0] _GEN_24 = _T_5 ? auto_stream_in_2_bits_data : _GEN_15; // @[Mux.scala 45:41]
  wire  _GEN_25 = _T_5 ? auto_stream_in_2_valid : _GEN_16; // @[Mux.scala 45:41]
  wire  _GEN_26 = _T_5 & auto_stream_out_0_ready; // @[Mux.scala 45:41]
  wire  _T_6 = sels_0 == 3'h3; // @[Mux.scala 45:28]
  wire  _GEN_30 = _T_6 ? 1'h0 : _GEN_21; // @[Mux.scala 45:41]
  wire [31:0] _GEN_33 = _T_6 ? 32'hffffffff : _GEN_24; // @[Mux.scala 45:41]
  wire  _GEN_34 = _T_6 | _GEN_25; // @[Mux.scala 45:41]
  wire  _T_7 = sels_0 == 3'h4; // @[Mux.scala 45:28]
  wire  _T_8 = sels_0 == sels_1; // @[Mux.scala 40:46]
  wire [2:0] _T_10 = _T_8 ? 3'h5 : sels_1; // @[Mux.scala 41:29]
  wire  _T_11 = _T_10 == 3'h0; // @[Mux.scala 45:28]
  wire  _T_12 = _T_10 == 3'h1; // @[Mux.scala 45:28]
  wire  _T_13 = _T_10 == 3'h2; // @[Mux.scala 45:28]
  wire  _T_17 = auto_register_in_aw_valid & auto_register_in_w_valid; // @[RegisterRouter.scala 40:39]
  wire  _T_18 = auto_register_in_ar_valid | _T_17; // @[RegisterRouter.scala 40:26]
  wire  _T_19 = ~auto_register_in_ar_valid; // @[RegisterRouter.scala 42:29]
  wire  _T_62_ready = Queue_io_enq_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 299:17]
  wire [29:0] _T_26 = auto_register_in_ar_valid ? auto_register_in_ar_bits_addr : auto_register_in_aw_bits_addr; // @[RegisterRouter.scala 48:19]
  wire [1:0] _T_66 = _T_26[3:2] & 2'h2; // @[RegisterRouter.scala 59:16]
  wire  _T_68 = _T_66 == 2'h0; // @[RegisterRouter.scala 59:16]
  wire  _T_20 = _T_62_ready & _T_19; // @[RegisterRouter.scala 42:26]
  wire [1:0] _T_29 = 2'h1 << auto_register_in_ar_bits_size[0]; // @[OneHot.scala 65:12]
  wire [1:0] _T_31 = _T_29 | 2'h1; // @[Misc.scala 200:81]
  wire  _T_32 = auto_register_in_ar_bits_size >= 3'h2; // @[Misc.scala 204:21]
  wire  _T_35 = ~auto_register_in_ar_bits_addr[1]; // @[Misc.scala 209:20]
  wire  _T_37 = _T_31[1] & _T_35; // @[Misc.scala 213:38]
  wire  _T_38 = _T_32 | _T_37; // @[Misc.scala 213:29]
  wire  _T_40 = _T_31[1] & auto_register_in_ar_bits_addr[1]; // @[Misc.scala 213:38]
  wire  _T_41 = _T_32 | _T_40; // @[Misc.scala 213:29]
  wire  _T_44 = ~auto_register_in_ar_bits_addr[0]; // @[Misc.scala 209:20]
  wire  _T_45 = _T_35 & _T_44; // @[Misc.scala 212:27]
  wire  _T_46 = _T_31[0] & _T_45; // @[Misc.scala 213:38]
  wire  _T_47 = _T_38 | _T_46; // @[Misc.scala 213:29]
  wire  _T_48 = _T_35 & auto_register_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  wire  _T_49 = _T_31[0] & _T_48; // @[Misc.scala 213:38]
  wire  _T_50 = _T_38 | _T_49; // @[Misc.scala 213:29]
  wire  _T_51 = auto_register_in_ar_bits_addr[1] & _T_44; // @[Misc.scala 212:27]
  wire  _T_52 = _T_31[0] & _T_51; // @[Misc.scala 213:38]
  wire  _T_53 = _T_41 | _T_52; // @[Misc.scala 213:29]
  wire  _T_54 = auto_register_in_ar_bits_addr[1] & auto_register_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  wire  _T_55 = _T_31[0] & _T_54; // @[Misc.scala 213:38]
  wire  _T_56 = _T_41 | _T_55; // @[Misc.scala 213:29]
  wire [3:0] _T_59 = {_T_56,_T_53,_T_50,_T_47}; // @[Cat.scala 29:58]
  wire [3:0] _T_61 = auto_register_in_ar_valid ? _T_59 : auto_register_in_w_bits_strb; // @[RegisterRouter.scala 54:25]
  wire [7:0] _T_80 = _T_61[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_82 = _T_61[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_84 = _T_61[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_86 = _T_61[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_89 = {_T_86,_T_84,_T_82,_T_80}; // @[Cat.scala 29:58]
  wire  _T_108 = _T_89[2:0] == 3'h7; // @[RegisterRouter.scala 59:16]
  wire  _T_161 = _T_18 & _T_62_ready; // @[RegisterRouter.scala 59:16]
  wire [1:0] _T_155 = 2'h1 << _T_26[2]; // @[OneHot.scala 58:35]
  wire  _T_178 = _T_161 & _T_19; // @[RegisterRouter.scala 59:16]
  wire  _T_185 = _T_178 & _T_155[1]; // @[RegisterRouter.scala 59:16]
  wire  _T_186 = _T_185 & _T_68; // @[RegisterRouter.scala 59:16]
  wire  _T_115 = _T_186 & _T_108; // @[RegisterRouter.scala 59:16]
  wire  _T_180 = _T_178 & _T_155[0]; // @[RegisterRouter.scala 59:16]
  wire  _T_181 = _T_180 & _T_68; // @[RegisterRouter.scala 59:16]
  wire  _T_138 = _T_181 & _T_108; // @[RegisterRouter.scala 59:16]
  wire  _GEN_101 = _T_26[2] ? _T_68 : _T_68; // @[MuxLiteral.scala 48:10]
  wire [2:0] _GEN_103 = _T_26[2] ? sels_1 : sels_0; // @[MuxLiteral.scala 48:10]
  wire [2:0] _T_235 = _GEN_101 ? _GEN_103 : 3'h0; // @[RegisterRouter.scala 59:16]
  wire  _T_236_bits_read = Queue_io_deq_bits_read; // @[Decoupled.scala 317:19 Decoupled.scala 318:14]
  wire  _T_236_valid = Queue_io_deq_valid; // @[Decoupled.scala 317:19 Decoupled.scala 319:15]
  wire  _T_239 = ~_T_236_bits_read; // @[RegisterRouter.scala 65:29]
  Queue Queue ( // @[Decoupled.scala 296:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_read(Queue_io_enq_bits_read),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_extra(Queue_io_enq_bits_extra),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_read(Queue_io_deq_bits_read),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_extra(Queue_io_deq_bits_extra)
  );
  assign auto_register_in_aw_ready = _T_20 & auto_register_in_w_valid; // @[LazyModule.scala 173:31]
  assign auto_register_in_w_ready = _T_20 & auto_register_in_aw_valid; // @[LazyModule.scala 173:31]
  assign auto_register_in_b_valid = _T_236_valid & _T_239; // @[LazyModule.scala 173:31]
  assign auto_register_in_b_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_register_in_ar_ready = Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_register_in_r_valid = _T_236_valid & _T_236_bits_read; // @[LazyModule.scala 173:31]
  assign auto_register_in_r_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_register_in_r_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 173:31]
  assign auto_stream_in_2_ready = _T_13 | _GEN_26; // @[LazyModule.scala 173:31]
  assign auto_stream_in_1_ready = _T_12 | _GEN_17; // @[LazyModule.scala 173:31]
  assign auto_stream_in_0_ready = _T_11 | _GEN_8; // @[LazyModule.scala 173:31]
  assign auto_stream_out_0_valid = _T_7 | _GEN_34; // @[LazyModule.scala 173:49]
  assign auto_stream_out_0_bits_data = _T_7 ? 32'h0 : _GEN_33; // @[LazyModule.scala 173:49]
  assign auto_stream_out_0_bits_last = _T_7 ? 1'h0 : _GEN_30; // @[LazyModule.scala 173:49]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_register_in_ar_valid | _T_17; // @[Decoupled.scala 297:22]
  assign Queue_io_enq_bits_read = auto_register_in_ar_valid; // @[Decoupled.scala 298:21]
  assign Queue_io_enq_bits_data = {{29'd0}, _T_235}; // @[Decoupled.scala 298:21]
  assign Queue_io_enq_bits_extra = auto_register_in_ar_valid ? auto_register_in_ar_bits_id : auto_register_in_aw_bits_id; // @[Decoupled.scala 298:21]
  assign Queue_io_deq_ready = _T_236_bits_read ? auto_register_in_r_ready : auto_register_in_b_ready; // @[Decoupled.scala 320:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  sels_0 = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  sels_1 = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      sels_0 <= 3'h5;
    end else if (_T_138) begin
      sels_0 <= auto_register_in_w_bits_data[2:0];
    end
    if (reset) begin
      sels_1 <= 3'h5;
    end else if (_T_115) begin
      sels_1 <= auto_register_in_w_bits_data[2:0];
    end
  end
endmodule
module AXI4StreamMux_1(
  input         clock,
  input         reset,
  output        auto_register_in_aw_ready,
  input         auto_register_in_aw_valid,
  input         auto_register_in_aw_bits_id,
  input  [29:0] auto_register_in_aw_bits_addr,
  output        auto_register_in_w_ready,
  input         auto_register_in_w_valid,
  input  [31:0] auto_register_in_w_bits_data,
  input  [3:0]  auto_register_in_w_bits_strb,
  input         auto_register_in_b_ready,
  output        auto_register_in_b_valid,
  output        auto_register_in_b_bits_id,
  output        auto_register_in_ar_ready,
  input         auto_register_in_ar_valid,
  input         auto_register_in_ar_bits_id,
  input  [29:0] auto_register_in_ar_bits_addr,
  input  [2:0]  auto_register_in_ar_bits_size,
  input         auto_register_in_r_ready,
  output        auto_register_in_r_valid,
  output        auto_register_in_r_bits_id,
  output [31:0] auto_register_in_r_bits_data,
  output        auto_stream_in_ready,
  input         auto_stream_in_valid,
  input  [31:0] auto_stream_in_bits_data,
  input         auto_stream_in_bits_last,
  input         auto_stream_out_1_ready,
  output        auto_stream_out_1_valid,
  output [31:0] auto_stream_out_1_bits_data,
  output        auto_stream_out_1_bits_last
);
  wire  Queue_clock; // @[Decoupled.scala 296:21]
  wire  Queue_reset; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_bits_read; // @[Decoupled.scala 296:21]
  wire [31:0] Queue_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_bits_extra; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_bits_read; // @[Decoupled.scala 296:21]
  wire [31:0] Queue_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_bits_extra; // @[Decoupled.scala 296:21]
  reg  sels_0; // @[Mux.scala 32:23]
  reg [31:0] _RAND_0;
  reg  sels_1; // @[Mux.scala 32:23]
  reg [31:0] _RAND_1;
  wire  _T_3 = ~sels_0; // @[Mux.scala 45:28]
  wire  _T_4 = sels_0 == sels_1; // @[Mux.scala 40:46]
  wire  _T_6 = _T_4 | sels_1; // @[Mux.scala 41:29]
  wire  _T_7 = ~_T_6; // @[Mux.scala 45:28]
  wire  _T_9 = auto_register_in_aw_valid & auto_register_in_w_valid; // @[RegisterRouter.scala 40:39]
  wire  _T_10 = auto_register_in_ar_valid | _T_9; // @[RegisterRouter.scala 40:26]
  wire  _T_11 = ~auto_register_in_ar_valid; // @[RegisterRouter.scala 42:29]
  wire  _T_54_ready = Queue_io_enq_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 299:17]
  wire [29:0] _T_18 = auto_register_in_ar_valid ? auto_register_in_ar_bits_addr : auto_register_in_aw_bits_addr; // @[RegisterRouter.scala 48:19]
  wire [1:0] _T_58 = _T_18[3:2] & 2'h2; // @[RegisterRouter.scala 59:16]
  wire  _T_60 = _T_58 == 2'h0; // @[RegisterRouter.scala 59:16]
  wire  _T_12 = _T_54_ready & _T_11; // @[RegisterRouter.scala 42:26]
  wire [1:0] _T_21 = 2'h1 << auto_register_in_ar_bits_size[0]; // @[OneHot.scala 65:12]
  wire [1:0] _T_23 = _T_21 | 2'h1; // @[Misc.scala 200:81]
  wire  _T_24 = auto_register_in_ar_bits_size >= 3'h2; // @[Misc.scala 204:21]
  wire  _T_27 = ~auto_register_in_ar_bits_addr[1]; // @[Misc.scala 209:20]
  wire  _T_29 = _T_23[1] & _T_27; // @[Misc.scala 213:38]
  wire  _T_30 = _T_24 | _T_29; // @[Misc.scala 213:29]
  wire  _T_32 = _T_23[1] & auto_register_in_ar_bits_addr[1]; // @[Misc.scala 213:38]
  wire  _T_33 = _T_24 | _T_32; // @[Misc.scala 213:29]
  wire  _T_36 = ~auto_register_in_ar_bits_addr[0]; // @[Misc.scala 209:20]
  wire  _T_37 = _T_27 & _T_36; // @[Misc.scala 212:27]
  wire  _T_38 = _T_23[0] & _T_37; // @[Misc.scala 213:38]
  wire  _T_39 = _T_30 | _T_38; // @[Misc.scala 213:29]
  wire  _T_40 = _T_27 & auto_register_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  wire  _T_41 = _T_23[0] & _T_40; // @[Misc.scala 213:38]
  wire  _T_42 = _T_30 | _T_41; // @[Misc.scala 213:29]
  wire  _T_43 = auto_register_in_ar_bits_addr[1] & _T_36; // @[Misc.scala 212:27]
  wire  _T_44 = _T_23[0] & _T_43; // @[Misc.scala 213:38]
  wire  _T_45 = _T_33 | _T_44; // @[Misc.scala 213:29]
  wire  _T_46 = auto_register_in_ar_bits_addr[1] & auto_register_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  wire  _T_47 = _T_23[0] & _T_46; // @[Misc.scala 213:38]
  wire  _T_48 = _T_33 | _T_47; // @[Misc.scala 213:29]
  wire [3:0] _T_51 = {_T_48,_T_45,_T_42,_T_39}; // @[Cat.scala 29:58]
  wire [3:0] _T_53 = auto_register_in_ar_valid ? _T_51 : auto_register_in_w_bits_strb; // @[RegisterRouter.scala 54:25]
  wire [7:0] _T_72 = _T_53[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_74 = _T_53[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_76 = _T_53[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_78 = _T_53[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_81 = {_T_78,_T_76,_T_74,_T_72}; // @[Cat.scala 29:58]
  wire  _T_153 = _T_10 & _T_54_ready; // @[RegisterRouter.scala 59:16]
  wire [1:0] _T_147 = 2'h1 << _T_18[2]; // @[OneHot.scala 58:35]
  wire  _T_170 = _T_153 & _T_11; // @[RegisterRouter.scala 59:16]
  wire  _T_177 = _T_170 & _T_147[1]; // @[RegisterRouter.scala 59:16]
  wire  _T_178 = _T_177 & _T_60; // @[RegisterRouter.scala 59:16]
  wire  _T_107 = _T_178 & _T_81[0]; // @[RegisterRouter.scala 59:16]
  wire  _GEN_18 = _T_107 ? auto_register_in_w_bits_data[0] : sels_1; // @[RegField.scala 134:88]
  wire  _T_172 = _T_170 & _T_147[0]; // @[RegisterRouter.scala 59:16]
  wire  _T_173 = _T_172 & _T_60; // @[RegisterRouter.scala 59:16]
  wire  _T_130 = _T_173 & _T_81[0]; // @[RegisterRouter.scala 59:16]
  wire  _GEN_19 = _T_130 ? auto_register_in_w_bits_data[0] : sels_0; // @[RegField.scala 134:88]
  wire  _GEN_29 = _T_18[2] ? _T_60 : _T_60; // @[MuxLiteral.scala 48:10]
  wire  _GEN_31 = _T_18[2] ? sels_1 : sels_0; // @[MuxLiteral.scala 48:10]
  wire  _T_227 = _GEN_29 & _GEN_31; // @[RegisterRouter.scala 59:16]
  wire  _T_228_bits_read = Queue_io_deq_bits_read; // @[Decoupled.scala 317:19 Decoupled.scala 318:14]
  wire  _T_228_valid = Queue_io_deq_valid; // @[Decoupled.scala 317:19 Decoupled.scala 319:15]
  wire  _T_231 = ~_T_228_bits_read; // @[RegisterRouter.scala 65:29]
  Queue Queue ( // @[Decoupled.scala 296:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_read(Queue_io_enq_bits_read),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_extra(Queue_io_enq_bits_extra),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_read(Queue_io_deq_bits_read),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_extra(Queue_io_deq_bits_extra)
  );
  assign auto_register_in_aw_ready = _T_12 & auto_register_in_w_valid; // @[LazyModule.scala 173:31]
  assign auto_register_in_w_ready = _T_12 & auto_register_in_aw_valid; // @[LazyModule.scala 173:31]
  assign auto_register_in_b_valid = _T_228_valid & _T_231; // @[LazyModule.scala 173:31]
  assign auto_register_in_b_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_register_in_ar_ready = Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_register_in_r_valid = _T_228_valid & _T_228_bits_read; // @[LazyModule.scala 173:31]
  assign auto_register_in_r_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_register_in_r_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 173:31]
  assign auto_stream_in_ready = _T_7 ? auto_stream_out_1_ready : _T_3; // @[LazyModule.scala 173:31]
  assign auto_stream_out_1_valid = _T_7 & auto_stream_in_valid; // @[LazyModule.scala 173:49]
  assign auto_stream_out_1_bits_data = auto_stream_in_bits_data; // @[LazyModule.scala 173:49]
  assign auto_stream_out_1_bits_last = auto_stream_in_bits_last; // @[LazyModule.scala 173:49]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_register_in_ar_valid | _T_9; // @[Decoupled.scala 297:22]
  assign Queue_io_enq_bits_read = auto_register_in_ar_valid; // @[Decoupled.scala 298:21]
  assign Queue_io_enq_bits_data = {{31'd0}, _T_227}; // @[Decoupled.scala 298:21]
  assign Queue_io_enq_bits_extra = auto_register_in_ar_valid ? auto_register_in_ar_bits_id : auto_register_in_aw_bits_id; // @[Decoupled.scala 298:21]
  assign Queue_io_deq_ready = _T_228_bits_read ? auto_register_in_r_ready : auto_register_in_b_ready; // @[Decoupled.scala 320:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  sels_0 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  sels_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    sels_0 <= reset | _GEN_19;
    sels_1 <= reset | _GEN_18;
  end
endmodule
module NCOTableStandardMode(
  input  [8:0]  io_phase,
  output [15:0] io_sinOut,
  output [15:0] io_cosOut
);
  wire [1:0] msbs = io_phase[8:7]; // @[NCOTable.scala 123:15]
  wire [6:0] addr = io_phase[6:0]; // @[NCOTable.scala 131:15]
  wire  _T_24 = 2'h0 == msbs; // @[Conditional.scala 37:30]
  wire [6:0] _T_26 = 7'h0 - addr; // @[NCOTable.scala 173:9]
  wire  _T_33 = 2'h1 == msbs; // @[Conditional.scala 37:30]
  wire  _T_42 = 2'h2 == msbs; // @[Conditional.scala 37:30]
  wire  _T_51 = 2'h3 == msbs; // @[Conditional.scala 37:30]
  wire [6:0] _GEN_1 = _T_51 ? addr : 7'h0; // @[Conditional.scala 39:67]
  wire [6:0] _GEN_7 = _T_42 ? _T_26 : _GEN_1; // @[Conditional.scala 39:67]
  wire [6:0] _GEN_15 = _T_33 ? addr : _GEN_7; // @[Conditional.scala 39:67]
  wire [6:0] cosAddr = _T_24 ? _T_26 : _GEN_15; // @[Conditional.scala 40:58]
  wire  _T_27 = cosAddr == 7'h0; // @[NCOTable.scala 199:27]
  wire  _T_28 = addr == 7'h0; // @[NCOTable.scala 199:43]
  wire  _T_29 = _T_27 & _T_28; // @[NCOTable.scala 199:35]
  wire [6:0] _GEN_0 = _T_51 ? _T_26 : 7'h0; // @[Conditional.scala 39:67]
  wire [6:0] _GEN_6 = _T_42 ? addr : _GEN_0; // @[Conditional.scala 39:67]
  wire [6:0] _GEN_14 = _T_33 ? _T_26 : _GEN_6; // @[Conditional.scala 39:67]
  wire [6:0] sinAddr = _T_24 ? addr : _GEN_14; // @[Conditional.scala 40:58]
  wire  _T_36 = sinAddr == 7'h0; // @[NCOTable.scala 209:27]
  wire  _T_38 = _T_36 & _T_28; // @[NCOTable.scala 209:35]
  wire  _GEN_4 = _T_51 & _T_38; // @[Conditional.scala 39:67]
  wire  _GEN_8 = _T_42 | _T_51; // @[Conditional.scala 39:67]
  wire  _GEN_10 = _T_42 & _T_29; // @[Conditional.scala 39:67]
  wire  _GEN_12 = _T_42 ? 1'h0 : _GEN_4; // @[Conditional.scala 39:67]
  wire  _GEN_16 = _T_33 ? 1'h0 : _GEN_8; // @[Conditional.scala 39:67]
  wire  _GEN_17 = _T_33 | _T_42; // @[Conditional.scala 39:67]
  wire  _GEN_18 = _T_33 ? _T_38 : _GEN_12; // @[Conditional.scala 39:67]
  wire  _GEN_20 = _T_33 ? 1'h0 : _GEN_10; // @[Conditional.scala 39:67]
  wire  sinNegative2 = _T_24 ? 1'h0 : _GEN_16; // @[Conditional.scala 40:58]
  wire  cosNegative2 = _T_24 ? 1'h0 : _GEN_17; // @[Conditional.scala 40:58]
  wire  _GEN_26 = _T_24 ? _T_29 : _GEN_20; // @[Conditional.scala 40:58]
  wire  _GEN_28 = _T_24 ? 1'h0 : _GEN_18; // @[Conditional.scala 40:58]
  wire [15:0] _GEN_31 = 7'h1 == sinAddr ? $signed(16'shc9) : $signed(16'sh0); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_32 = 7'h2 == sinAddr ? $signed(16'sh192) : $signed(_GEN_31); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_33 = 7'h3 == sinAddr ? $signed(16'sh25b) : $signed(_GEN_32); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_34 = 7'h4 == sinAddr ? $signed(16'sh324) : $signed(_GEN_33); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_35 = 7'h5 == sinAddr ? $signed(16'sh3ed) : $signed(_GEN_34); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_36 = 7'h6 == sinAddr ? $signed(16'sh4b5) : $signed(_GEN_35); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_37 = 7'h7 == sinAddr ? $signed(16'sh57e) : $signed(_GEN_36); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_38 = 7'h8 == sinAddr ? $signed(16'sh646) : $signed(_GEN_37); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_39 = 7'h9 == sinAddr ? $signed(16'sh70e) : $signed(_GEN_38); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_40 = 7'ha == sinAddr ? $signed(16'sh7d6) : $signed(_GEN_39); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_41 = 7'hb == sinAddr ? $signed(16'sh89d) : $signed(_GEN_40); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_42 = 7'hc == sinAddr ? $signed(16'sh964) : $signed(_GEN_41); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_43 = 7'hd == sinAddr ? $signed(16'sha2b) : $signed(_GEN_42); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_44 = 7'he == sinAddr ? $signed(16'shaf1) : $signed(_GEN_43); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_45 = 7'hf == sinAddr ? $signed(16'shbb7) : $signed(_GEN_44); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_46 = 7'h10 == sinAddr ? $signed(16'shc7c) : $signed(_GEN_45); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_47 = 7'h11 == sinAddr ? $signed(16'shd41) : $signed(_GEN_46); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_48 = 7'h12 == sinAddr ? $signed(16'she06) : $signed(_GEN_47); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_49 = 7'h13 == sinAddr ? $signed(16'sheca) : $signed(_GEN_48); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_50 = 7'h14 == sinAddr ? $signed(16'shf8d) : $signed(_GEN_49); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_51 = 7'h15 == sinAddr ? $signed(16'sh1050) : $signed(_GEN_50); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_52 = 7'h16 == sinAddr ? $signed(16'sh1112) : $signed(_GEN_51); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_53 = 7'h17 == sinAddr ? $signed(16'sh11d3) : $signed(_GEN_52); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_54 = 7'h18 == sinAddr ? $signed(16'sh1294) : $signed(_GEN_53); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_55 = 7'h19 == sinAddr ? $signed(16'sh1354) : $signed(_GEN_54); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_56 = 7'h1a == sinAddr ? $signed(16'sh1413) : $signed(_GEN_55); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_57 = 7'h1b == sinAddr ? $signed(16'sh14d2) : $signed(_GEN_56); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_58 = 7'h1c == sinAddr ? $signed(16'sh1590) : $signed(_GEN_57); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_59 = 7'h1d == sinAddr ? $signed(16'sh164c) : $signed(_GEN_58); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_60 = 7'h1e == sinAddr ? $signed(16'sh1709) : $signed(_GEN_59); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_61 = 7'h1f == sinAddr ? $signed(16'sh17c4) : $signed(_GEN_60); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_62 = 7'h20 == sinAddr ? $signed(16'sh187e) : $signed(_GEN_61); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_63 = 7'h21 == sinAddr ? $signed(16'sh1937) : $signed(_GEN_62); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_64 = 7'h22 == sinAddr ? $signed(16'sh19ef) : $signed(_GEN_63); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_65 = 7'h23 == sinAddr ? $signed(16'sh1aa7) : $signed(_GEN_64); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_66 = 7'h24 == sinAddr ? $signed(16'sh1b5d) : $signed(_GEN_65); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_67 = 7'h25 == sinAddr ? $signed(16'sh1c12) : $signed(_GEN_66); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_68 = 7'h26 == sinAddr ? $signed(16'sh1cc6) : $signed(_GEN_67); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_69 = 7'h27 == sinAddr ? $signed(16'sh1d79) : $signed(_GEN_68); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_70 = 7'h28 == sinAddr ? $signed(16'sh1e2b) : $signed(_GEN_69); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_71 = 7'h29 == sinAddr ? $signed(16'sh1edc) : $signed(_GEN_70); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_72 = 7'h2a == sinAddr ? $signed(16'sh1f8c) : $signed(_GEN_71); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_73 = 7'h2b == sinAddr ? $signed(16'sh203a) : $signed(_GEN_72); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_74 = 7'h2c == sinAddr ? $signed(16'sh20e7) : $signed(_GEN_73); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_75 = 7'h2d == sinAddr ? $signed(16'sh2193) : $signed(_GEN_74); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_76 = 7'h2e == sinAddr ? $signed(16'sh223d) : $signed(_GEN_75); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_77 = 7'h2f == sinAddr ? $signed(16'sh22e7) : $signed(_GEN_76); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_78 = 7'h30 == sinAddr ? $signed(16'sh238e) : $signed(_GEN_77); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_79 = 7'h31 == sinAddr ? $signed(16'sh2435) : $signed(_GEN_78); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_80 = 7'h32 == sinAddr ? $signed(16'sh24da) : $signed(_GEN_79); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_81 = 7'h33 == sinAddr ? $signed(16'sh257e) : $signed(_GEN_80); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_82 = 7'h34 == sinAddr ? $signed(16'sh2620) : $signed(_GEN_81); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_83 = 7'h35 == sinAddr ? $signed(16'sh26c1) : $signed(_GEN_82); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_84 = 7'h36 == sinAddr ? $signed(16'sh2760) : $signed(_GEN_83); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_85 = 7'h37 == sinAddr ? $signed(16'sh27fe) : $signed(_GEN_84); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_86 = 7'h38 == sinAddr ? $signed(16'sh289a) : $signed(_GEN_85); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_87 = 7'h39 == sinAddr ? $signed(16'sh2935) : $signed(_GEN_86); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_88 = 7'h3a == sinAddr ? $signed(16'sh29ce) : $signed(_GEN_87); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_89 = 7'h3b == sinAddr ? $signed(16'sh2a65) : $signed(_GEN_88); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_90 = 7'h3c == sinAddr ? $signed(16'sh2afb) : $signed(_GEN_89); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_91 = 7'h3d == sinAddr ? $signed(16'sh2b8f) : $signed(_GEN_90); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_92 = 7'h3e == sinAddr ? $signed(16'sh2c21) : $signed(_GEN_91); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_93 = 7'h3f == sinAddr ? $signed(16'sh2cb2) : $signed(_GEN_92); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_94 = 7'h40 == sinAddr ? $signed(16'sh2d41) : $signed(_GEN_93); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_95 = 7'h41 == sinAddr ? $signed(16'sh2dcf) : $signed(_GEN_94); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_96 = 7'h42 == sinAddr ? $signed(16'sh2e5a) : $signed(_GEN_95); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_97 = 7'h43 == sinAddr ? $signed(16'sh2ee4) : $signed(_GEN_96); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_98 = 7'h44 == sinAddr ? $signed(16'sh2f6c) : $signed(_GEN_97); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_99 = 7'h45 == sinAddr ? $signed(16'sh2ff2) : $signed(_GEN_98); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_100 = 7'h46 == sinAddr ? $signed(16'sh3076) : $signed(_GEN_99); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_101 = 7'h47 == sinAddr ? $signed(16'sh30f9) : $signed(_GEN_100); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_102 = 7'h48 == sinAddr ? $signed(16'sh3179) : $signed(_GEN_101); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_103 = 7'h49 == sinAddr ? $signed(16'sh31f8) : $signed(_GEN_102); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_104 = 7'h4a == sinAddr ? $signed(16'sh3274) : $signed(_GEN_103); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_105 = 7'h4b == sinAddr ? $signed(16'sh32ef) : $signed(_GEN_104); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_106 = 7'h4c == sinAddr ? $signed(16'sh3368) : $signed(_GEN_105); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_107 = 7'h4d == sinAddr ? $signed(16'sh33df) : $signed(_GEN_106); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_108 = 7'h4e == sinAddr ? $signed(16'sh3453) : $signed(_GEN_107); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_109 = 7'h4f == sinAddr ? $signed(16'sh34c6) : $signed(_GEN_108); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_110 = 7'h50 == sinAddr ? $signed(16'sh3537) : $signed(_GEN_109); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_111 = 7'h51 == sinAddr ? $signed(16'sh35a5) : $signed(_GEN_110); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_112 = 7'h52 == sinAddr ? $signed(16'sh3612) : $signed(_GEN_111); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_113 = 7'h53 == sinAddr ? $signed(16'sh367d) : $signed(_GEN_112); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_114 = 7'h54 == sinAddr ? $signed(16'sh36e5) : $signed(_GEN_113); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_115 = 7'h55 == sinAddr ? $signed(16'sh374b) : $signed(_GEN_114); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_116 = 7'h56 == sinAddr ? $signed(16'sh37b0) : $signed(_GEN_115); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_117 = 7'h57 == sinAddr ? $signed(16'sh3812) : $signed(_GEN_116); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_118 = 7'h58 == sinAddr ? $signed(16'sh3871) : $signed(_GEN_117); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_119 = 7'h59 == sinAddr ? $signed(16'sh38cf) : $signed(_GEN_118); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_120 = 7'h5a == sinAddr ? $signed(16'sh392b) : $signed(_GEN_119); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_121 = 7'h5b == sinAddr ? $signed(16'sh3984) : $signed(_GEN_120); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_122 = 7'h5c == sinAddr ? $signed(16'sh39db) : $signed(_GEN_121); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_123 = 7'h5d == sinAddr ? $signed(16'sh3a30) : $signed(_GEN_122); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_124 = 7'h5e == sinAddr ? $signed(16'sh3a82) : $signed(_GEN_123); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_125 = 7'h5f == sinAddr ? $signed(16'sh3ad3) : $signed(_GEN_124); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_126 = 7'h60 == sinAddr ? $signed(16'sh3b21) : $signed(_GEN_125); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_127 = 7'h61 == sinAddr ? $signed(16'sh3b6d) : $signed(_GEN_126); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_128 = 7'h62 == sinAddr ? $signed(16'sh3bb6) : $signed(_GEN_127); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_129 = 7'h63 == sinAddr ? $signed(16'sh3bfd) : $signed(_GEN_128); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_130 = 7'h64 == sinAddr ? $signed(16'sh3c42) : $signed(_GEN_129); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_131 = 7'h65 == sinAddr ? $signed(16'sh3c85) : $signed(_GEN_130); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_132 = 7'h66 == sinAddr ? $signed(16'sh3cc5) : $signed(_GEN_131); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_133 = 7'h67 == sinAddr ? $signed(16'sh3d03) : $signed(_GEN_132); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_134 = 7'h68 == sinAddr ? $signed(16'sh3d3f) : $signed(_GEN_133); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_135 = 7'h69 == sinAddr ? $signed(16'sh3d78) : $signed(_GEN_134); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_136 = 7'h6a == sinAddr ? $signed(16'sh3daf) : $signed(_GEN_135); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_137 = 7'h6b == sinAddr ? $signed(16'sh3de3) : $signed(_GEN_136); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_138 = 7'h6c == sinAddr ? $signed(16'sh3e15) : $signed(_GEN_137); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_139 = 7'h6d == sinAddr ? $signed(16'sh3e45) : $signed(_GEN_138); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_140 = 7'h6e == sinAddr ? $signed(16'sh3e72) : $signed(_GEN_139); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_141 = 7'h6f == sinAddr ? $signed(16'sh3e9d) : $signed(_GEN_140); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_142 = 7'h70 == sinAddr ? $signed(16'sh3ec5) : $signed(_GEN_141); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_143 = 7'h71 == sinAddr ? $signed(16'sh3eeb) : $signed(_GEN_142); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_144 = 7'h72 == sinAddr ? $signed(16'sh3f0f) : $signed(_GEN_143); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_145 = 7'h73 == sinAddr ? $signed(16'sh3f30) : $signed(_GEN_144); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_146 = 7'h74 == sinAddr ? $signed(16'sh3f4f) : $signed(_GEN_145); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_147 = 7'h75 == sinAddr ? $signed(16'sh3f6b) : $signed(_GEN_146); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_148 = 7'h76 == sinAddr ? $signed(16'sh3f85) : $signed(_GEN_147); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_149 = 7'h77 == sinAddr ? $signed(16'sh3f9c) : $signed(_GEN_148); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_150 = 7'h78 == sinAddr ? $signed(16'sh3fb1) : $signed(_GEN_149); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_151 = 7'h79 == sinAddr ? $signed(16'sh3fc4) : $signed(_GEN_150); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_152 = 7'h7a == sinAddr ? $signed(16'sh3fd4) : $signed(_GEN_151); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_153 = 7'h7b == sinAddr ? $signed(16'sh3fe1) : $signed(_GEN_152); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_154 = 7'h7c == sinAddr ? $signed(16'sh3fec) : $signed(_GEN_153); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_155 = 7'h7d == sinAddr ? $signed(16'sh3ff5) : $signed(_GEN_154); // @[NCOTable.scala 260:64]
  wire [15:0] _GEN_156 = 7'h7e == sinAddr ? $signed(16'sh3ffb) : $signed(_GEN_155); // @[NCOTable.scala 260:64]
  wire [15:0] _T_65 = 7'h7f == sinAddr ? $signed(16'sh3fff) : $signed(_GEN_156); // @[NCOTable.scala 260:64]
  wire [15:0] sinTableOut = _GEN_28 ? $signed(16'sh4000) : $signed(_T_65); // @[NCOTable.scala 260:23]
  wire [15:0] _GEN_159 = 7'h1 == cosAddr ? $signed(16'shc9) : $signed(16'sh0); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_160 = 7'h2 == cosAddr ? $signed(16'sh192) : $signed(_GEN_159); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_161 = 7'h3 == cosAddr ? $signed(16'sh25b) : $signed(_GEN_160); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_162 = 7'h4 == cosAddr ? $signed(16'sh324) : $signed(_GEN_161); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_163 = 7'h5 == cosAddr ? $signed(16'sh3ed) : $signed(_GEN_162); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_164 = 7'h6 == cosAddr ? $signed(16'sh4b5) : $signed(_GEN_163); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_165 = 7'h7 == cosAddr ? $signed(16'sh57e) : $signed(_GEN_164); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_166 = 7'h8 == cosAddr ? $signed(16'sh646) : $signed(_GEN_165); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_167 = 7'h9 == cosAddr ? $signed(16'sh70e) : $signed(_GEN_166); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_168 = 7'ha == cosAddr ? $signed(16'sh7d6) : $signed(_GEN_167); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_169 = 7'hb == cosAddr ? $signed(16'sh89d) : $signed(_GEN_168); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_170 = 7'hc == cosAddr ? $signed(16'sh964) : $signed(_GEN_169); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_171 = 7'hd == cosAddr ? $signed(16'sha2b) : $signed(_GEN_170); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_172 = 7'he == cosAddr ? $signed(16'shaf1) : $signed(_GEN_171); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_173 = 7'hf == cosAddr ? $signed(16'shbb7) : $signed(_GEN_172); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_174 = 7'h10 == cosAddr ? $signed(16'shc7c) : $signed(_GEN_173); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_175 = 7'h11 == cosAddr ? $signed(16'shd41) : $signed(_GEN_174); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_176 = 7'h12 == cosAddr ? $signed(16'she06) : $signed(_GEN_175); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_177 = 7'h13 == cosAddr ? $signed(16'sheca) : $signed(_GEN_176); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_178 = 7'h14 == cosAddr ? $signed(16'shf8d) : $signed(_GEN_177); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_179 = 7'h15 == cosAddr ? $signed(16'sh1050) : $signed(_GEN_178); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_180 = 7'h16 == cosAddr ? $signed(16'sh1112) : $signed(_GEN_179); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_181 = 7'h17 == cosAddr ? $signed(16'sh11d3) : $signed(_GEN_180); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_182 = 7'h18 == cosAddr ? $signed(16'sh1294) : $signed(_GEN_181); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_183 = 7'h19 == cosAddr ? $signed(16'sh1354) : $signed(_GEN_182); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_184 = 7'h1a == cosAddr ? $signed(16'sh1413) : $signed(_GEN_183); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_185 = 7'h1b == cosAddr ? $signed(16'sh14d2) : $signed(_GEN_184); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_186 = 7'h1c == cosAddr ? $signed(16'sh1590) : $signed(_GEN_185); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_187 = 7'h1d == cosAddr ? $signed(16'sh164c) : $signed(_GEN_186); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_188 = 7'h1e == cosAddr ? $signed(16'sh1709) : $signed(_GEN_187); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_189 = 7'h1f == cosAddr ? $signed(16'sh17c4) : $signed(_GEN_188); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_190 = 7'h20 == cosAddr ? $signed(16'sh187e) : $signed(_GEN_189); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_191 = 7'h21 == cosAddr ? $signed(16'sh1937) : $signed(_GEN_190); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_192 = 7'h22 == cosAddr ? $signed(16'sh19ef) : $signed(_GEN_191); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_193 = 7'h23 == cosAddr ? $signed(16'sh1aa7) : $signed(_GEN_192); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_194 = 7'h24 == cosAddr ? $signed(16'sh1b5d) : $signed(_GEN_193); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_195 = 7'h25 == cosAddr ? $signed(16'sh1c12) : $signed(_GEN_194); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_196 = 7'h26 == cosAddr ? $signed(16'sh1cc6) : $signed(_GEN_195); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_197 = 7'h27 == cosAddr ? $signed(16'sh1d79) : $signed(_GEN_196); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_198 = 7'h28 == cosAddr ? $signed(16'sh1e2b) : $signed(_GEN_197); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_199 = 7'h29 == cosAddr ? $signed(16'sh1edc) : $signed(_GEN_198); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_200 = 7'h2a == cosAddr ? $signed(16'sh1f8c) : $signed(_GEN_199); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_201 = 7'h2b == cosAddr ? $signed(16'sh203a) : $signed(_GEN_200); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_202 = 7'h2c == cosAddr ? $signed(16'sh20e7) : $signed(_GEN_201); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_203 = 7'h2d == cosAddr ? $signed(16'sh2193) : $signed(_GEN_202); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_204 = 7'h2e == cosAddr ? $signed(16'sh223d) : $signed(_GEN_203); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_205 = 7'h2f == cosAddr ? $signed(16'sh22e7) : $signed(_GEN_204); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_206 = 7'h30 == cosAddr ? $signed(16'sh238e) : $signed(_GEN_205); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_207 = 7'h31 == cosAddr ? $signed(16'sh2435) : $signed(_GEN_206); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_208 = 7'h32 == cosAddr ? $signed(16'sh24da) : $signed(_GEN_207); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_209 = 7'h33 == cosAddr ? $signed(16'sh257e) : $signed(_GEN_208); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_210 = 7'h34 == cosAddr ? $signed(16'sh2620) : $signed(_GEN_209); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_211 = 7'h35 == cosAddr ? $signed(16'sh26c1) : $signed(_GEN_210); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_212 = 7'h36 == cosAddr ? $signed(16'sh2760) : $signed(_GEN_211); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_213 = 7'h37 == cosAddr ? $signed(16'sh27fe) : $signed(_GEN_212); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_214 = 7'h38 == cosAddr ? $signed(16'sh289a) : $signed(_GEN_213); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_215 = 7'h39 == cosAddr ? $signed(16'sh2935) : $signed(_GEN_214); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_216 = 7'h3a == cosAddr ? $signed(16'sh29ce) : $signed(_GEN_215); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_217 = 7'h3b == cosAddr ? $signed(16'sh2a65) : $signed(_GEN_216); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_218 = 7'h3c == cosAddr ? $signed(16'sh2afb) : $signed(_GEN_217); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_219 = 7'h3d == cosAddr ? $signed(16'sh2b8f) : $signed(_GEN_218); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_220 = 7'h3e == cosAddr ? $signed(16'sh2c21) : $signed(_GEN_219); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_221 = 7'h3f == cosAddr ? $signed(16'sh2cb2) : $signed(_GEN_220); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_222 = 7'h40 == cosAddr ? $signed(16'sh2d41) : $signed(_GEN_221); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_223 = 7'h41 == cosAddr ? $signed(16'sh2dcf) : $signed(_GEN_222); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_224 = 7'h42 == cosAddr ? $signed(16'sh2e5a) : $signed(_GEN_223); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_225 = 7'h43 == cosAddr ? $signed(16'sh2ee4) : $signed(_GEN_224); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_226 = 7'h44 == cosAddr ? $signed(16'sh2f6c) : $signed(_GEN_225); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_227 = 7'h45 == cosAddr ? $signed(16'sh2ff2) : $signed(_GEN_226); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_228 = 7'h46 == cosAddr ? $signed(16'sh3076) : $signed(_GEN_227); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_229 = 7'h47 == cosAddr ? $signed(16'sh30f9) : $signed(_GEN_228); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_230 = 7'h48 == cosAddr ? $signed(16'sh3179) : $signed(_GEN_229); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_231 = 7'h49 == cosAddr ? $signed(16'sh31f8) : $signed(_GEN_230); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_232 = 7'h4a == cosAddr ? $signed(16'sh3274) : $signed(_GEN_231); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_233 = 7'h4b == cosAddr ? $signed(16'sh32ef) : $signed(_GEN_232); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_234 = 7'h4c == cosAddr ? $signed(16'sh3368) : $signed(_GEN_233); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_235 = 7'h4d == cosAddr ? $signed(16'sh33df) : $signed(_GEN_234); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_236 = 7'h4e == cosAddr ? $signed(16'sh3453) : $signed(_GEN_235); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_237 = 7'h4f == cosAddr ? $signed(16'sh34c6) : $signed(_GEN_236); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_238 = 7'h50 == cosAddr ? $signed(16'sh3537) : $signed(_GEN_237); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_239 = 7'h51 == cosAddr ? $signed(16'sh35a5) : $signed(_GEN_238); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_240 = 7'h52 == cosAddr ? $signed(16'sh3612) : $signed(_GEN_239); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_241 = 7'h53 == cosAddr ? $signed(16'sh367d) : $signed(_GEN_240); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_242 = 7'h54 == cosAddr ? $signed(16'sh36e5) : $signed(_GEN_241); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_243 = 7'h55 == cosAddr ? $signed(16'sh374b) : $signed(_GEN_242); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_244 = 7'h56 == cosAddr ? $signed(16'sh37b0) : $signed(_GEN_243); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_245 = 7'h57 == cosAddr ? $signed(16'sh3812) : $signed(_GEN_244); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_246 = 7'h58 == cosAddr ? $signed(16'sh3871) : $signed(_GEN_245); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_247 = 7'h59 == cosAddr ? $signed(16'sh38cf) : $signed(_GEN_246); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_248 = 7'h5a == cosAddr ? $signed(16'sh392b) : $signed(_GEN_247); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_249 = 7'h5b == cosAddr ? $signed(16'sh3984) : $signed(_GEN_248); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_250 = 7'h5c == cosAddr ? $signed(16'sh39db) : $signed(_GEN_249); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_251 = 7'h5d == cosAddr ? $signed(16'sh3a30) : $signed(_GEN_250); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_252 = 7'h5e == cosAddr ? $signed(16'sh3a82) : $signed(_GEN_251); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_253 = 7'h5f == cosAddr ? $signed(16'sh3ad3) : $signed(_GEN_252); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_254 = 7'h60 == cosAddr ? $signed(16'sh3b21) : $signed(_GEN_253); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_255 = 7'h61 == cosAddr ? $signed(16'sh3b6d) : $signed(_GEN_254); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_256 = 7'h62 == cosAddr ? $signed(16'sh3bb6) : $signed(_GEN_255); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_257 = 7'h63 == cosAddr ? $signed(16'sh3bfd) : $signed(_GEN_256); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_258 = 7'h64 == cosAddr ? $signed(16'sh3c42) : $signed(_GEN_257); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_259 = 7'h65 == cosAddr ? $signed(16'sh3c85) : $signed(_GEN_258); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_260 = 7'h66 == cosAddr ? $signed(16'sh3cc5) : $signed(_GEN_259); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_261 = 7'h67 == cosAddr ? $signed(16'sh3d03) : $signed(_GEN_260); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_262 = 7'h68 == cosAddr ? $signed(16'sh3d3f) : $signed(_GEN_261); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_263 = 7'h69 == cosAddr ? $signed(16'sh3d78) : $signed(_GEN_262); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_264 = 7'h6a == cosAddr ? $signed(16'sh3daf) : $signed(_GEN_263); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_265 = 7'h6b == cosAddr ? $signed(16'sh3de3) : $signed(_GEN_264); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_266 = 7'h6c == cosAddr ? $signed(16'sh3e15) : $signed(_GEN_265); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_267 = 7'h6d == cosAddr ? $signed(16'sh3e45) : $signed(_GEN_266); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_268 = 7'h6e == cosAddr ? $signed(16'sh3e72) : $signed(_GEN_267); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_269 = 7'h6f == cosAddr ? $signed(16'sh3e9d) : $signed(_GEN_268); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_270 = 7'h70 == cosAddr ? $signed(16'sh3ec5) : $signed(_GEN_269); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_271 = 7'h71 == cosAddr ? $signed(16'sh3eeb) : $signed(_GEN_270); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_272 = 7'h72 == cosAddr ? $signed(16'sh3f0f) : $signed(_GEN_271); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_273 = 7'h73 == cosAddr ? $signed(16'sh3f30) : $signed(_GEN_272); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_274 = 7'h74 == cosAddr ? $signed(16'sh3f4f) : $signed(_GEN_273); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_275 = 7'h75 == cosAddr ? $signed(16'sh3f6b) : $signed(_GEN_274); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_276 = 7'h76 == cosAddr ? $signed(16'sh3f85) : $signed(_GEN_275); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_277 = 7'h77 == cosAddr ? $signed(16'sh3f9c) : $signed(_GEN_276); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_278 = 7'h78 == cosAddr ? $signed(16'sh3fb1) : $signed(_GEN_277); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_279 = 7'h79 == cosAddr ? $signed(16'sh3fc4) : $signed(_GEN_278); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_280 = 7'h7a == cosAddr ? $signed(16'sh3fd4) : $signed(_GEN_279); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_281 = 7'h7b == cosAddr ? $signed(16'sh3fe1) : $signed(_GEN_280); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_282 = 7'h7c == cosAddr ? $signed(16'sh3fec) : $signed(_GEN_281); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_283 = 7'h7d == cosAddr ? $signed(16'sh3ff5) : $signed(_GEN_282); // @[NCOTable.scala 261:64]
  wire [15:0] _GEN_284 = 7'h7e == cosAddr ? $signed(16'sh3ffb) : $signed(_GEN_283); // @[NCOTable.scala 261:64]
  wire [15:0] _T_71 = 7'h7f == cosAddr ? $signed(16'sh3fff) : $signed(_GEN_284); // @[NCOTable.scala 261:64]
  wire [15:0] cosTableOut = _GEN_26 ? $signed(16'sh4000) : $signed(_T_71); // @[NCOTable.scala 261:23]
  wire [15:0] _T_75 = 16'sh0 - $signed(sinTableOut); // @[FixedPointTypeClass.scala 39:43]
  wire [15:0] _T_78 = 16'sh0 - $signed(cosTableOut); // @[FixedPointTypeClass.scala 39:43]
  assign io_sinOut = sinNegative2 ? $signed(_T_75) : $signed(sinTableOut); // @[NCOTable.scala 314:13]
  assign io_cosOut = cosNegative2 ? $signed(_T_78) : $signed(cosTableOut); // @[NCOTable.scala 315:13]
endmodule
module NCOTable(
  input  [8:0]  io_phase,
  output [15:0] io_sinOut,
  output [15:0] io_cosOut
);
  wire [8:0] tableNCO_io_phase; // @[NCOTable.scala 473:13]
  wire [15:0] tableNCO_io_sinOut; // @[NCOTable.scala 473:13]
  wire [15:0] tableNCO_io_cosOut; // @[NCOTable.scala 473:13]
  NCOTableStandardMode tableNCO ( // @[NCOTable.scala 473:13]
    .io_phase(tableNCO_io_phase),
    .io_sinOut(tableNCO_io_sinOut),
    .io_cosOut(tableNCO_io_cosOut)
  );
  assign io_sinOut = tableNCO_io_sinOut; // @[NCOTable.scala 478:13]
  assign io_cosOut = tableNCO_io_cosOut; // @[NCOTable.scala 479:13]
  assign tableNCO_io_phase = io_phase; // @[NCOTable.scala 477:21]
endmodule
module Queue_6(
  input   clock,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input   io_enq_bits,
  input   io_deq_ready,
  output  io_deq_valid,
  output  io_deq_bits
);
  reg  _T [0:1]; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_0;
  wire  _T__T_18_data; // @[Decoupled.scala 218:24]
  wire  _T__T_18_addr; // @[Decoupled.scala 218:24]
  wire  _T__T_10_data; // @[Decoupled.scala 218:24]
  wire  _T__T_10_addr; // @[Decoupled.scala 218:24]
  wire  _T__T_10_mask; // @[Decoupled.scala 218:24]
  wire  _T__T_10_en; // @[Decoupled.scala 218:24]
  reg  value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_1;
  reg  value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_2;
  reg  _T_1; // @[Decoupled.scala 221:35]
  reg [31:0] _RAND_3;
  wire  _T_2 = value == value_1; // @[Decoupled.scala 223:41]
  wire  _T_3 = ~_T_1; // @[Decoupled.scala 224:36]
  wire  _T_4 = _T_2 & _T_3; // @[Decoupled.scala 224:33]
  wire  _T_5 = _T_2 & _T_1; // @[Decoupled.scala 225:32]
  wire  _T_6 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  _T_8 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire  _T_12 = value + 1'h1; // @[Counter.scala 39:22]
  wire  _T_14 = value_1 + 1'h1; // @[Counter.scala 39:22]
  wire  _T_15 = _T_6 != _T_8; // @[Decoupled.scala 236:16]
  wire  _T_17 = ~_T_5; // @[Decoupled.scala 241:19]
  assign _T__T_18_addr = value_1;
  assign _T__T_18_data = _T[_T__T_18_addr]; // @[Decoupled.scala 218:24]
  assign _T__T_10_data = io_enq_bits;
  assign _T__T_10_addr = value;
  assign _T__T_10_mask = 1'h1;
  assign _T__T_10_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = io_deq_ready | _T_17; // @[Decoupled.scala 241:16 Decoupled.scala 254:40]
  assign io_deq_valid = ~_T_4; // @[Decoupled.scala 240:16]
  assign io_deq_bits = _T__T_18_data; // @[Decoupled.scala 242:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T[initvar] = _RAND_0[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  value = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  value_1 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_1 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T__T_10_en & _T__T_10_mask) begin
      _T[_T__T_10_addr] <= _T__T_10_data; // @[Decoupled.scala 218:24]
    end
    if (reset) begin
      value <= 1'h0;
    end else if (_T_6) begin
      value <= _T_12;
    end
    if (reset) begin
      value_1 <= 1'h0;
    end else if (_T_8) begin
      value_1 <= _T_14;
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else if (_T_15) begin
      _T_1 <= _T_6;
    end
  end
endmodule
module AXI4NCOLazyModuleBlock(
  input         clock,
  input         reset,
  input         auto_stream_out_ready,
  output        auto_stream_out_valid,
  output [31:0] auto_stream_out_bits_data,
  output        auto_stream_out_bits_last,
  output        auto_freq_in_ready,
  input         auto_freq_in_valid,
  input  [31:0] auto_freq_in_bits_data,
  input         auto_freq_in_bits_last
);
  wire [8:0] phaseConverter_io_phase; // @[NCOLazyModuleBlock.scala 35:32]
  wire [15:0] phaseConverter_io_sinOut; // @[NCOLazyModuleBlock.scala 35:32]
  wire [15:0] phaseConverter_io_cosOut; // @[NCOLazyModuleBlock.scala 35:32]
  wire  Queue_clock; // @[Skid.scala 21:23]
  wire  Queue_reset; // @[Skid.scala 21:23]
  wire  Queue_io_enq_ready; // @[Skid.scala 21:23]
  wire  Queue_io_enq_valid; // @[Skid.scala 21:23]
  wire  Queue_io_enq_bits; // @[Skid.scala 21:23]
  wire  Queue_io_deq_ready; // @[Skid.scala 21:23]
  wire  Queue_io_deq_valid; // @[Skid.scala 21:23]
  wire  Queue_io_deq_bits; // @[Skid.scala 21:23]
  reg [8:0] phaseCounter; // @[NCOLazyModuleBlock.scala 36:33]
  reg [31:0] _RAND_0;
  reg [1:0] _T_35; // @[NCOLazyModuleBlock.scala 213:33]
  reg [31:0] _RAND_1;
  wire  _T_52 = _T_35 < 2'h2; // @[NCOLazyModuleBlock.scala 223:48]
  wire  _T_53 = _T_35 == 2'h2; // @[NCOLazyModuleBlock.scala 223:78]
  wire  _T_54 = _T_53 & auto_stream_out_ready; // @[NCOLazyModuleBlock.scala 223:92]
  wire  _T_55 = _T_52 | _T_54; // @[NCOLazyModuleBlock.scala 223:61]
  wire  _T_5 = _T_55 & auto_freq_in_valid; // @[Decoupled.scala 40:37]
  wire [31:0] _GEN_15 = {{23'd0}, phaseCounter}; // @[NCOLazyModuleBlock.scala 190:40]
  wire [31:0] _T_7 = _GEN_15 + auto_freq_in_bits_data; // @[NCOLazyModuleBlock.scala 190:40]
  wire [31:0] _GEN_0 = _T_5 ? _T_7 : {{23'd0}, phaseCounter}; // @[NCOLazyModuleBlock.scala 189:40]
  wire [16:0] _T_8 = {{8'd0}, phaseCounter}; // @[NCOLazyModuleBlock.scala 199:47]
  reg  queueCounter; // @[Skid.scala 22:31]
  reg [31:0] _RAND_2;
  wire  _T_26 = queueCounter < 1'h1; // @[Skid.scala 29:31]
  wire  _T_28 = queueCounter & auto_stream_out_ready; // @[Skid.scala 29:75]
  wire  _T_29 = _T_26 | _T_28; // @[Skid.scala 29:44]
  wire  _T_14 = _T_29 & auto_freq_in_valid; // @[Decoupled.scala 40:37]
  wire [1:0] _T_15 = queueCounter + _T_14; // @[Skid.scala 23:34]
  wire  _T_11_valid = Queue_io_deq_valid; // @[NCOLazyModuleBlock.scala 202:29 Skid.scala 31:15]
  wire  _T_16 = auto_stream_out_ready & _T_11_valid; // @[Decoupled.scala 40:37]
  wire [1:0] _GEN_16 = {{1'd0}, _T_16}; // @[Skid.scala 23:47]
  wire [2:0] _T_17 = _T_15 - _GEN_16; // @[Skid.scala 23:47]
  reg  _T_20; // @[Reg.scala 27:20]
  reg [31:0] _RAND_3;
  wire  _T_21 = ~Queue_io_enq_valid; // @[Skid.scala 26:12]
  wire  _T_22 = _T_21 | Queue_io_enq_ready; // @[Skid.scala 26:32]
  wire  _T_24 = _T_22 | reset; // @[Skid.scala 26:11]
  wire  _T_25 = ~_T_24; // @[Skid.scala 26:11]
  reg  ioout_bits_last; // @[NCOLazyModuleBlock.scala 207:28]
  reg [31:0] _RAND_4;
  reg  _T_31; // @[NCOLazyModuleBlock.scala 208:30]
  reg [31:0] _RAND_5;
  wire  _T_11_bits = Queue_io_deq_bits; // @[NCOLazyModuleBlock.scala 202:29 Skid.scala 32:14]
  wire  _GEN_2 = _T_11_bits | _T_31; // @[NCOLazyModuleBlock.scala 209:30]
  wire  _T_32 = ~_T_31; // @[NCOLazyModuleBlock.scala 210:32]
  wire  _T_33 = _T_11_bits & _T_32; // @[NCOLazyModuleBlock.scala 210:29]
  wire  _T_57 = _T_35 == 2'h1; // @[NCOLazyModuleBlock.scala 224:65]
  reg [1:0] _T_46; // @[NCOLazyModuleBlock.scala 218:64]
  reg [31:0] _RAND_6;
  wire  _T_47 = _T_35 != _T_46; // @[NCOLazyModuleBlock.scala 218:53]
  reg [1:0] _T_48; // @[NCOLazyModuleBlock.scala 218:87]
  reg [31:0] _RAND_7;
  reg [1:0] _T_41; // @[NCOLazyModuleBlock.scala 215:42]
  reg [31:0] _RAND_8;
  wire [1:0] _T_49 = _T_47 ? _T_48 : _T_41; // @[NCOLazyModuleBlock.scala 218:39]
  wire  _T_58 = _T_49 == 2'h2; // @[NCOLazyModuleBlock.scala 224:104]
  wire  _T_59 = _T_57 & _T_58; // @[NCOLazyModuleBlock.scala 224:74]
  wire  _T_60 = _T_53 | _T_59; // @[NCOLazyModuleBlock.scala 224:47]
  wire  ioout_valid = _T_60 & auto_stream_out_ready; // @[NCOLazyModuleBlock.scala 224:115]
  wire [1:0] _GEN_17 = {{1'd0}, _T_5}; // @[NCOLazyModuleBlock.scala 214:36]
  wire [2:0] _T_37 = _T_35 + _GEN_17; // @[NCOLazyModuleBlock.scala 214:36]
  wire  _T_38 = auto_stream_out_ready & ioout_valid; // @[Decoupled.scala 40:37]
  wire [2:0] _GEN_18 = {{2'd0}, _T_38}; // @[NCOLazyModuleBlock.scala 214:64]
  wire [3:0] _T_39 = _T_37 - _GEN_18; // @[NCOLazyModuleBlock.scala 214:64]
  reg [1:0] _T_42; // @[NCOLazyModuleBlock.scala 216:37]
  reg [31:0] _RAND_9;
  wire  _T_43 = _T_35 != _T_42; // @[NCOLazyModuleBlock.scala 216:26]
  reg [1:0] _T_44; // @[NCOLazyModuleBlock.scala 216:86]
  reg [31:0] _RAND_10;
  reg  _T_50; // @[NCOLazyModuleBlock.scala 220:27]
  reg [31:0] _RAND_11;
  reg [15:0] _T_64; // @[NCOLazyModuleBlock.scala 226:36]
  reg [31:0] _RAND_12;
  reg [15:0] _T_67; // @[NCOLazyModuleBlock.scala 227:36]
  reg [31:0] _RAND_13;
  reg [15:0] _T_70; // @[NCOLazyModuleBlock.scala 229:37]
  reg [31:0] _RAND_14;
  reg [15:0] _T_73; // @[NCOLazyModuleBlock.scala 230:37]
  reg [31:0] _RAND_15;
  wire  _T_76 = _T_5 & _T_50; // @[NCOLazyModuleBlock.scala 258:39]
  wire [31:0] _T_79 = {_T_67,_T_64}; // @[Cat.scala 29:58]
  wire  _T_81 = ~_T_50; // @[NCOLazyModuleBlock.scala 260:48]
  wire  _T_82 = _T_5 & _T_81; // @[NCOLazyModuleBlock.scala 260:45]
  wire [31:0] _T_85 = {_T_73,_T_70}; // @[Cat.scala 29:58]
  wire  _T_87 = ~_T_5; // @[NCOLazyModuleBlock.scala 262:20]
  wire  _T_88 = _T_87 & _T_50; // @[NCOLazyModuleBlock.scala 262:46]
  wire [31:0] _GEN_11 = _T_88 ? _T_79 : _T_85; // @[NCOLazyModuleBlock.scala 262:56]
  wire [31:0] _GEN_12 = _T_82 ? _T_85 : _GEN_11; // @[NCOLazyModuleBlock.scala 260:56]
  wire [31:0] _GEN_13 = _T_76 ? _T_79 : _GEN_12; // @[NCOLazyModuleBlock.scala 258:49]
  NCOTable phaseConverter ( // @[NCOLazyModuleBlock.scala 35:32]
    .io_phase(phaseConverter_io_phase),
    .io_sinOut(phaseConverter_io_sinOut),
    .io_cosOut(phaseConverter_io_cosOut)
  );
  Queue_6 Queue ( // @[Skid.scala 21:23]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits(Queue_io_enq_bits),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits(Queue_io_deq_bits)
  );
  assign auto_stream_out_valid = _T_60 & auto_stream_out_ready; // @[LazyModule.scala 173:49]
  assign auto_stream_out_bits_data = _T_53 ? _GEN_13 : _T_79; // @[LazyModule.scala 173:49]
  assign auto_stream_out_bits_last = ioout_bits_last; // @[LazyModule.scala 173:49]
  assign auto_freq_in_ready = _T_52 | _T_54; // @[LazyModule.scala 173:31]
  assign phaseConverter_io_phase = _T_8[8:0]; // @[NCOLazyModuleBlock.scala 199:31]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = _T_20; // @[Skid.scala 25:24]
  assign Queue_io_enq_bits = auto_freq_in_bits_last & _T_5; // @[NCOLazyModuleBlock.scala 206:41]
  assign Queue_io_deq_ready = auto_stream_out_ready; // @[Skid.scala 30:24]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  phaseCounter = _RAND_0[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_35 = _RAND_1[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  queueCounter = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_20 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  ioout_bits_last = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_31 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_46 = _RAND_6[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_48 = _RAND_7[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_41 = _RAND_8[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_42 = _RAND_9[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_44 = _RAND_10[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_50 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_64 = _RAND_12[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_67 = _RAND_13[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_70 = _RAND_14[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_73 = _RAND_15[15:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      phaseCounter <= 9'h0;
    end else begin
      phaseCounter <= _GEN_0[8:0];
    end
    if (reset) begin
      _T_35 <= 2'h0;
    end else begin
      _T_35 <= _T_39[1:0];
    end
    if (reset) begin
      queueCounter <= 1'h0;
    end else begin
      queueCounter <= _T_17[0];
    end
    if (reset) begin
      _T_20 <= 1'h0;
    end else begin
      _T_20 <= _T_14;
    end
    if (reset) begin
      ioout_bits_last <= 1'h0;
    end else begin
      ioout_bits_last <= _T_33;
    end
    if (reset) begin
      _T_31 <= 1'h0;
    end else begin
      _T_31 <= _GEN_2;
    end
    _T_46 <= _T_35;
    _T_48 <= _T_35;
    if (reset) begin
      _T_41 <= 2'h0;
    end else if (_T_43) begin
      _T_41 <= _T_44;
    end
    _T_42 <= _T_35;
    _T_44 <= _T_35;
    if (reset) begin
      _T_50 <= 1'h0;
    end else begin
      _T_50 <= _T_5;
    end
    if (reset) begin
      _T_64 <= 16'sh0;
    end else if (_T_50) begin
      _T_64 <= phaseConverter_io_sinOut;
    end
    if (reset) begin
      _T_67 <= 16'sh0;
    end else if (_T_50) begin
      _T_67 <= phaseConverter_io_cosOut;
    end
    if (reset) begin
      _T_70 <= 16'sh0;
    end else if (_T_50) begin
      _T_70 <= _T_64;
    end
    if (reset) begin
      _T_73 <= 16'sh0;
    end else if (_T_50) begin
      _T_73 <= _T_67;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_25) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Skid.scala:26 assert(!queue.io.enq.valid || queue.io.enq.ready) // we control in.ready such that the queue can't fill up!\n"); // @[Skid.scala 26:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_25) begin
          $fatal; // @[Skid.scala 26:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module AXI4Splitter_2(
  input         clock,
  input         reset,
  output        auto_mem_in_aw_ready,
  input         auto_mem_in_aw_valid,
  input         auto_mem_in_aw_bits_id,
  input  [29:0] auto_mem_in_aw_bits_addr,
  output        auto_mem_in_w_ready,
  input         auto_mem_in_w_valid,
  input  [31:0] auto_mem_in_w_bits_data,
  input  [3:0]  auto_mem_in_w_bits_strb,
  input         auto_mem_in_b_ready,
  output        auto_mem_in_b_valid,
  output        auto_mem_in_b_bits_id,
  output        auto_mem_in_ar_ready,
  input         auto_mem_in_ar_valid,
  input         auto_mem_in_ar_bits_id,
  input  [29:0] auto_mem_in_ar_bits_addr,
  input  [2:0]  auto_mem_in_ar_bits_size,
  input         auto_mem_in_r_ready,
  output        auto_mem_in_r_valid,
  output        auto_mem_in_r_bits_id,
  output [31:0] auto_mem_in_r_bits_data,
  output        auto_stream_in_ready,
  input         auto_stream_in_valid,
  input  [31:0] auto_stream_in_bits_data,
  input         auto_stream_in_bits_last,
  input         auto_stream_out_1_ready,
  output        auto_stream_out_1_valid,
  output [31:0] auto_stream_out_1_bits_data,
  output        auto_stream_out_1_bits_last,
  input         auto_stream_out_0_ready,
  output        auto_stream_out_0_valid,
  output [31:0] auto_stream_out_0_bits_data,
  output        auto_stream_out_0_bits_last
);
  wire  Queue_clock; // @[Decoupled.scala 296:21]
  wire  Queue_reset; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_bits_read; // @[Decoupled.scala 296:21]
  wire [31:0] Queue_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_bits_extra; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_bits_read; // @[Decoupled.scala 296:21]
  wire [31:0] Queue_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_bits_extra; // @[Decoupled.scala 296:21]
  reg [31:0] ctrlReg; // @[Splitter.scala 27:26]
  reg [31:0] _RAND_0;
  reg [31:0] maskReg; // @[Splitter.scala 28:26]
  reg [31:0] _RAND_1;
  wire  _T_4 = auto_mem_in_aw_valid & auto_mem_in_w_valid; // @[RegisterRouter.scala 40:39]
  wire  _T_5 = auto_mem_in_ar_valid | _T_4; // @[RegisterRouter.scala 40:26]
  wire  _T_6 = ~auto_mem_in_ar_valid; // @[RegisterRouter.scala 42:29]
  wire  _T_49_ready = Queue_io_enq_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 299:17]
  wire [29:0] _T_13 = auto_mem_in_ar_valid ? auto_mem_in_ar_bits_addr : auto_mem_in_aw_bits_addr; // @[RegisterRouter.scala 48:19]
  wire [1:0] _T_53 = _T_13[3:2] & 2'h2; // @[RegisterRouter.scala 59:16]
  wire  _T_55 = _T_53 == 2'h0; // @[RegisterRouter.scala 59:16]
  wire  _T_7 = _T_49_ready & _T_6; // @[RegisterRouter.scala 42:26]
  wire [1:0] _T_16 = 2'h1 << auto_mem_in_ar_bits_size[0]; // @[OneHot.scala 65:12]
  wire [1:0] _T_18 = _T_16 | 2'h1; // @[Misc.scala 200:81]
  wire  _T_19 = auto_mem_in_ar_bits_size >= 3'h2; // @[Misc.scala 204:21]
  wire  _T_22 = ~auto_mem_in_ar_bits_addr[1]; // @[Misc.scala 209:20]
  wire  _T_24 = _T_18[1] & _T_22; // @[Misc.scala 213:38]
  wire  _T_25 = _T_19 | _T_24; // @[Misc.scala 213:29]
  wire  _T_27 = _T_18[1] & auto_mem_in_ar_bits_addr[1]; // @[Misc.scala 213:38]
  wire  _T_28 = _T_19 | _T_27; // @[Misc.scala 213:29]
  wire  _T_31 = ~auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 209:20]
  wire  _T_32 = _T_22 & _T_31; // @[Misc.scala 212:27]
  wire  _T_33 = _T_18[0] & _T_32; // @[Misc.scala 213:38]
  wire  _T_34 = _T_25 | _T_33; // @[Misc.scala 213:29]
  wire  _T_35 = _T_22 & auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  wire  _T_36 = _T_18[0] & _T_35; // @[Misc.scala 213:38]
  wire  _T_37 = _T_25 | _T_36; // @[Misc.scala 213:29]
  wire  _T_38 = auto_mem_in_ar_bits_addr[1] & _T_31; // @[Misc.scala 212:27]
  wire  _T_39 = _T_18[0] & _T_38; // @[Misc.scala 213:38]
  wire  _T_40 = _T_28 | _T_39; // @[Misc.scala 213:29]
  wire  _T_41 = auto_mem_in_ar_bits_addr[1] & auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  wire  _T_42 = _T_18[0] & _T_41; // @[Misc.scala 213:38]
  wire  _T_43 = _T_28 | _T_42; // @[Misc.scala 213:29]
  wire [3:0] _T_46 = {_T_43,_T_40,_T_37,_T_34}; // @[Cat.scala 29:58]
  wire [3:0] _T_48 = auto_mem_in_ar_valid ? _T_46 : auto_mem_in_w_bits_strb; // @[RegisterRouter.scala 54:25]
  wire [7:0] _T_67 = _T_48[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_69 = _T_48[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_71 = _T_48[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_73 = _T_48[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_76 = {_T_73,_T_71,_T_69,_T_67}; // @[Cat.scala 29:58]
  wire  _T_95 = _T_76 == 32'hffffffff; // @[RegisterRouter.scala 59:16]
  wire  _T_148 = _T_5 & _T_49_ready; // @[RegisterRouter.scala 59:16]
  wire [1:0] _T_142 = 2'h1 << _T_13[2]; // @[OneHot.scala 58:35]
  wire  _T_165 = _T_148 & _T_6; // @[RegisterRouter.scala 59:16]
  wire  _T_172 = _T_165 & _T_142[1]; // @[RegisterRouter.scala 59:16]
  wire  _T_173 = _T_172 & _T_55; // @[RegisterRouter.scala 59:16]
  wire  _T_102 = _T_173 & _T_95; // @[RegisterRouter.scala 59:16]
  wire  _T_167 = _T_165 & _T_142[0]; // @[RegisterRouter.scala 59:16]
  wire  _T_168 = _T_167 & _T_55; // @[RegisterRouter.scala 59:16]
  wire  _T_125 = _T_168 & _T_95; // @[RegisterRouter.scala 59:16]
  wire  _GEN_11 = _T_13[2] ? _T_55 : _T_55; // @[MuxLiteral.scala 48:10]
  wire [31:0] _GEN_13 = _T_13[2] ? maskReg : ctrlReg; // @[MuxLiteral.scala 48:10]
  wire  _T_223_bits_read = Queue_io_deq_bits_read; // @[Decoupled.scala 317:19 Decoupled.scala 318:14]
  wire  _T_223_valid = Queue_io_deq_valid; // @[Decoupled.scala 317:19 Decoupled.scala 319:15]
  wire  _T_226 = ~_T_223_bits_read; // @[RegisterRouter.scala 65:29]
  wire  readyOR = auto_stream_out_0_ready | auto_stream_out_1_ready; // @[Splitter.scala 45:34]
  wire  readyAND = auto_stream_out_0_ready & auto_stream_out_1_ready; // @[Splitter.scala 46:34]
  wire  _T_229 = ctrlReg == 32'h0; // @[Splitter.scala 49:19]
  wire  _T_230 = ctrlReg == 32'h1; // @[Splitter.scala 52:24]
  wire  _GEN_14 = _T_230 & readyOR; // @[Splitter.scala 52:33]
  wire  _T_233 = ~maskReg[0]; // @[Splitter.scala 62:34]
  wire  _T_237 = ~maskReg[1]; // @[Splitter.scala 62:34]
  Queue Queue ( // @[Decoupled.scala 296:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_read(Queue_io_enq_bits_read),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_extra(Queue_io_enq_bits_extra),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_read(Queue_io_deq_bits_read),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_extra(Queue_io_deq_bits_extra)
  );
  assign auto_mem_in_aw_ready = _T_7 & auto_mem_in_w_valid; // @[LazyModule.scala 173:31]
  assign auto_mem_in_w_ready = _T_7 & auto_mem_in_aw_valid; // @[LazyModule.scala 173:31]
  assign auto_mem_in_b_valid = _T_223_valid & _T_226; // @[LazyModule.scala 173:31]
  assign auto_mem_in_b_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_mem_in_ar_ready = Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_valid = _T_223_valid & _T_223_bits_read; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 173:31]
  assign auto_stream_in_ready = _T_229 ? readyAND : _GEN_14; // @[LazyModule.scala 173:31]
  assign auto_stream_out_1_valid = auto_stream_in_valid & _T_237; // @[LazyModule.scala 173:49]
  assign auto_stream_out_1_bits_data = auto_stream_in_bits_data; // @[LazyModule.scala 173:49]
  assign auto_stream_out_1_bits_last = auto_stream_in_bits_last; // @[LazyModule.scala 173:49]
  assign auto_stream_out_0_valid = auto_stream_in_valid & _T_233; // @[LazyModule.scala 173:49]
  assign auto_stream_out_0_bits_data = auto_stream_in_bits_data; // @[LazyModule.scala 173:49]
  assign auto_stream_out_0_bits_last = auto_stream_in_bits_last; // @[LazyModule.scala 173:49]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_mem_in_ar_valid | _T_4; // @[Decoupled.scala 297:22]
  assign Queue_io_enq_bits_read = auto_mem_in_ar_valid; // @[Decoupled.scala 298:21]
  assign Queue_io_enq_bits_data = _GEN_11 ? _GEN_13 : 32'h0; // @[Decoupled.scala 298:21]
  assign Queue_io_enq_bits_extra = auto_mem_in_ar_valid ? auto_mem_in_ar_bits_id : auto_mem_in_aw_bits_id; // @[Decoupled.scala 298:21]
  assign Queue_io_deq_ready = _T_223_bits_read ? auto_mem_in_r_ready : auto_mem_in_b_ready; // @[Decoupled.scala 320:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ctrlReg = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  maskReg = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      ctrlReg <= 32'h0;
    end else if (_T_125) begin
      ctrlReg <= auto_mem_in_w_bits_data;
    end
    if (reset) begin
      maskReg <= 32'h0;
    end else if (_T_102) begin
      maskReg <= auto_mem_in_w_bits_data;
    end
  end
endmodule
module AXI4StreamMux_2(
  input         clock,
  input         reset,
  output        auto_register_in_aw_ready,
  input         auto_register_in_aw_valid,
  input         auto_register_in_aw_bits_id,
  input  [29:0] auto_register_in_aw_bits_addr,
  output        auto_register_in_w_ready,
  input         auto_register_in_w_valid,
  input  [31:0] auto_register_in_w_bits_data,
  input  [3:0]  auto_register_in_w_bits_strb,
  input         auto_register_in_b_ready,
  output        auto_register_in_b_valid,
  output        auto_register_in_b_bits_id,
  output        auto_register_in_ar_ready,
  input         auto_register_in_ar_valid,
  input         auto_register_in_ar_bits_id,
  input  [29:0] auto_register_in_ar_bits_addr,
  input  [2:0]  auto_register_in_ar_bits_size,
  input         auto_register_in_r_ready,
  output        auto_register_in_r_valid,
  output        auto_register_in_r_bits_id,
  output [31:0] auto_register_in_r_bits_data,
  output        auto_stream_in_2_ready,
  input         auto_stream_in_2_valid,
  input  [31:0] auto_stream_in_2_bits_data,
  input         auto_stream_in_2_bits_last,
  output        auto_stream_in_1_ready,
  input         auto_stream_in_1_valid,
  input  [31:0] auto_stream_in_1_bits_data,
  input         auto_stream_in_1_bits_last,
  output        auto_stream_in_0_ready,
  input         auto_stream_in_0_valid,
  input  [31:0] auto_stream_in_0_bits_data,
  input         auto_stream_in_0_bits_last,
  input         auto_stream_out_0_ready,
  output        auto_stream_out_0_valid,
  output [31:0] auto_stream_out_0_bits_data,
  output        auto_stream_out_0_bits_last
);
  wire  Queue_clock; // @[Decoupled.scala 296:21]
  wire  Queue_reset; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_bits_read; // @[Decoupled.scala 296:21]
  wire [31:0] Queue_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_bits_extra; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_bits_read; // @[Decoupled.scala 296:21]
  wire [31:0] Queue_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_bits_extra; // @[Decoupled.scala 296:21]
  reg [2:0] sels_0; // @[Mux.scala 32:23]
  reg [31:0] _RAND_0;
  reg [2:0] sels_1; // @[Mux.scala 32:23]
  reg [31:0] _RAND_1;
  wire  _T_3 = sels_0 == 3'h0; // @[Mux.scala 45:28]
  wire  _GEN_7 = _T_3 & auto_stream_in_0_valid; // @[Mux.scala 45:41]
  wire  _GEN_8 = _T_3 & auto_stream_out_0_ready; // @[Mux.scala 45:41]
  wire  _T_4 = sels_0 == 3'h1; // @[Mux.scala 45:28]
  wire  _GEN_12 = _T_4 ? auto_stream_in_1_bits_last : auto_stream_in_0_bits_last; // @[Mux.scala 45:41]
  wire [31:0] _GEN_15 = _T_4 ? auto_stream_in_1_bits_data : auto_stream_in_0_bits_data; // @[Mux.scala 45:41]
  wire  _GEN_16 = _T_4 ? auto_stream_in_1_valid : _GEN_7; // @[Mux.scala 45:41]
  wire  _GEN_17 = _T_4 & auto_stream_out_0_ready; // @[Mux.scala 45:41]
  wire  _T_5 = sels_0 == 3'h2; // @[Mux.scala 45:28]
  wire  _GEN_21 = _T_5 ? auto_stream_in_2_bits_last : _GEN_12; // @[Mux.scala 45:41]
  wire [31:0] _GEN_24 = _T_5 ? auto_stream_in_2_bits_data : _GEN_15; // @[Mux.scala 45:41]
  wire  _GEN_25 = _T_5 ? auto_stream_in_2_valid : _GEN_16; // @[Mux.scala 45:41]
  wire  _GEN_26 = _T_5 & auto_stream_out_0_ready; // @[Mux.scala 45:41]
  wire  _T_6 = sels_0 == 3'h3; // @[Mux.scala 45:28]
  wire  _GEN_30 = _T_6 ? 1'h0 : _GEN_21; // @[Mux.scala 45:41]
  wire [31:0] _GEN_33 = _T_6 ? 32'hffffffff : _GEN_24; // @[Mux.scala 45:41]
  wire  _GEN_34 = _T_6 | _GEN_25; // @[Mux.scala 45:41]
  wire  _T_7 = sels_0 == 3'h4; // @[Mux.scala 45:28]
  wire  _T_8 = sels_0 == sels_1; // @[Mux.scala 40:46]
  wire [2:0] _T_10 = _T_8 ? 3'h5 : sels_1; // @[Mux.scala 41:29]
  wire  _T_11 = _T_10 == 3'h0; // @[Mux.scala 45:28]
  wire  _T_12 = _T_10 == 3'h1; // @[Mux.scala 45:28]
  wire  _T_13 = _T_10 == 3'h2; // @[Mux.scala 45:28]
  wire  _T_17 = auto_register_in_aw_valid & auto_register_in_w_valid; // @[RegisterRouter.scala 40:39]
  wire  _T_18 = auto_register_in_ar_valid | _T_17; // @[RegisterRouter.scala 40:26]
  wire  _T_19 = ~auto_register_in_ar_valid; // @[RegisterRouter.scala 42:29]
  wire  _T_62_ready = Queue_io_enq_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 299:17]
  wire [29:0] _T_26 = auto_register_in_ar_valid ? auto_register_in_ar_bits_addr : auto_register_in_aw_bits_addr; // @[RegisterRouter.scala 48:19]
  wire [1:0] _T_66 = _T_26[3:2] & 2'h2; // @[RegisterRouter.scala 59:16]
  wire  _T_68 = _T_66 == 2'h0; // @[RegisterRouter.scala 59:16]
  wire  _T_20 = _T_62_ready & _T_19; // @[RegisterRouter.scala 42:26]
  wire [1:0] _T_29 = 2'h1 << auto_register_in_ar_bits_size[0]; // @[OneHot.scala 65:12]
  wire [1:0] _T_31 = _T_29 | 2'h1; // @[Misc.scala 200:81]
  wire  _T_32 = auto_register_in_ar_bits_size >= 3'h2; // @[Misc.scala 204:21]
  wire  _T_35 = ~auto_register_in_ar_bits_addr[1]; // @[Misc.scala 209:20]
  wire  _T_37 = _T_31[1] & _T_35; // @[Misc.scala 213:38]
  wire  _T_38 = _T_32 | _T_37; // @[Misc.scala 213:29]
  wire  _T_40 = _T_31[1] & auto_register_in_ar_bits_addr[1]; // @[Misc.scala 213:38]
  wire  _T_41 = _T_32 | _T_40; // @[Misc.scala 213:29]
  wire  _T_44 = ~auto_register_in_ar_bits_addr[0]; // @[Misc.scala 209:20]
  wire  _T_45 = _T_35 & _T_44; // @[Misc.scala 212:27]
  wire  _T_46 = _T_31[0] & _T_45; // @[Misc.scala 213:38]
  wire  _T_47 = _T_38 | _T_46; // @[Misc.scala 213:29]
  wire  _T_48 = _T_35 & auto_register_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  wire  _T_49 = _T_31[0] & _T_48; // @[Misc.scala 213:38]
  wire  _T_50 = _T_38 | _T_49; // @[Misc.scala 213:29]
  wire  _T_51 = auto_register_in_ar_bits_addr[1] & _T_44; // @[Misc.scala 212:27]
  wire  _T_52 = _T_31[0] & _T_51; // @[Misc.scala 213:38]
  wire  _T_53 = _T_41 | _T_52; // @[Misc.scala 213:29]
  wire  _T_54 = auto_register_in_ar_bits_addr[1] & auto_register_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  wire  _T_55 = _T_31[0] & _T_54; // @[Misc.scala 213:38]
  wire  _T_56 = _T_41 | _T_55; // @[Misc.scala 213:29]
  wire [3:0] _T_59 = {_T_56,_T_53,_T_50,_T_47}; // @[Cat.scala 29:58]
  wire [3:0] _T_61 = auto_register_in_ar_valid ? _T_59 : auto_register_in_w_bits_strb; // @[RegisterRouter.scala 54:25]
  wire [7:0] _T_80 = _T_61[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_82 = _T_61[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_84 = _T_61[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_86 = _T_61[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_89 = {_T_86,_T_84,_T_82,_T_80}; // @[Cat.scala 29:58]
  wire  _T_108 = _T_89[2:0] == 3'h7; // @[RegisterRouter.scala 59:16]
  wire  _T_161 = _T_18 & _T_62_ready; // @[RegisterRouter.scala 59:16]
  wire [1:0] _T_155 = 2'h1 << _T_26[2]; // @[OneHot.scala 58:35]
  wire  _T_178 = _T_161 & _T_19; // @[RegisterRouter.scala 59:16]
  wire  _T_185 = _T_178 & _T_155[1]; // @[RegisterRouter.scala 59:16]
  wire  _T_186 = _T_185 & _T_68; // @[RegisterRouter.scala 59:16]
  wire  _T_115 = _T_186 & _T_108; // @[RegisterRouter.scala 59:16]
  wire  _T_180 = _T_178 & _T_155[0]; // @[RegisterRouter.scala 59:16]
  wire  _T_181 = _T_180 & _T_68; // @[RegisterRouter.scala 59:16]
  wire  _T_138 = _T_181 & _T_108; // @[RegisterRouter.scala 59:16]
  wire  _GEN_101 = _T_26[2] ? _T_68 : _T_68; // @[MuxLiteral.scala 48:10]
  wire [2:0] _GEN_103 = _T_26[2] ? sels_1 : sels_0; // @[MuxLiteral.scala 48:10]
  wire [2:0] _T_235 = _GEN_101 ? _GEN_103 : 3'h0; // @[RegisterRouter.scala 59:16]
  wire  _T_236_bits_read = Queue_io_deq_bits_read; // @[Decoupled.scala 317:19 Decoupled.scala 318:14]
  wire  _T_236_valid = Queue_io_deq_valid; // @[Decoupled.scala 317:19 Decoupled.scala 319:15]
  wire  _T_239 = ~_T_236_bits_read; // @[RegisterRouter.scala 65:29]
  Queue Queue ( // @[Decoupled.scala 296:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_read(Queue_io_enq_bits_read),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_extra(Queue_io_enq_bits_extra),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_read(Queue_io_deq_bits_read),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_extra(Queue_io_deq_bits_extra)
  );
  assign auto_register_in_aw_ready = _T_20 & auto_register_in_w_valid; // @[LazyModule.scala 173:31]
  assign auto_register_in_w_ready = _T_20 & auto_register_in_aw_valid; // @[LazyModule.scala 173:31]
  assign auto_register_in_b_valid = _T_236_valid & _T_239; // @[LazyModule.scala 173:31]
  assign auto_register_in_b_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_register_in_ar_ready = Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_register_in_r_valid = _T_236_valid & _T_236_bits_read; // @[LazyModule.scala 173:31]
  assign auto_register_in_r_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_register_in_r_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 173:31]
  assign auto_stream_in_2_ready = _T_13 | _GEN_26; // @[LazyModule.scala 173:31]
  assign auto_stream_in_1_ready = _T_12 | _GEN_17; // @[LazyModule.scala 173:31]
  assign auto_stream_in_0_ready = _T_11 | _GEN_8; // @[LazyModule.scala 173:31]
  assign auto_stream_out_0_valid = _T_7 | _GEN_34; // @[LazyModule.scala 173:49]
  assign auto_stream_out_0_bits_data = _T_7 ? 32'h0 : _GEN_33; // @[LazyModule.scala 173:49]
  assign auto_stream_out_0_bits_last = _T_7 ? 1'h0 : _GEN_30; // @[LazyModule.scala 173:49]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_register_in_ar_valid | _T_17; // @[Decoupled.scala 297:22]
  assign Queue_io_enq_bits_read = auto_register_in_ar_valid; // @[Decoupled.scala 298:21]
  assign Queue_io_enq_bits_data = {{29'd0}, _T_235}; // @[Decoupled.scala 298:21]
  assign Queue_io_enq_bits_extra = auto_register_in_ar_valid ? auto_register_in_ar_bits_id : auto_register_in_aw_bits_id; // @[Decoupled.scala 298:21]
  assign Queue_io_deq_ready = _T_236_bits_read ? auto_register_in_r_ready : auto_register_in_b_ready; // @[Decoupled.scala 320:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  sels_0 = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  sels_1 = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      sels_0 <= 3'h5;
    end else if (_T_138) begin
      sels_0 <= auto_register_in_w_bits_data[2:0];
    end
    if (reset) begin
      sels_1 <= 3'h5;
    end else if (_T_115) begin
      sels_1 <= auto_register_in_w_bits_data[2:0];
    end
  end
endmodule
module SDFStageRadix22(
  input         clock,
  input         reset,
  input  [15:0] io_in_real,
  input  [15:0] io_in_imag,
  output [15:0] io_out_real,
  output [15:0] io_out_imag,
  input  [6:0]  io_cntr,
  input         io_en
);
  wire  load_input = io_cntr < 7'h40; // @[SDFChainRadix22.scala 426:66]
  reg [15:0] shift_out_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_0;
  wire [16:0] butt_outputs_1_real = $signed(shift_out_real) - $signed(io_in_real); // @[FixedPointTypeClass.scala 33:22]
  wire [17:0] _T_236 = {$signed(butt_outputs_1_real), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_238 = _T_236[17:1]; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_241 = $signed(_T_238) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] butterfly_outputs_1_real = _T_241[16:1]; // @[FixedPointTypeClass.scala 176:41]
  reg [15:0] shift_out_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1;
  wire [16:0] butt_outputs_1_imag = $signed(shift_out_imag) - $signed(io_in_imag); // @[FixedPointTypeClass.scala 33:22]
  wire [17:0] _T_243 = {$signed(butt_outputs_1_imag), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_245 = _T_243[17:1]; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_248 = $signed(_T_245) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] butterfly_outputs_1_imag = _T_248[16:1]; // @[FixedPointTypeClass.scala 176:41]
  reg [15:0] _T_21_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2;
  reg [15:0] _T_21_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3;
  reg [15:0] _T_24_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4;
  reg [15:0] _T_24_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5;
  reg [15:0] _T_27_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6;
  reg [15:0] _T_27_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7;
  reg [15:0] _T_30_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8;
  reg [15:0] _T_30_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9;
  reg [15:0] _T_33_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10;
  reg [15:0] _T_33_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11;
  reg [15:0] _T_36_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12;
  reg [15:0] _T_36_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_13;
  reg [15:0] _T_39_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_14;
  reg [15:0] _T_39_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_15;
  reg [15:0] _T_42_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_16;
  reg [15:0] _T_42_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_17;
  reg [15:0] _T_45_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_18;
  reg [15:0] _T_45_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_19;
  reg [15:0] _T_48_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_20;
  reg [15:0] _T_48_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_21;
  reg [15:0] _T_51_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_22;
  reg [15:0] _T_51_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_23;
  reg [15:0] _T_54_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_24;
  reg [15:0] _T_54_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_25;
  reg [15:0] _T_57_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_26;
  reg [15:0] _T_57_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_27;
  reg [15:0] _T_60_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_28;
  reg [15:0] _T_60_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_29;
  reg [15:0] _T_63_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_30;
  reg [15:0] _T_63_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_31;
  reg [15:0] _T_66_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_32;
  reg [15:0] _T_66_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_33;
  reg [15:0] _T_69_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_34;
  reg [15:0] _T_69_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_35;
  reg [15:0] _T_72_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_36;
  reg [15:0] _T_72_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_37;
  reg [15:0] _T_75_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_38;
  reg [15:0] _T_75_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_39;
  reg [15:0] _T_78_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_40;
  reg [15:0] _T_78_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_41;
  reg [15:0] _T_81_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_42;
  reg [15:0] _T_81_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_43;
  reg [15:0] _T_84_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_44;
  reg [15:0] _T_84_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_45;
  reg [15:0] _T_87_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_46;
  reg [15:0] _T_87_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_47;
  reg [15:0] _T_90_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_48;
  reg [15:0] _T_90_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_49;
  reg [15:0] _T_93_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_50;
  reg [15:0] _T_93_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_51;
  reg [15:0] _T_96_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_52;
  reg [15:0] _T_96_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_53;
  reg [15:0] _T_99_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_54;
  reg [15:0] _T_99_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_55;
  reg [15:0] _T_102_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_56;
  reg [15:0] _T_102_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_57;
  reg [15:0] _T_105_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_58;
  reg [15:0] _T_105_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_59;
  reg [15:0] _T_108_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_60;
  reg [15:0] _T_108_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_61;
  reg [15:0] _T_111_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_62;
  reg [15:0] _T_111_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_63;
  reg [15:0] _T_114_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_64;
  reg [15:0] _T_114_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_65;
  reg [15:0] _T_117_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_66;
  reg [15:0] _T_117_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_67;
  reg [15:0] _T_120_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_68;
  reg [15:0] _T_120_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_69;
  reg [15:0] _T_123_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_70;
  reg [15:0] _T_123_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_71;
  reg [15:0] _T_126_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_72;
  reg [15:0] _T_126_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_73;
  reg [15:0] _T_129_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_74;
  reg [15:0] _T_129_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_75;
  reg [15:0] _T_132_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_76;
  reg [15:0] _T_132_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_77;
  reg [15:0] _T_135_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_78;
  reg [15:0] _T_135_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_79;
  reg [15:0] _T_138_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_80;
  reg [15:0] _T_138_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_81;
  reg [15:0] _T_141_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_82;
  reg [15:0] _T_141_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_83;
  reg [15:0] _T_144_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_84;
  reg [15:0] _T_144_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_85;
  reg [15:0] _T_147_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_86;
  reg [15:0] _T_147_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_87;
  reg [15:0] _T_150_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_88;
  reg [15:0] _T_150_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_89;
  reg [15:0] _T_153_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_90;
  reg [15:0] _T_153_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_91;
  reg [15:0] _T_156_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_92;
  reg [15:0] _T_156_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_93;
  reg [15:0] _T_159_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_94;
  reg [15:0] _T_159_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_95;
  reg [15:0] _T_162_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_96;
  reg [15:0] _T_162_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_97;
  reg [15:0] _T_165_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_98;
  reg [15:0] _T_165_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_99;
  reg [15:0] _T_168_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_100;
  reg [15:0] _T_168_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_101;
  reg [15:0] _T_171_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_102;
  reg [15:0] _T_171_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_103;
  reg [15:0] _T_174_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_104;
  reg [15:0] _T_174_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_105;
  reg [15:0] _T_177_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_106;
  reg [15:0] _T_177_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_107;
  reg [15:0] _T_180_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_108;
  reg [15:0] _T_180_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_109;
  reg [15:0] _T_183_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_110;
  reg [15:0] _T_183_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_111;
  reg [15:0] _T_186_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_112;
  reg [15:0] _T_186_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_113;
  reg [15:0] _T_189_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_114;
  reg [15:0] _T_189_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_115;
  reg [15:0] _T_192_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_116;
  reg [15:0] _T_192_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_117;
  reg [15:0] _T_195_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_118;
  reg [15:0] _T_195_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_119;
  reg [15:0] _T_198_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_120;
  reg [15:0] _T_198_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_121;
  reg [15:0] _T_201_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_122;
  reg [15:0] _T_201_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_123;
  reg [15:0] _T_204_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_124;
  reg [15:0] _T_204_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_125;
  reg [15:0] _T_207_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_126;
  reg [15:0] _T_207_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_127;
  wire [16:0] butt_outputs_0_real = $signed(shift_out_real) + $signed(io_in_real); // @[FixedPointTypeClass.scala 24:22]
  wire [16:0] butt_outputs_0_imag = $signed(shift_out_imag) + $signed(io_in_imag); // @[FixedPointTypeClass.scala 24:22]
  wire [17:0] _T_219 = {$signed(butt_outputs_0_real), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_221 = _T_219[17:1]; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_224 = $signed(_T_221) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  wire [17:0] _T_226 = {$signed(butt_outputs_0_imag), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_228 = _T_226[17:1]; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_231 = $signed(_T_228) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  reg [15:0] feedback_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_128;
  reg [15:0] feedback_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_129;
  reg [15:0] butt_out_0_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_130;
  reg [15:0] butt_out_0_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_131;
  reg  load_output; // @[Reg.scala 27:20]
  reg [31:0] _RAND_132;
  assign io_out_real = load_output ? $signed(feedback_real) : $signed(butt_out_0_real); // @[SDFChainRadix22.scala 422:10]
  assign io_out_imag = load_output ? $signed(feedback_imag) : $signed(butt_out_0_imag); // @[SDFChainRadix22.scala 422:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  shift_out_real = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  shift_out_imag = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_21_real = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_21_imag = _RAND_3[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_24_real = _RAND_4[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_24_imag = _RAND_5[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_27_real = _RAND_6[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_27_imag = _RAND_7[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_30_real = _RAND_8[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_30_imag = _RAND_9[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_33_real = _RAND_10[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_33_imag = _RAND_11[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_36_real = _RAND_12[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_36_imag = _RAND_13[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_39_real = _RAND_14[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_39_imag = _RAND_15[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_42_real = _RAND_16[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_42_imag = _RAND_17[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_45_real = _RAND_18[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_45_imag = _RAND_19[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_48_real = _RAND_20[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_48_imag = _RAND_21[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_51_real = _RAND_22[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_51_imag = _RAND_23[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_54_real = _RAND_24[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_54_imag = _RAND_25[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_57_real = _RAND_26[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T_57_imag = _RAND_27[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_60_real = _RAND_28[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_60_imag = _RAND_29[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_63_real = _RAND_30[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T_63_imag = _RAND_31[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _T_66_real = _RAND_32[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _T_66_imag = _RAND_33[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _T_69_real = _RAND_34[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _T_69_imag = _RAND_35[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _T_72_real = _RAND_36[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _T_72_imag = _RAND_37[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _T_75_real = _RAND_38[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _T_75_imag = _RAND_39[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _T_78_real = _RAND_40[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  _T_78_imag = _RAND_41[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  _T_81_real = _RAND_42[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  _T_81_imag = _RAND_43[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  _T_84_real = _RAND_44[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  _T_84_imag = _RAND_45[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  _T_87_real = _RAND_46[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  _T_87_imag = _RAND_47[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  _T_90_real = _RAND_48[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  _T_90_imag = _RAND_49[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  _T_93_real = _RAND_50[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  _T_93_imag = _RAND_51[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  _T_96_real = _RAND_52[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  _T_96_imag = _RAND_53[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  _T_99_real = _RAND_54[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  _T_99_imag = _RAND_55[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  _T_102_real = _RAND_56[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  _T_102_imag = _RAND_57[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  _T_105_real = _RAND_58[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  _T_105_imag = _RAND_59[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  _T_108_real = _RAND_60[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  _T_108_imag = _RAND_61[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  _T_111_real = _RAND_62[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  _T_111_imag = _RAND_63[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  _T_114_real = _RAND_64[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  _T_114_imag = _RAND_65[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  _T_117_real = _RAND_66[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  _T_117_imag = _RAND_67[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  _T_120_real = _RAND_68[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  _T_120_imag = _RAND_69[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  _T_123_real = _RAND_70[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  _T_123_imag = _RAND_71[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  _T_126_real = _RAND_72[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  _T_126_imag = _RAND_73[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  _T_129_real = _RAND_74[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  _T_129_imag = _RAND_75[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  _T_132_real = _RAND_76[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  _T_132_imag = _RAND_77[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  _T_135_real = _RAND_78[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  _T_135_imag = _RAND_79[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  _T_138_real = _RAND_80[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  _T_138_imag = _RAND_81[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  _T_141_real = _RAND_82[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  _T_141_imag = _RAND_83[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  _T_144_real = _RAND_84[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  _T_144_imag = _RAND_85[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  _T_147_real = _RAND_86[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  _T_147_imag = _RAND_87[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  _T_150_real = _RAND_88[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  _T_150_imag = _RAND_89[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  _T_153_real = _RAND_90[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  _T_153_imag = _RAND_91[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  _T_156_real = _RAND_92[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  _T_156_imag = _RAND_93[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  _T_159_real = _RAND_94[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  _T_159_imag = _RAND_95[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  _T_162_real = _RAND_96[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  _T_162_imag = _RAND_97[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  _T_165_real = _RAND_98[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  _T_165_imag = _RAND_99[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  _T_168_real = _RAND_100[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  _T_168_imag = _RAND_101[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  _T_171_real = _RAND_102[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  _T_171_imag = _RAND_103[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  _T_174_real = _RAND_104[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  _T_174_imag = _RAND_105[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  _T_177_real = _RAND_106[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  _T_177_imag = _RAND_107[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  _T_180_real = _RAND_108[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  _T_180_imag = _RAND_109[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  _T_183_real = _RAND_110[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  _T_183_imag = _RAND_111[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  _T_186_real = _RAND_112[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  _T_186_imag = _RAND_113[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  _T_189_real = _RAND_114[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  _T_189_imag = _RAND_115[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  _T_192_real = _RAND_116[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  _T_192_imag = _RAND_117[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  _T_195_real = _RAND_118[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  _T_195_imag = _RAND_119[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  _T_198_real = _RAND_120[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  _T_198_imag = _RAND_121[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  _T_201_real = _RAND_122[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  _T_201_imag = _RAND_123[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  _T_204_real = _RAND_124[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  _T_204_imag = _RAND_125[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  _T_207_real = _RAND_126[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  _T_207_imag = _RAND_127[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  feedback_real = _RAND_128[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{`RANDOM}};
  feedback_imag = _RAND_129[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{`RANDOM}};
  butt_out_0_real = _RAND_130[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{`RANDOM}};
  butt_out_0_imag = _RAND_131[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{`RANDOM}};
  load_output = _RAND_132[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (io_en) begin
      shift_out_real <= _T_207_real;
    end
    if (io_en) begin
      shift_out_imag <= _T_207_imag;
    end
    if (io_en) begin
      if (load_input) begin
        _T_21_real <= io_in_real;
      end else begin
        _T_21_real <= butterfly_outputs_1_real;
      end
    end
    if (io_en) begin
      if (load_input) begin
        _T_21_imag <= io_in_imag;
      end else begin
        _T_21_imag <= butterfly_outputs_1_imag;
      end
    end
    if (io_en) begin
      _T_24_real <= _T_21_real;
    end
    if (io_en) begin
      _T_24_imag <= _T_21_imag;
    end
    if (io_en) begin
      _T_27_real <= _T_24_real;
    end
    if (io_en) begin
      _T_27_imag <= _T_24_imag;
    end
    if (io_en) begin
      _T_30_real <= _T_27_real;
    end
    if (io_en) begin
      _T_30_imag <= _T_27_imag;
    end
    if (io_en) begin
      _T_33_real <= _T_30_real;
    end
    if (io_en) begin
      _T_33_imag <= _T_30_imag;
    end
    if (io_en) begin
      _T_36_real <= _T_33_real;
    end
    if (io_en) begin
      _T_36_imag <= _T_33_imag;
    end
    if (io_en) begin
      _T_39_real <= _T_36_real;
    end
    if (io_en) begin
      _T_39_imag <= _T_36_imag;
    end
    if (io_en) begin
      _T_42_real <= _T_39_real;
    end
    if (io_en) begin
      _T_42_imag <= _T_39_imag;
    end
    if (io_en) begin
      _T_45_real <= _T_42_real;
    end
    if (io_en) begin
      _T_45_imag <= _T_42_imag;
    end
    if (io_en) begin
      _T_48_real <= _T_45_real;
    end
    if (io_en) begin
      _T_48_imag <= _T_45_imag;
    end
    if (io_en) begin
      _T_51_real <= _T_48_real;
    end
    if (io_en) begin
      _T_51_imag <= _T_48_imag;
    end
    if (io_en) begin
      _T_54_real <= _T_51_real;
    end
    if (io_en) begin
      _T_54_imag <= _T_51_imag;
    end
    if (io_en) begin
      _T_57_real <= _T_54_real;
    end
    if (io_en) begin
      _T_57_imag <= _T_54_imag;
    end
    if (io_en) begin
      _T_60_real <= _T_57_real;
    end
    if (io_en) begin
      _T_60_imag <= _T_57_imag;
    end
    if (io_en) begin
      _T_63_real <= _T_60_real;
    end
    if (io_en) begin
      _T_63_imag <= _T_60_imag;
    end
    if (io_en) begin
      _T_66_real <= _T_63_real;
    end
    if (io_en) begin
      _T_66_imag <= _T_63_imag;
    end
    if (io_en) begin
      _T_69_real <= _T_66_real;
    end
    if (io_en) begin
      _T_69_imag <= _T_66_imag;
    end
    if (io_en) begin
      _T_72_real <= _T_69_real;
    end
    if (io_en) begin
      _T_72_imag <= _T_69_imag;
    end
    if (io_en) begin
      _T_75_real <= _T_72_real;
    end
    if (io_en) begin
      _T_75_imag <= _T_72_imag;
    end
    if (io_en) begin
      _T_78_real <= _T_75_real;
    end
    if (io_en) begin
      _T_78_imag <= _T_75_imag;
    end
    if (io_en) begin
      _T_81_real <= _T_78_real;
    end
    if (io_en) begin
      _T_81_imag <= _T_78_imag;
    end
    if (io_en) begin
      _T_84_real <= _T_81_real;
    end
    if (io_en) begin
      _T_84_imag <= _T_81_imag;
    end
    if (io_en) begin
      _T_87_real <= _T_84_real;
    end
    if (io_en) begin
      _T_87_imag <= _T_84_imag;
    end
    if (io_en) begin
      _T_90_real <= _T_87_real;
    end
    if (io_en) begin
      _T_90_imag <= _T_87_imag;
    end
    if (io_en) begin
      _T_93_real <= _T_90_real;
    end
    if (io_en) begin
      _T_93_imag <= _T_90_imag;
    end
    if (io_en) begin
      _T_96_real <= _T_93_real;
    end
    if (io_en) begin
      _T_96_imag <= _T_93_imag;
    end
    if (io_en) begin
      _T_99_real <= _T_96_real;
    end
    if (io_en) begin
      _T_99_imag <= _T_96_imag;
    end
    if (io_en) begin
      _T_102_real <= _T_99_real;
    end
    if (io_en) begin
      _T_102_imag <= _T_99_imag;
    end
    if (io_en) begin
      _T_105_real <= _T_102_real;
    end
    if (io_en) begin
      _T_105_imag <= _T_102_imag;
    end
    if (io_en) begin
      _T_108_real <= _T_105_real;
    end
    if (io_en) begin
      _T_108_imag <= _T_105_imag;
    end
    if (io_en) begin
      _T_111_real <= _T_108_real;
    end
    if (io_en) begin
      _T_111_imag <= _T_108_imag;
    end
    if (io_en) begin
      _T_114_real <= _T_111_real;
    end
    if (io_en) begin
      _T_114_imag <= _T_111_imag;
    end
    if (io_en) begin
      _T_117_real <= _T_114_real;
    end
    if (io_en) begin
      _T_117_imag <= _T_114_imag;
    end
    if (io_en) begin
      _T_120_real <= _T_117_real;
    end
    if (io_en) begin
      _T_120_imag <= _T_117_imag;
    end
    if (io_en) begin
      _T_123_real <= _T_120_real;
    end
    if (io_en) begin
      _T_123_imag <= _T_120_imag;
    end
    if (io_en) begin
      _T_126_real <= _T_123_real;
    end
    if (io_en) begin
      _T_126_imag <= _T_123_imag;
    end
    if (io_en) begin
      _T_129_real <= _T_126_real;
    end
    if (io_en) begin
      _T_129_imag <= _T_126_imag;
    end
    if (io_en) begin
      _T_132_real <= _T_129_real;
    end
    if (io_en) begin
      _T_132_imag <= _T_129_imag;
    end
    if (io_en) begin
      _T_135_real <= _T_132_real;
    end
    if (io_en) begin
      _T_135_imag <= _T_132_imag;
    end
    if (io_en) begin
      _T_138_real <= _T_135_real;
    end
    if (io_en) begin
      _T_138_imag <= _T_135_imag;
    end
    if (io_en) begin
      _T_141_real <= _T_138_real;
    end
    if (io_en) begin
      _T_141_imag <= _T_138_imag;
    end
    if (io_en) begin
      _T_144_real <= _T_141_real;
    end
    if (io_en) begin
      _T_144_imag <= _T_141_imag;
    end
    if (io_en) begin
      _T_147_real <= _T_144_real;
    end
    if (io_en) begin
      _T_147_imag <= _T_144_imag;
    end
    if (io_en) begin
      _T_150_real <= _T_147_real;
    end
    if (io_en) begin
      _T_150_imag <= _T_147_imag;
    end
    if (io_en) begin
      _T_153_real <= _T_150_real;
    end
    if (io_en) begin
      _T_153_imag <= _T_150_imag;
    end
    if (io_en) begin
      _T_156_real <= _T_153_real;
    end
    if (io_en) begin
      _T_156_imag <= _T_153_imag;
    end
    if (io_en) begin
      _T_159_real <= _T_156_real;
    end
    if (io_en) begin
      _T_159_imag <= _T_156_imag;
    end
    if (io_en) begin
      _T_162_real <= _T_159_real;
    end
    if (io_en) begin
      _T_162_imag <= _T_159_imag;
    end
    if (io_en) begin
      _T_165_real <= _T_162_real;
    end
    if (io_en) begin
      _T_165_imag <= _T_162_imag;
    end
    if (io_en) begin
      _T_168_real <= _T_165_real;
    end
    if (io_en) begin
      _T_168_imag <= _T_165_imag;
    end
    if (io_en) begin
      _T_171_real <= _T_168_real;
    end
    if (io_en) begin
      _T_171_imag <= _T_168_imag;
    end
    if (io_en) begin
      _T_174_real <= _T_171_real;
    end
    if (io_en) begin
      _T_174_imag <= _T_171_imag;
    end
    if (io_en) begin
      _T_177_real <= _T_174_real;
    end
    if (io_en) begin
      _T_177_imag <= _T_174_imag;
    end
    if (io_en) begin
      _T_180_real <= _T_177_real;
    end
    if (io_en) begin
      _T_180_imag <= _T_177_imag;
    end
    if (io_en) begin
      _T_183_real <= _T_180_real;
    end
    if (io_en) begin
      _T_183_imag <= _T_180_imag;
    end
    if (io_en) begin
      _T_186_real <= _T_183_real;
    end
    if (io_en) begin
      _T_186_imag <= _T_183_imag;
    end
    if (io_en) begin
      _T_189_real <= _T_186_real;
    end
    if (io_en) begin
      _T_189_imag <= _T_186_imag;
    end
    if (io_en) begin
      _T_192_real <= _T_189_real;
    end
    if (io_en) begin
      _T_192_imag <= _T_189_imag;
    end
    if (io_en) begin
      _T_195_real <= _T_192_real;
    end
    if (io_en) begin
      _T_195_imag <= _T_192_imag;
    end
    if (io_en) begin
      _T_198_real <= _T_195_real;
    end
    if (io_en) begin
      _T_198_imag <= _T_195_imag;
    end
    if (io_en) begin
      _T_201_real <= _T_198_real;
    end
    if (io_en) begin
      _T_201_imag <= _T_198_imag;
    end
    if (io_en) begin
      _T_204_real <= _T_201_real;
    end
    if (io_en) begin
      _T_204_imag <= _T_201_imag;
    end
    if (io_en) begin
      _T_207_real <= _T_204_real;
    end
    if (io_en) begin
      _T_207_imag <= _T_204_imag;
    end
    feedback_real <= shift_out_real;
    feedback_imag <= shift_out_imag;
    butt_out_0_real <= _T_224[16:1];
    butt_out_0_imag <= _T_231[16:1];
    if (reset) begin
      load_output <= 1'h0;
    end else begin
      load_output <= load_input;
    end
  end
endmodule
module SDFStageRadix22_1(
  input         clock,
  input         reset,
  input  [15:0] io_in_real,
  input  [15:0] io_in_imag,
  output [15:0] io_out_real,
  output [15:0] io_out_imag,
  input  [6:0]  io_cntr,
  input         io_en
);
  wire  load_input = io_cntr < 7'h20; // @[SDFChainRadix22.scala 426:66]
  reg [15:0] shift_out_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_0;
  wire [16:0] butt_outputs_1_real = $signed(shift_out_real) - $signed(io_in_real); // @[FixedPointTypeClass.scala 33:22]
  wire [17:0] _T_140 = {$signed(butt_outputs_1_real), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_142 = _T_140[17:1]; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_145 = $signed(_T_142) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] butterfly_outputs_1_real = _T_145[16:1]; // @[FixedPointTypeClass.scala 176:41]
  reg [15:0] shift_out_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1;
  wire [16:0] butt_outputs_1_imag = $signed(shift_out_imag) - $signed(io_in_imag); // @[FixedPointTypeClass.scala 33:22]
  wire [17:0] _T_147 = {$signed(butt_outputs_1_imag), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_149 = _T_147[17:1]; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_152 = $signed(_T_149) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] butterfly_outputs_1_imag = _T_152[16:1]; // @[FixedPointTypeClass.scala 176:41]
  reg [15:0] _T_21_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2;
  reg [15:0] _T_21_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3;
  reg [15:0] _T_24_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4;
  reg [15:0] _T_24_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5;
  reg [15:0] _T_27_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6;
  reg [15:0] _T_27_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7;
  reg [15:0] _T_30_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8;
  reg [15:0] _T_30_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9;
  reg [15:0] _T_33_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10;
  reg [15:0] _T_33_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11;
  reg [15:0] _T_36_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12;
  reg [15:0] _T_36_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_13;
  reg [15:0] _T_39_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_14;
  reg [15:0] _T_39_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_15;
  reg [15:0] _T_42_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_16;
  reg [15:0] _T_42_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_17;
  reg [15:0] _T_45_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_18;
  reg [15:0] _T_45_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_19;
  reg [15:0] _T_48_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_20;
  reg [15:0] _T_48_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_21;
  reg [15:0] _T_51_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_22;
  reg [15:0] _T_51_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_23;
  reg [15:0] _T_54_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_24;
  reg [15:0] _T_54_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_25;
  reg [15:0] _T_57_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_26;
  reg [15:0] _T_57_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_27;
  reg [15:0] _T_60_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_28;
  reg [15:0] _T_60_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_29;
  reg [15:0] _T_63_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_30;
  reg [15:0] _T_63_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_31;
  reg [15:0] _T_66_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_32;
  reg [15:0] _T_66_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_33;
  reg [15:0] _T_69_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_34;
  reg [15:0] _T_69_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_35;
  reg [15:0] _T_72_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_36;
  reg [15:0] _T_72_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_37;
  reg [15:0] _T_75_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_38;
  reg [15:0] _T_75_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_39;
  reg [15:0] _T_78_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_40;
  reg [15:0] _T_78_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_41;
  reg [15:0] _T_81_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_42;
  reg [15:0] _T_81_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_43;
  reg [15:0] _T_84_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_44;
  reg [15:0] _T_84_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_45;
  reg [15:0] _T_87_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_46;
  reg [15:0] _T_87_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_47;
  reg [15:0] _T_90_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_48;
  reg [15:0] _T_90_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_49;
  reg [15:0] _T_93_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_50;
  reg [15:0] _T_93_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_51;
  reg [15:0] _T_96_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_52;
  reg [15:0] _T_96_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_53;
  reg [15:0] _T_99_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_54;
  reg [15:0] _T_99_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_55;
  reg [15:0] _T_102_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_56;
  reg [15:0] _T_102_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_57;
  reg [15:0] _T_105_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_58;
  reg [15:0] _T_105_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_59;
  reg [15:0] _T_108_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_60;
  reg [15:0] _T_108_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_61;
  reg [15:0] _T_111_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_62;
  reg [15:0] _T_111_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_63;
  wire [16:0] butt_outputs_0_real = $signed(shift_out_real) + $signed(io_in_real); // @[FixedPointTypeClass.scala 24:22]
  wire [16:0] butt_outputs_0_imag = $signed(shift_out_imag) + $signed(io_in_imag); // @[FixedPointTypeClass.scala 24:22]
  wire [17:0] _T_123 = {$signed(butt_outputs_0_real), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_125 = _T_123[17:1]; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_128 = $signed(_T_125) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  wire [17:0] _T_130 = {$signed(butt_outputs_0_imag), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_132 = _T_130[17:1]; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_135 = $signed(_T_132) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  reg [15:0] feedback_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_64;
  reg [15:0] feedback_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_65;
  reg [15:0] butt_out_0_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_66;
  reg [15:0] butt_out_0_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_67;
  reg  load_output; // @[Reg.scala 27:20]
  reg [31:0] _RAND_68;
  assign io_out_real = load_output ? $signed(feedback_real) : $signed(butt_out_0_real); // @[SDFChainRadix22.scala 422:10]
  assign io_out_imag = load_output ? $signed(feedback_imag) : $signed(butt_out_0_imag); // @[SDFChainRadix22.scala 422:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  shift_out_real = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  shift_out_imag = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_21_real = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_21_imag = _RAND_3[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_24_real = _RAND_4[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_24_imag = _RAND_5[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_27_real = _RAND_6[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_27_imag = _RAND_7[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_30_real = _RAND_8[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_30_imag = _RAND_9[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_33_real = _RAND_10[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_33_imag = _RAND_11[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_36_real = _RAND_12[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_36_imag = _RAND_13[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_39_real = _RAND_14[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_39_imag = _RAND_15[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_42_real = _RAND_16[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_42_imag = _RAND_17[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_45_real = _RAND_18[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_45_imag = _RAND_19[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_48_real = _RAND_20[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_48_imag = _RAND_21[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_51_real = _RAND_22[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_51_imag = _RAND_23[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_54_real = _RAND_24[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_54_imag = _RAND_25[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_57_real = _RAND_26[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T_57_imag = _RAND_27[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_60_real = _RAND_28[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_60_imag = _RAND_29[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_63_real = _RAND_30[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T_63_imag = _RAND_31[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _T_66_real = _RAND_32[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _T_66_imag = _RAND_33[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _T_69_real = _RAND_34[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _T_69_imag = _RAND_35[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _T_72_real = _RAND_36[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _T_72_imag = _RAND_37[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _T_75_real = _RAND_38[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _T_75_imag = _RAND_39[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _T_78_real = _RAND_40[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  _T_78_imag = _RAND_41[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  _T_81_real = _RAND_42[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  _T_81_imag = _RAND_43[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  _T_84_real = _RAND_44[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  _T_84_imag = _RAND_45[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  _T_87_real = _RAND_46[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  _T_87_imag = _RAND_47[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  _T_90_real = _RAND_48[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  _T_90_imag = _RAND_49[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  _T_93_real = _RAND_50[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  _T_93_imag = _RAND_51[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  _T_96_real = _RAND_52[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  _T_96_imag = _RAND_53[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  _T_99_real = _RAND_54[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  _T_99_imag = _RAND_55[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  _T_102_real = _RAND_56[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  _T_102_imag = _RAND_57[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  _T_105_real = _RAND_58[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  _T_105_imag = _RAND_59[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  _T_108_real = _RAND_60[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  _T_108_imag = _RAND_61[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  _T_111_real = _RAND_62[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  _T_111_imag = _RAND_63[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  feedback_real = _RAND_64[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  feedback_imag = _RAND_65[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  butt_out_0_real = _RAND_66[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  butt_out_0_imag = _RAND_67[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  load_output = _RAND_68[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (io_en) begin
      shift_out_real <= _T_111_real;
    end
    if (io_en) begin
      shift_out_imag <= _T_111_imag;
    end
    if (io_en) begin
      if (load_input) begin
        _T_21_real <= io_in_real;
      end else begin
        _T_21_real <= butterfly_outputs_1_real;
      end
    end
    if (io_en) begin
      if (load_input) begin
        _T_21_imag <= io_in_imag;
      end else begin
        _T_21_imag <= butterfly_outputs_1_imag;
      end
    end
    if (io_en) begin
      _T_24_real <= _T_21_real;
    end
    if (io_en) begin
      _T_24_imag <= _T_21_imag;
    end
    if (io_en) begin
      _T_27_real <= _T_24_real;
    end
    if (io_en) begin
      _T_27_imag <= _T_24_imag;
    end
    if (io_en) begin
      _T_30_real <= _T_27_real;
    end
    if (io_en) begin
      _T_30_imag <= _T_27_imag;
    end
    if (io_en) begin
      _T_33_real <= _T_30_real;
    end
    if (io_en) begin
      _T_33_imag <= _T_30_imag;
    end
    if (io_en) begin
      _T_36_real <= _T_33_real;
    end
    if (io_en) begin
      _T_36_imag <= _T_33_imag;
    end
    if (io_en) begin
      _T_39_real <= _T_36_real;
    end
    if (io_en) begin
      _T_39_imag <= _T_36_imag;
    end
    if (io_en) begin
      _T_42_real <= _T_39_real;
    end
    if (io_en) begin
      _T_42_imag <= _T_39_imag;
    end
    if (io_en) begin
      _T_45_real <= _T_42_real;
    end
    if (io_en) begin
      _T_45_imag <= _T_42_imag;
    end
    if (io_en) begin
      _T_48_real <= _T_45_real;
    end
    if (io_en) begin
      _T_48_imag <= _T_45_imag;
    end
    if (io_en) begin
      _T_51_real <= _T_48_real;
    end
    if (io_en) begin
      _T_51_imag <= _T_48_imag;
    end
    if (io_en) begin
      _T_54_real <= _T_51_real;
    end
    if (io_en) begin
      _T_54_imag <= _T_51_imag;
    end
    if (io_en) begin
      _T_57_real <= _T_54_real;
    end
    if (io_en) begin
      _T_57_imag <= _T_54_imag;
    end
    if (io_en) begin
      _T_60_real <= _T_57_real;
    end
    if (io_en) begin
      _T_60_imag <= _T_57_imag;
    end
    if (io_en) begin
      _T_63_real <= _T_60_real;
    end
    if (io_en) begin
      _T_63_imag <= _T_60_imag;
    end
    if (io_en) begin
      _T_66_real <= _T_63_real;
    end
    if (io_en) begin
      _T_66_imag <= _T_63_imag;
    end
    if (io_en) begin
      _T_69_real <= _T_66_real;
    end
    if (io_en) begin
      _T_69_imag <= _T_66_imag;
    end
    if (io_en) begin
      _T_72_real <= _T_69_real;
    end
    if (io_en) begin
      _T_72_imag <= _T_69_imag;
    end
    if (io_en) begin
      _T_75_real <= _T_72_real;
    end
    if (io_en) begin
      _T_75_imag <= _T_72_imag;
    end
    if (io_en) begin
      _T_78_real <= _T_75_real;
    end
    if (io_en) begin
      _T_78_imag <= _T_75_imag;
    end
    if (io_en) begin
      _T_81_real <= _T_78_real;
    end
    if (io_en) begin
      _T_81_imag <= _T_78_imag;
    end
    if (io_en) begin
      _T_84_real <= _T_81_real;
    end
    if (io_en) begin
      _T_84_imag <= _T_81_imag;
    end
    if (io_en) begin
      _T_87_real <= _T_84_real;
    end
    if (io_en) begin
      _T_87_imag <= _T_84_imag;
    end
    if (io_en) begin
      _T_90_real <= _T_87_real;
    end
    if (io_en) begin
      _T_90_imag <= _T_87_imag;
    end
    if (io_en) begin
      _T_93_real <= _T_90_real;
    end
    if (io_en) begin
      _T_93_imag <= _T_90_imag;
    end
    if (io_en) begin
      _T_96_real <= _T_93_real;
    end
    if (io_en) begin
      _T_96_imag <= _T_93_imag;
    end
    if (io_en) begin
      _T_99_real <= _T_96_real;
    end
    if (io_en) begin
      _T_99_imag <= _T_96_imag;
    end
    if (io_en) begin
      _T_102_real <= _T_99_real;
    end
    if (io_en) begin
      _T_102_imag <= _T_99_imag;
    end
    if (io_en) begin
      _T_105_real <= _T_102_real;
    end
    if (io_en) begin
      _T_105_imag <= _T_102_imag;
    end
    if (io_en) begin
      _T_108_real <= _T_105_real;
    end
    if (io_en) begin
      _T_108_imag <= _T_105_imag;
    end
    if (io_en) begin
      _T_111_real <= _T_108_real;
    end
    if (io_en) begin
      _T_111_imag <= _T_108_imag;
    end
    feedback_real <= shift_out_real;
    feedback_imag <= shift_out_imag;
    butt_out_0_real <= _T_128[16:1];
    butt_out_0_imag <= _T_135[16:1];
    if (reset) begin
      load_output <= 1'h0;
    end else begin
      load_output <= load_input;
    end
  end
endmodule
module SDFStageRadix22_2(
  input         clock,
  input         reset,
  input  [15:0] io_in_real,
  input  [15:0] io_in_imag,
  output [15:0] io_out_real,
  output [15:0] io_out_imag,
  input  [6:0]  io_cntr,
  input         io_en
);
  wire  load_input = io_cntr < 7'h10; // @[SDFChainRadix22.scala 426:66]
  reg [15:0] shift_out_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_0;
  wire [16:0] butt_outputs_1_real = $signed(shift_out_real) - $signed(io_in_real); // @[FixedPointTypeClass.scala 33:22]
  wire [17:0] _T_92 = {$signed(butt_outputs_1_real), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_94 = _T_92[17:1]; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_97 = $signed(_T_94) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] butterfly_outputs_1_real = _T_97[16:1]; // @[FixedPointTypeClass.scala 176:41]
  reg [15:0] shift_out_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1;
  wire [16:0] butt_outputs_1_imag = $signed(shift_out_imag) - $signed(io_in_imag); // @[FixedPointTypeClass.scala 33:22]
  wire [17:0] _T_99 = {$signed(butt_outputs_1_imag), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_101 = _T_99[17:1]; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_104 = $signed(_T_101) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] butterfly_outputs_1_imag = _T_104[16:1]; // @[FixedPointTypeClass.scala 176:41]
  reg [15:0] _T_21_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2;
  reg [15:0] _T_21_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3;
  reg [15:0] _T_24_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4;
  reg [15:0] _T_24_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5;
  reg [15:0] _T_27_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6;
  reg [15:0] _T_27_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7;
  reg [15:0] _T_30_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8;
  reg [15:0] _T_30_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9;
  reg [15:0] _T_33_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10;
  reg [15:0] _T_33_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11;
  reg [15:0] _T_36_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12;
  reg [15:0] _T_36_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_13;
  reg [15:0] _T_39_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_14;
  reg [15:0] _T_39_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_15;
  reg [15:0] _T_42_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_16;
  reg [15:0] _T_42_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_17;
  reg [15:0] _T_45_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_18;
  reg [15:0] _T_45_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_19;
  reg [15:0] _T_48_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_20;
  reg [15:0] _T_48_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_21;
  reg [15:0] _T_51_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_22;
  reg [15:0] _T_51_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_23;
  reg [15:0] _T_54_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_24;
  reg [15:0] _T_54_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_25;
  reg [15:0] _T_57_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_26;
  reg [15:0] _T_57_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_27;
  reg [15:0] _T_60_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_28;
  reg [15:0] _T_60_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_29;
  reg [15:0] _T_63_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_30;
  reg [15:0] _T_63_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_31;
  wire [16:0] butt_outputs_0_real = $signed(shift_out_real) + $signed(io_in_real); // @[FixedPointTypeClass.scala 24:22]
  wire [16:0] butt_outputs_0_imag = $signed(shift_out_imag) + $signed(io_in_imag); // @[FixedPointTypeClass.scala 24:22]
  wire [17:0] _T_75 = {$signed(butt_outputs_0_real), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_77 = _T_75[17:1]; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_80 = $signed(_T_77) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  wire [17:0] _T_82 = {$signed(butt_outputs_0_imag), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_84 = _T_82[17:1]; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_87 = $signed(_T_84) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  reg [15:0] feedback_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_32;
  reg [15:0] feedback_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_33;
  reg [15:0] butt_out_0_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_34;
  reg [15:0] butt_out_0_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_35;
  reg  load_output; // @[Reg.scala 27:20]
  reg [31:0] _RAND_36;
  assign io_out_real = load_output ? $signed(feedback_real) : $signed(butt_out_0_real); // @[SDFChainRadix22.scala 422:10]
  assign io_out_imag = load_output ? $signed(feedback_imag) : $signed(butt_out_0_imag); // @[SDFChainRadix22.scala 422:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  shift_out_real = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  shift_out_imag = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_21_real = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_21_imag = _RAND_3[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_24_real = _RAND_4[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_24_imag = _RAND_5[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_27_real = _RAND_6[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_27_imag = _RAND_7[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_30_real = _RAND_8[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_30_imag = _RAND_9[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_33_real = _RAND_10[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_33_imag = _RAND_11[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_36_real = _RAND_12[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_36_imag = _RAND_13[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_39_real = _RAND_14[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_39_imag = _RAND_15[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_42_real = _RAND_16[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_42_imag = _RAND_17[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_45_real = _RAND_18[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_45_imag = _RAND_19[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_48_real = _RAND_20[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_48_imag = _RAND_21[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_51_real = _RAND_22[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_51_imag = _RAND_23[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_54_real = _RAND_24[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_54_imag = _RAND_25[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_57_real = _RAND_26[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T_57_imag = _RAND_27[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_60_real = _RAND_28[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_60_imag = _RAND_29[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_63_real = _RAND_30[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T_63_imag = _RAND_31[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  feedback_real = _RAND_32[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  feedback_imag = _RAND_33[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  butt_out_0_real = _RAND_34[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  butt_out_0_imag = _RAND_35[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  load_output = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (io_en) begin
      shift_out_real <= _T_63_real;
    end
    if (io_en) begin
      shift_out_imag <= _T_63_imag;
    end
    if (io_en) begin
      if (load_input) begin
        _T_21_real <= io_in_real;
      end else begin
        _T_21_real <= butterfly_outputs_1_real;
      end
    end
    if (io_en) begin
      if (load_input) begin
        _T_21_imag <= io_in_imag;
      end else begin
        _T_21_imag <= butterfly_outputs_1_imag;
      end
    end
    if (io_en) begin
      _T_24_real <= _T_21_real;
    end
    if (io_en) begin
      _T_24_imag <= _T_21_imag;
    end
    if (io_en) begin
      _T_27_real <= _T_24_real;
    end
    if (io_en) begin
      _T_27_imag <= _T_24_imag;
    end
    if (io_en) begin
      _T_30_real <= _T_27_real;
    end
    if (io_en) begin
      _T_30_imag <= _T_27_imag;
    end
    if (io_en) begin
      _T_33_real <= _T_30_real;
    end
    if (io_en) begin
      _T_33_imag <= _T_30_imag;
    end
    if (io_en) begin
      _T_36_real <= _T_33_real;
    end
    if (io_en) begin
      _T_36_imag <= _T_33_imag;
    end
    if (io_en) begin
      _T_39_real <= _T_36_real;
    end
    if (io_en) begin
      _T_39_imag <= _T_36_imag;
    end
    if (io_en) begin
      _T_42_real <= _T_39_real;
    end
    if (io_en) begin
      _T_42_imag <= _T_39_imag;
    end
    if (io_en) begin
      _T_45_real <= _T_42_real;
    end
    if (io_en) begin
      _T_45_imag <= _T_42_imag;
    end
    if (io_en) begin
      _T_48_real <= _T_45_real;
    end
    if (io_en) begin
      _T_48_imag <= _T_45_imag;
    end
    if (io_en) begin
      _T_51_real <= _T_48_real;
    end
    if (io_en) begin
      _T_51_imag <= _T_48_imag;
    end
    if (io_en) begin
      _T_54_real <= _T_51_real;
    end
    if (io_en) begin
      _T_54_imag <= _T_51_imag;
    end
    if (io_en) begin
      _T_57_real <= _T_54_real;
    end
    if (io_en) begin
      _T_57_imag <= _T_54_imag;
    end
    if (io_en) begin
      _T_60_real <= _T_57_real;
    end
    if (io_en) begin
      _T_60_imag <= _T_57_imag;
    end
    if (io_en) begin
      _T_63_real <= _T_60_real;
    end
    if (io_en) begin
      _T_63_imag <= _T_60_imag;
    end
    feedback_real <= shift_out_real;
    feedback_imag <= shift_out_imag;
    butt_out_0_real <= _T_80[16:1];
    butt_out_0_imag <= _T_87[16:1];
    if (reset) begin
      load_output <= 1'h0;
    end else begin
      load_output <= load_input;
    end
  end
endmodule
module SDFStageRadix22_3(
  input         clock,
  input         reset,
  input  [15:0] io_in_real,
  input  [15:0] io_in_imag,
  output [15:0] io_out_real,
  output [15:0] io_out_imag,
  input  [6:0]  io_cntr,
  input         io_en
);
  wire  load_input = io_cntr < 7'h8; // @[SDFChainRadix22.scala 426:66]
  reg [15:0] shift_out_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_0;
  wire [16:0] butt_outputs_1_real = $signed(shift_out_real) - $signed(io_in_real); // @[FixedPointTypeClass.scala 33:22]
  wire [17:0] _T_68 = {$signed(butt_outputs_1_real), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_70 = _T_68[17:1]; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_73 = $signed(_T_70) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] butterfly_outputs_1_real = _T_73[16:1]; // @[FixedPointTypeClass.scala 176:41]
  reg [15:0] shift_out_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1;
  wire [16:0] butt_outputs_1_imag = $signed(shift_out_imag) - $signed(io_in_imag); // @[FixedPointTypeClass.scala 33:22]
  wire [17:0] _T_75 = {$signed(butt_outputs_1_imag), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_77 = _T_75[17:1]; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_80 = $signed(_T_77) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] butterfly_outputs_1_imag = _T_80[16:1]; // @[FixedPointTypeClass.scala 176:41]
  reg [15:0] _T_21_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2;
  reg [15:0] _T_21_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3;
  reg [15:0] _T_24_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4;
  reg [15:0] _T_24_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5;
  reg [15:0] _T_27_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6;
  reg [15:0] _T_27_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7;
  reg [15:0] _T_30_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8;
  reg [15:0] _T_30_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9;
  reg [15:0] _T_33_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10;
  reg [15:0] _T_33_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11;
  reg [15:0] _T_36_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12;
  reg [15:0] _T_36_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_13;
  reg [15:0] _T_39_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_14;
  reg [15:0] _T_39_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_15;
  wire [16:0] butt_outputs_0_real = $signed(shift_out_real) + $signed(io_in_real); // @[FixedPointTypeClass.scala 24:22]
  wire [16:0] butt_outputs_0_imag = $signed(shift_out_imag) + $signed(io_in_imag); // @[FixedPointTypeClass.scala 24:22]
  wire [17:0] _T_51 = {$signed(butt_outputs_0_real), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_53 = _T_51[17:1]; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_56 = $signed(_T_53) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  wire [17:0] _T_58 = {$signed(butt_outputs_0_imag), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_60 = _T_58[17:1]; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_63 = $signed(_T_60) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  reg [15:0] feedback_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_16;
  reg [15:0] feedback_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_17;
  reg [15:0] butt_out_0_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_18;
  reg [15:0] butt_out_0_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_19;
  reg  load_output; // @[Reg.scala 27:20]
  reg [31:0] _RAND_20;
  assign io_out_real = load_output ? $signed(feedback_real) : $signed(butt_out_0_real); // @[SDFChainRadix22.scala 422:10]
  assign io_out_imag = load_output ? $signed(feedback_imag) : $signed(butt_out_0_imag); // @[SDFChainRadix22.scala 422:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  shift_out_real = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  shift_out_imag = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_21_real = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_21_imag = _RAND_3[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_24_real = _RAND_4[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_24_imag = _RAND_5[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_27_real = _RAND_6[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_27_imag = _RAND_7[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_30_real = _RAND_8[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_30_imag = _RAND_9[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_33_real = _RAND_10[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_33_imag = _RAND_11[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_36_real = _RAND_12[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_36_imag = _RAND_13[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_39_real = _RAND_14[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_39_imag = _RAND_15[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  feedback_real = _RAND_16[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  feedback_imag = _RAND_17[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  butt_out_0_real = _RAND_18[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  butt_out_0_imag = _RAND_19[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  load_output = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (io_en) begin
      shift_out_real <= _T_39_real;
    end
    if (io_en) begin
      shift_out_imag <= _T_39_imag;
    end
    if (io_en) begin
      if (load_input) begin
        _T_21_real <= io_in_real;
      end else begin
        _T_21_real <= butterfly_outputs_1_real;
      end
    end
    if (io_en) begin
      if (load_input) begin
        _T_21_imag <= io_in_imag;
      end else begin
        _T_21_imag <= butterfly_outputs_1_imag;
      end
    end
    if (io_en) begin
      _T_24_real <= _T_21_real;
    end
    if (io_en) begin
      _T_24_imag <= _T_21_imag;
    end
    if (io_en) begin
      _T_27_real <= _T_24_real;
    end
    if (io_en) begin
      _T_27_imag <= _T_24_imag;
    end
    if (io_en) begin
      _T_30_real <= _T_27_real;
    end
    if (io_en) begin
      _T_30_imag <= _T_27_imag;
    end
    if (io_en) begin
      _T_33_real <= _T_30_real;
    end
    if (io_en) begin
      _T_33_imag <= _T_30_imag;
    end
    if (io_en) begin
      _T_36_real <= _T_33_real;
    end
    if (io_en) begin
      _T_36_imag <= _T_33_imag;
    end
    if (io_en) begin
      _T_39_real <= _T_36_real;
    end
    if (io_en) begin
      _T_39_imag <= _T_36_imag;
    end
    feedback_real <= shift_out_real;
    feedback_imag <= shift_out_imag;
    butt_out_0_real <= _T_56[16:1];
    butt_out_0_imag <= _T_63[16:1];
    if (reset) begin
      load_output <= 1'h0;
    end else begin
      load_output <= load_input;
    end
  end
endmodule
module SDFStageRadix22_4(
  input         clock,
  input         reset,
  input  [15:0] io_in_real,
  input  [15:0] io_in_imag,
  output [15:0] io_out_real,
  output [15:0] io_out_imag,
  input  [6:0]  io_cntr,
  input         io_en
);
  wire  load_input = io_cntr < 7'h4; // @[SDFChainRadix22.scala 426:66]
  reg [15:0] shift_out_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_0;
  wire [16:0] butt_outputs_1_real = $signed(shift_out_real) - $signed(io_in_real); // @[FixedPointTypeClass.scala 33:22]
  wire [17:0] _T_56 = {$signed(butt_outputs_1_real), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_58 = _T_56[17:1]; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_61 = $signed(_T_58) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] butterfly_outputs_1_real = _T_61[16:1]; // @[FixedPointTypeClass.scala 176:41]
  reg [15:0] shift_out_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1;
  wire [16:0] butt_outputs_1_imag = $signed(shift_out_imag) - $signed(io_in_imag); // @[FixedPointTypeClass.scala 33:22]
  wire [17:0] _T_63 = {$signed(butt_outputs_1_imag), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_65 = _T_63[17:1]; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_68 = $signed(_T_65) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] butterfly_outputs_1_imag = _T_68[16:1]; // @[FixedPointTypeClass.scala 176:41]
  reg [15:0] _T_21_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2;
  reg [15:0] _T_21_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3;
  reg [15:0] _T_24_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4;
  reg [15:0] _T_24_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5;
  reg [15:0] _T_27_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6;
  reg [15:0] _T_27_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7;
  wire [16:0] butt_outputs_0_real = $signed(shift_out_real) + $signed(io_in_real); // @[FixedPointTypeClass.scala 24:22]
  wire [16:0] butt_outputs_0_imag = $signed(shift_out_imag) + $signed(io_in_imag); // @[FixedPointTypeClass.scala 24:22]
  wire [17:0] _T_39 = {$signed(butt_outputs_0_real), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_41 = _T_39[17:1]; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_44 = $signed(_T_41) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  wire [17:0] _T_46 = {$signed(butt_outputs_0_imag), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_48 = _T_46[17:1]; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_51 = $signed(_T_48) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  reg [15:0] feedback_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8;
  reg [15:0] feedback_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9;
  reg [15:0] butt_out_0_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10;
  reg [15:0] butt_out_0_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11;
  reg  load_output; // @[Reg.scala 27:20]
  reg [31:0] _RAND_12;
  assign io_out_real = load_output ? $signed(feedback_real) : $signed(butt_out_0_real); // @[SDFChainRadix22.scala 422:10]
  assign io_out_imag = load_output ? $signed(feedback_imag) : $signed(butt_out_0_imag); // @[SDFChainRadix22.scala 422:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  shift_out_real = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  shift_out_imag = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_21_real = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_21_imag = _RAND_3[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_24_real = _RAND_4[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_24_imag = _RAND_5[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_27_real = _RAND_6[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_27_imag = _RAND_7[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  feedback_real = _RAND_8[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  feedback_imag = _RAND_9[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  butt_out_0_real = _RAND_10[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  butt_out_0_imag = _RAND_11[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  load_output = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (io_en) begin
      shift_out_real <= _T_27_real;
    end
    if (io_en) begin
      shift_out_imag <= _T_27_imag;
    end
    if (io_en) begin
      if (load_input) begin
        _T_21_real <= io_in_real;
      end else begin
        _T_21_real <= butterfly_outputs_1_real;
      end
    end
    if (io_en) begin
      if (load_input) begin
        _T_21_imag <= io_in_imag;
      end else begin
        _T_21_imag <= butterfly_outputs_1_imag;
      end
    end
    if (io_en) begin
      _T_24_real <= _T_21_real;
    end
    if (io_en) begin
      _T_24_imag <= _T_21_imag;
    end
    if (io_en) begin
      _T_27_real <= _T_24_real;
    end
    if (io_en) begin
      _T_27_imag <= _T_24_imag;
    end
    feedback_real <= shift_out_real;
    feedback_imag <= shift_out_imag;
    butt_out_0_real <= _T_44[16:1];
    butt_out_0_imag <= _T_51[16:1];
    if (reset) begin
      load_output <= 1'h0;
    end else begin
      load_output <= load_input;
    end
  end
endmodule
module SDFStageRadix22_5(
  input         clock,
  input         reset,
  input  [15:0] io_in_real,
  input  [15:0] io_in_imag,
  output [15:0] io_out_real,
  output [15:0] io_out_imag,
  input  [6:0]  io_cntr,
  input         io_en
);
  wire  load_input = io_cntr < 7'h2; // @[SDFChainRadix22.scala 426:66]
  reg [15:0] shift_out_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_0;
  wire [16:0] butt_outputs_1_real = $signed(shift_out_real) - $signed(io_in_real); // @[FixedPointTypeClass.scala 33:22]
  wire [17:0] _T_50 = {$signed(butt_outputs_1_real), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_52 = _T_50[17:1]; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_55 = $signed(_T_52) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] butterfly_outputs_1_real = _T_55[16:1]; // @[FixedPointTypeClass.scala 176:41]
  reg [15:0] shift_out_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1;
  wire [16:0] butt_outputs_1_imag = $signed(shift_out_imag) - $signed(io_in_imag); // @[FixedPointTypeClass.scala 33:22]
  wire [17:0] _T_57 = {$signed(butt_outputs_1_imag), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_59 = _T_57[17:1]; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_62 = $signed(_T_59) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] butterfly_outputs_1_imag = _T_62[16:1]; // @[FixedPointTypeClass.scala 176:41]
  reg [15:0] _T_21_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2;
  reg [15:0] _T_21_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3;
  wire [16:0] butt_outputs_0_real = $signed(shift_out_real) + $signed(io_in_real); // @[FixedPointTypeClass.scala 24:22]
  wire [16:0] butt_outputs_0_imag = $signed(shift_out_imag) + $signed(io_in_imag); // @[FixedPointTypeClass.scala 24:22]
  wire [17:0] _T_33 = {$signed(butt_outputs_0_real), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_35 = _T_33[17:1]; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_38 = $signed(_T_35) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  wire [17:0] _T_40 = {$signed(butt_outputs_0_imag), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_42 = _T_40[17:1]; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_45 = $signed(_T_42) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  reg [15:0] feedback_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4;
  reg [15:0] feedback_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5;
  reg [15:0] butt_out_0_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6;
  reg [15:0] butt_out_0_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7;
  reg  load_output; // @[Reg.scala 27:20]
  reg [31:0] _RAND_8;
  assign io_out_real = load_output ? $signed(feedback_real) : $signed(butt_out_0_real); // @[SDFChainRadix22.scala 422:10]
  assign io_out_imag = load_output ? $signed(feedback_imag) : $signed(butt_out_0_imag); // @[SDFChainRadix22.scala 422:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  shift_out_real = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  shift_out_imag = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_21_real = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_21_imag = _RAND_3[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  feedback_real = _RAND_4[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  feedback_imag = _RAND_5[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  butt_out_0_real = _RAND_6[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  butt_out_0_imag = _RAND_7[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  load_output = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (io_en) begin
      shift_out_real <= _T_21_real;
    end
    if (io_en) begin
      shift_out_imag <= _T_21_imag;
    end
    if (io_en) begin
      if (load_input) begin
        _T_21_real <= io_in_real;
      end else begin
        _T_21_real <= butterfly_outputs_1_real;
      end
    end
    if (io_en) begin
      if (load_input) begin
        _T_21_imag <= io_in_imag;
      end else begin
        _T_21_imag <= butterfly_outputs_1_imag;
      end
    end
    feedback_real <= shift_out_real;
    feedback_imag <= shift_out_imag;
    butt_out_0_real <= _T_38[16:1];
    butt_out_0_imag <= _T_45[16:1];
    if (reset) begin
      load_output <= 1'h0;
    end else begin
      load_output <= load_input;
    end
  end
endmodule
module SDFStageRadix22_6(
  input         clock,
  input         reset,
  input  [15:0] io_in_real,
  input  [15:0] io_in_imag,
  output [15:0] io_out_real,
  output [15:0] io_out_imag,
  input  [6:0]  io_cntr,
  input         io_en
);
  wire  load_input = io_cntr < 7'h1; // @[SDFChainRadix22.scala 426:66]
  reg [15:0] shift_out_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_0;
  wire [16:0] butt_outputs_1_real = $signed(shift_out_real) - $signed(io_in_real); // @[FixedPointTypeClass.scala 33:22]
  wire [17:0] _T_47 = {$signed(butt_outputs_1_real), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_49 = _T_47[17:1]; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_52 = $signed(_T_49) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] butterfly_outputs_1_real = _T_52[16:1]; // @[FixedPointTypeClass.scala 176:41]
  reg [15:0] shift_out_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1;
  wire [16:0] butt_outputs_1_imag = $signed(shift_out_imag) - $signed(io_in_imag); // @[FixedPointTypeClass.scala 33:22]
  wire [17:0] _T_54 = {$signed(butt_outputs_1_imag), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_56 = _T_54[17:1]; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_59 = $signed(_T_56) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  wire [15:0] butterfly_outputs_1_imag = _T_59[16:1]; // @[FixedPointTypeClass.scala 176:41]
  wire [16:0] butt_outputs_0_real = $signed(shift_out_real) + $signed(io_in_real); // @[FixedPointTypeClass.scala 24:22]
  wire [16:0] butt_outputs_0_imag = $signed(shift_out_imag) + $signed(io_in_imag); // @[FixedPointTypeClass.scala 24:22]
  wire [17:0] _T_30 = {$signed(butt_outputs_0_real), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_32 = _T_30[17:1]; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_35 = $signed(_T_32) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  wire [17:0] _T_37 = {$signed(butt_outputs_0_imag), 1'h0}; // @[FixedPointTypeClass.scala 129:22 FixedPointTypeClass.scala 130:12]
  wire [16:0] _T_39 = _T_37[17:1]; // @[FixedPointTypeClass.scala 133:23]
  wire [16:0] _T_42 = $signed(_T_39) + 17'sh1; // @[FixedPointTypeClass.scala 20:58]
  reg [15:0] feedback_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2;
  reg [15:0] feedback_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3;
  reg [15:0] butt_out_0_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4;
  reg [15:0] butt_out_0_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5;
  reg  load_output; // @[Reg.scala 27:20]
  reg [31:0] _RAND_6;
  assign io_out_real = load_output ? $signed(feedback_real) : $signed(butt_out_0_real); // @[SDFChainRadix22.scala 422:10]
  assign io_out_imag = load_output ? $signed(feedback_imag) : $signed(butt_out_0_imag); // @[SDFChainRadix22.scala 422:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  shift_out_real = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  shift_out_imag = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  feedback_real = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  feedback_imag = _RAND_3[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  butt_out_0_real = _RAND_4[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  butt_out_0_imag = _RAND_5[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  load_output = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (io_en) begin
      if (load_input) begin
        shift_out_real <= io_in_real;
      end else begin
        shift_out_real <= butterfly_outputs_1_real;
      end
    end
    if (io_en) begin
      if (load_input) begin
        shift_out_imag <= io_in_imag;
      end else begin
        shift_out_imag <= butterfly_outputs_1_imag;
      end
    end
    feedback_real <= shift_out_real;
    feedback_imag <= shift_out_imag;
    butt_out_0_real <= _T_35[16:1];
    butt_out_0_imag <= _T_42[16:1];
    if (reset) begin
      load_output <= 1'h0;
    end else begin
      load_output <= load_input;
    end
  end
endmodule
module Queue_10(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [15:0] io_enq_bits_real,
  input  [15:0] io_enq_bits_imag,
  input         io_deq_ready,
  output        io_deq_valid,
  output [15:0] io_deq_bits_real,
  output [15:0] io_deq_bits_imag
);
  reg [15:0] _T_4_real [0:28]; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_0;
  wire [15:0] _T_4_real__T_26_data; // @[Decoupled.scala 218:24]
  wire [4:0] _T_4_real__T_26_addr; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_1;
  wire [15:0] _T_4_real__T_16_data; // @[Decoupled.scala 218:24]
  wire [4:0] _T_4_real__T_16_addr; // @[Decoupled.scala 218:24]
  wire  _T_4_real__T_16_mask; // @[Decoupled.scala 218:24]
  wire  _T_4_real__T_16_en; // @[Decoupled.scala 218:24]
  reg [15:0] _T_4_imag [0:28]; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_2;
  wire [15:0] _T_4_imag__T_26_data; // @[Decoupled.scala 218:24]
  wire [4:0] _T_4_imag__T_26_addr; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_3;
  wire [15:0] _T_4_imag__T_16_data; // @[Decoupled.scala 218:24]
  wire [4:0] _T_4_imag__T_16_addr; // @[Decoupled.scala 218:24]
  wire  _T_4_imag__T_16_mask; // @[Decoupled.scala 218:24]
  wire  _T_4_imag__T_16_en; // @[Decoupled.scala 218:24]
  reg [4:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_4;
  reg [4:0] value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  reg  _T_5; // @[Decoupled.scala 221:35]
  reg [31:0] _RAND_6;
  wire  _T_6 = value == value_1; // @[Decoupled.scala 223:41]
  wire  _T_7 = ~_T_5; // @[Decoupled.scala 224:36]
  wire  _T_8 = _T_6 & _T_7; // @[Decoupled.scala 224:33]
  wire  _T_9 = _T_6 & _T_5; // @[Decoupled.scala 225:32]
  wire  _T_10 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  _T_12 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire  wrap = value == 5'h1c; // @[Counter.scala 38:24]
  wire [4:0] _T_18 = value + 5'h1; // @[Counter.scala 39:22]
  wire  _GEN_12 = io_deq_ready ? 1'h0 : _T_10; // @[Decoupled.scala 249:27]
  wire  _GEN_16 = _T_8 ? _GEN_12 : _T_10; // @[Decoupled.scala 246:18]
  wire  wrap_1 = value_1 == 5'h1c; // @[Counter.scala 38:24]
  wire [4:0] _T_20 = value_1 + 5'h1; // @[Counter.scala 39:22]
  wire  _GEN_15 = _T_8 ? 1'h0 : _T_12; // @[Decoupled.scala 246:18]
  wire  _T_21 = _GEN_16 != _GEN_15; // @[Decoupled.scala 236:16]
  wire  _T_22 = ~_T_8; // @[Decoupled.scala 240:19]
  wire  _T_23 = ~_T_9; // @[Decoupled.scala 241:19]
  assign _T_4_real__T_26_addr = value_1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_4_real__T_26_data = _T_4_real[_T_4_real__T_26_addr]; // @[Decoupled.scala 218:24]
  `else
  assign _T_4_real__T_26_data = _T_4_real__T_26_addr >= 5'h1d ? _RAND_1[15:0] : _T_4_real[_T_4_real__T_26_addr]; // @[Decoupled.scala 218:24]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_4_real__T_16_data = io_enq_bits_real;
  assign _T_4_real__T_16_addr = value;
  assign _T_4_real__T_16_mask = 1'h1;
  assign _T_4_real__T_16_en = _T_8 ? _GEN_12 : _T_10;
  assign _T_4_imag__T_26_addr = value_1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_4_imag__T_26_data = _T_4_imag[_T_4_imag__T_26_addr]; // @[Decoupled.scala 218:24]
  `else
  assign _T_4_imag__T_26_data = _T_4_imag__T_26_addr >= 5'h1d ? _RAND_3[15:0] : _T_4_imag[_T_4_imag__T_26_addr]; // @[Decoupled.scala 218:24]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_4_imag__T_16_data = io_enq_bits_imag;
  assign _T_4_imag__T_16_addr = value;
  assign _T_4_imag__T_16_mask = 1'h1;
  assign _T_4_imag__T_16_en = _T_8 ? _GEN_12 : _T_10;
  assign io_enq_ready = io_deq_ready | _T_23; // @[Decoupled.scala 241:16 Decoupled.scala 254:40]
  assign io_deq_valid = io_enq_valid | _T_22; // @[Decoupled.scala 240:16 Decoupled.scala 245:40]
  assign io_deq_bits_real = _T_8 ? $signed(io_enq_bits_real) : $signed(_T_4_real__T_26_data); // @[Decoupled.scala 242:15 Decoupled.scala 247:19]
  assign io_deq_bits_imag = _T_8 ? $signed(io_enq_bits_imag) : $signed(_T_4_imag__T_26_data); // @[Decoupled.scala 242:15 Decoupled.scala 247:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 29; initvar = initvar+1)
    _T_4_real[initvar] = _RAND_0[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  _RAND_2 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 29; initvar = initvar+1)
    _T_4_imag[initvar] = _RAND_2[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  value = _RAND_4[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value_1 = _RAND_5[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_5 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T_4_real__T_16_en & _T_4_real__T_16_mask) begin
      _T_4_real[_T_4_real__T_16_addr] <= _T_4_real__T_16_data; // @[Decoupled.scala 218:24]
    end
    if(_T_4_imag__T_16_en & _T_4_imag__T_16_mask) begin
      _T_4_imag[_T_4_imag__T_16_addr] <= _T_4_imag__T_16_data; // @[Decoupled.scala 218:24]
    end
    if (reset) begin
      value <= 5'h0;
    end else if (_GEN_16) begin
      if (wrap) begin
        value <= 5'h0;
      end else begin
        value <= _T_18;
      end
    end
    if (reset) begin
      value_1 <= 5'h0;
    end else if (_GEN_15) begin
      if (wrap_1) begin
        value_1 <= 5'h0;
      end else begin
        value_1 <= _T_20;
      end
    end
    if (reset) begin
      _T_5 <= 1'h0;
    end else if (_T_21) begin
      if (_T_8) begin
        if (io_deq_ready) begin
          _T_5 <= 1'h0;
        end else begin
          _T_5 <= _T_10;
        end
      end else begin
        _T_5 <= _T_10;
      end
    end
  end
endmodule
module SDFChainRadix22(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [15:0] io_in_bits_real,
  input  [15:0] io_in_bits_imag,
  input         io_out_ready,
  output        io_out_valid,
  output [15:0] io_out_bits_real,
  output [15:0] io_out_bits_imag,
  output        io_lastOut,
  input         io_lastIn,
  input  [6:0]  io_fftSize,
  output        io_busy
);
  wire  sdf_stages_0_clock; // @[SDFChainRadix22.scala 155:25]
  wire  sdf_stages_0_reset; // @[SDFChainRadix22.scala 155:25]
  wire [15:0] sdf_stages_0_io_in_real; // @[SDFChainRadix22.scala 155:25]
  wire [15:0] sdf_stages_0_io_in_imag; // @[SDFChainRadix22.scala 155:25]
  wire [15:0] sdf_stages_0_io_out_real; // @[SDFChainRadix22.scala 155:25]
  wire [15:0] sdf_stages_0_io_out_imag; // @[SDFChainRadix22.scala 155:25]
  wire [6:0] sdf_stages_0_io_cntr; // @[SDFChainRadix22.scala 155:25]
  wire  sdf_stages_0_io_en; // @[SDFChainRadix22.scala 155:25]
  wire  sdf_stages_1_clock; // @[SDFChainRadix22.scala 155:25]
  wire  sdf_stages_1_reset; // @[SDFChainRadix22.scala 155:25]
  wire [15:0] sdf_stages_1_io_in_real; // @[SDFChainRadix22.scala 155:25]
  wire [15:0] sdf_stages_1_io_in_imag; // @[SDFChainRadix22.scala 155:25]
  wire [15:0] sdf_stages_1_io_out_real; // @[SDFChainRadix22.scala 155:25]
  wire [15:0] sdf_stages_1_io_out_imag; // @[SDFChainRadix22.scala 155:25]
  wire [6:0] sdf_stages_1_io_cntr; // @[SDFChainRadix22.scala 155:25]
  wire  sdf_stages_1_io_en; // @[SDFChainRadix22.scala 155:25]
  wire  sdf_stages_2_clock; // @[SDFChainRadix22.scala 155:25]
  wire  sdf_stages_2_reset; // @[SDFChainRadix22.scala 155:25]
  wire [15:0] sdf_stages_2_io_in_real; // @[SDFChainRadix22.scala 155:25]
  wire [15:0] sdf_stages_2_io_in_imag; // @[SDFChainRadix22.scala 155:25]
  wire [15:0] sdf_stages_2_io_out_real; // @[SDFChainRadix22.scala 155:25]
  wire [15:0] sdf_stages_2_io_out_imag; // @[SDFChainRadix22.scala 155:25]
  wire [6:0] sdf_stages_2_io_cntr; // @[SDFChainRadix22.scala 155:25]
  wire  sdf_stages_2_io_en; // @[SDFChainRadix22.scala 155:25]
  wire  sdf_stages_3_clock; // @[SDFChainRadix22.scala 155:25]
  wire  sdf_stages_3_reset; // @[SDFChainRadix22.scala 155:25]
  wire [15:0] sdf_stages_3_io_in_real; // @[SDFChainRadix22.scala 155:25]
  wire [15:0] sdf_stages_3_io_in_imag; // @[SDFChainRadix22.scala 155:25]
  wire [15:0] sdf_stages_3_io_out_real; // @[SDFChainRadix22.scala 155:25]
  wire [15:0] sdf_stages_3_io_out_imag; // @[SDFChainRadix22.scala 155:25]
  wire [6:0] sdf_stages_3_io_cntr; // @[SDFChainRadix22.scala 155:25]
  wire  sdf_stages_3_io_en; // @[SDFChainRadix22.scala 155:25]
  wire  sdf_stages_4_clock; // @[SDFChainRadix22.scala 155:25]
  wire  sdf_stages_4_reset; // @[SDFChainRadix22.scala 155:25]
  wire [15:0] sdf_stages_4_io_in_real; // @[SDFChainRadix22.scala 155:25]
  wire [15:0] sdf_stages_4_io_in_imag; // @[SDFChainRadix22.scala 155:25]
  wire [15:0] sdf_stages_4_io_out_real; // @[SDFChainRadix22.scala 155:25]
  wire [15:0] sdf_stages_4_io_out_imag; // @[SDFChainRadix22.scala 155:25]
  wire [6:0] sdf_stages_4_io_cntr; // @[SDFChainRadix22.scala 155:25]
  wire  sdf_stages_4_io_en; // @[SDFChainRadix22.scala 155:25]
  wire  sdf_stages_5_clock; // @[SDFChainRadix22.scala 155:25]
  wire  sdf_stages_5_reset; // @[SDFChainRadix22.scala 155:25]
  wire [15:0] sdf_stages_5_io_in_real; // @[SDFChainRadix22.scala 155:25]
  wire [15:0] sdf_stages_5_io_in_imag; // @[SDFChainRadix22.scala 155:25]
  wire [15:0] sdf_stages_5_io_out_real; // @[SDFChainRadix22.scala 155:25]
  wire [15:0] sdf_stages_5_io_out_imag; // @[SDFChainRadix22.scala 155:25]
  wire [6:0] sdf_stages_5_io_cntr; // @[SDFChainRadix22.scala 155:25]
  wire  sdf_stages_5_io_en; // @[SDFChainRadix22.scala 155:25]
  wire  sdf_stages_6_clock; // @[SDFChainRadix22.scala 155:25]
  wire  sdf_stages_6_reset; // @[SDFChainRadix22.scala 155:25]
  wire [15:0] sdf_stages_6_io_in_real; // @[SDFChainRadix22.scala 155:25]
  wire [15:0] sdf_stages_6_io_in_imag; // @[SDFChainRadix22.scala 155:25]
  wire [15:0] sdf_stages_6_io_out_real; // @[SDFChainRadix22.scala 155:25]
  wire [15:0] sdf_stages_6_io_out_imag; // @[SDFChainRadix22.scala 155:25]
  wire [6:0] sdf_stages_6_io_cntr; // @[SDFChainRadix22.scala 155:25]
  wire  sdf_stages_6_io_en; // @[SDFChainRadix22.scala 155:25]
  wire  outQueue_clock; // @[SDFChainRadix22.scala 356:25]
  wire  outQueue_reset; // @[SDFChainRadix22.scala 356:25]
  wire  outQueue_io_enq_ready; // @[SDFChainRadix22.scala 356:25]
  wire  outQueue_io_enq_valid; // @[SDFChainRadix22.scala 356:25]
  wire [15:0] outQueue_io_enq_bits_real; // @[SDFChainRadix22.scala 356:25]
  wire [15:0] outQueue_io_enq_bits_imag; // @[SDFChainRadix22.scala 356:25]
  wire  outQueue_io_deq_ready; // @[SDFChainRadix22.scala 356:25]
  wire  outQueue_io_deq_valid; // @[SDFChainRadix22.scala 356:25]
  wire [15:0] outQueue_io_deq_bits_real; // @[SDFChainRadix22.scala 356:25]
  wire [15:0] outQueue_io_deq_bits_imag; // @[SDFChainRadix22.scala 356:25]
  reg [6:0] regNumStages; // @[SDFChainRadix22.scala 41:29]
  reg [31:0] _RAND_0;
  reg [1:0] state; // @[SDFChainRadix22.scala 52:22]
  reg [31:0] _RAND_1;
  reg  initialOutDone; // @[SDFChainRadix22.scala 55:31]
  reg [31:0] _RAND_2;
  reg [7:0] cnt; // @[SDFChainRadix22.scala 56:20]
  reg [31:0] _RAND_3;
  wire [6:0] _T_39 = regNumStages - 7'h1; // @[SDFChainRadix22.scala 69:39]
  wire [128:0] _T_40 = 129'h2 << _T_39; // @[SDFChainRadix22.scala 69:23]
  wire  _T_41 = io_in_ready & io_in_valid; // @[Decoupled.scala 40:37]
  wire  fireLast = io_lastIn & _T_41; // @[SDFChainRadix22.scala 75:28]
  wire  _T_42 = 2'h0 == state; // @[Conditional.scala 37:30]
  wire [1:0] _GEN_0 = _T_41 ? 2'h1 : state; // @[SDFChainRadix22.scala 82:27]
  wire  _T_45 = 2'h1 == state; // @[Conditional.scala 37:30]
  wire [1:0] _GEN_1 = fireLast ? 2'h2 : state; // @[SDFChainRadix22.scala 85:23]
  wire  _T_46 = 2'h2 == state; // @[Conditional.scala 37:30]
  wire [1:0] _GEN_2 = io_lastOut ? 2'h0 : state; // @[SDFChainRadix22.scala 90:25]
  wire [1:0] _GEN_3 = _T_46 ? _GEN_2 : state; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_4 = _T_45 ? _GEN_1 : _GEN_3; // @[Conditional.scala 39:67]
  wire [1:0] state_next = _T_42 ? _GEN_0 : _GEN_4; // @[Conditional.scala 40:58]
  reg [6:0] cntValidOut; // @[SDFChainRadix22.scala 99:28]
  reg [31:0] _RAND_4;
  reg  lastWait; // @[SDFChainRadix22.scala 100:25]
  reg [31:0] _RAND_5;
  reg  lastIndeed; // @[SDFChainRadix22.scala 101:27]
  reg [31:0] _RAND_6;
  reg  initialInDone; // @[SDFChainRadix22.scala 102:30]
  reg [31:0] _RAND_7;
  reg  initialInDonePrev; // @[SDFChainRadix22.scala 103:34]
  reg [31:0] _RAND_8;
  wire [7:0] numPoints = _T_40[7:0]; // @[SDFChainRadix22.scala 46:23 SDFChainRadix22.scala 69:15]
  wire [7:0] _T_48 = numPoints - 8'h1; // @[SDFChainRadix22.scala 104:44]
  wire [7:0] _GEN_939 = {{1'd0}, cntValidOut}; // @[SDFChainRadix22.scala 104:29]
  wire  _T_49 = _GEN_939 == _T_48; // @[SDFChainRadix22.scala 104:29]
  wire  _T_50 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  wire  pktEnd = _T_49 & _T_50; // @[SDFChainRadix22.scala 104:52]
  wire  _T_51 = state_next == 2'h0; // @[SDFChainRadix22.scala 106:20]
  wire  _T_54 = cnt == _T_48; // @[SDFChainRadix22.scala 109:18]
  wire  _T_56 = _T_54 & _T_41; // @[SDFChainRadix22.scala 109:40]
  wire  _GEN_15 = _T_56 | initialInDone; // @[SDFChainRadix22.scala 109:57]
  wire  _T_58 = initialInDone & initialInDonePrev; // @[SDFChainRadix22.scala 117:41]
  wire  _T_59 = fireLast & _T_58; // @[SDFChainRadix22.scala 117:23]
  wire  _GEN_17 = _T_59 | lastWait; // @[SDFChainRadix22.scala 117:64]
  wire  _T_61 = _T_51 & pktEnd; // @[SDFChainRadix22.scala 121:30]
  wire [6:0] _T_64 = cntValidOut + 7'h1; // @[SDFChainRadix22.scala 125:32]
  wire  _T_66 = lastWait & pktEnd; // @[SDFChainRadix22.scala 131:23]
  wire  _GEN_21 = _T_66 | lastIndeed; // @[SDFChainRadix22.scala 131:34]
  wire  _T_67 = lastIndeed & pktEnd; // @[SDFChainRadix22.scala 135:132]
  wire  _T_68 = state == 2'h2; // @[SDFChainRadix22.scala 135:159]
  wire  _T_69 = pktEnd & _T_68; // @[SDFChainRadix22.scala 135:150]
  wire [6:0] _T_71 = 7'h7 - regNumStages; // @[SDFChainRadix22.scala 138:62]
  wire [6:0] _GEN_24 = 3'h1 == _T_71[2:0] ? 7'h40 : 7'h0; // @[SDFChainRadix22.scala 138:25]
  wire [6:0] _GEN_25 = 3'h2 == _T_71[2:0] ? 7'h60 : _GEN_24; // @[SDFChainRadix22.scala 138:25]
  wire [6:0] _GEN_26 = 3'h3 == _T_71[2:0] ? 7'h70 : _GEN_25; // @[SDFChainRadix22.scala 138:25]
  wire [6:0] _GEN_27 = 3'h4 == _T_71[2:0] ? 7'h78 : _GEN_26; // @[SDFChainRadix22.scala 138:25]
  wire [6:0] _GEN_28 = 3'h5 == _T_71[2:0] ? 7'h7c : _GEN_27; // @[SDFChainRadix22.scala 138:25]
  wire [6:0] _GEN_29 = 3'h6 == _T_71[2:0] ? 7'h7e : _GEN_28; // @[SDFChainRadix22.scala 138:25]
  wire [6:0] cumulativeDelayWire = 3'h7 == _T_71[2:0] ? 7'h7f : _GEN_29; // @[SDFChainRadix22.scala 138:25]
  wire  activeStages_0 = _T_71 <= 7'h0; // @[SDFChainRadix22.scala 146:48]
  wire  activeStages_1 = _T_71 <= 7'h1; // @[SDFChainRadix22.scala 146:48]
  wire  activeStages_2 = _T_71 <= 7'h2; // @[SDFChainRadix22.scala 146:48]
  wire  activeStages_3 = _T_71 <= 7'h3; // @[SDFChainRadix22.scala 146:48]
  wire  activeStages_4 = _T_71 <= 7'h4; // @[SDFChainRadix22.scala 146:48]
  wire  activeStages_5 = _T_71 <= 7'h5; // @[SDFChainRadix22.scala 146:48]
  wire  activeStages_6 = _T_71 <= 7'h6; // @[SDFChainRadix22.scala 146:48]
  wire  _T_103 = _T_68 & io_out_ready; // @[SDFChainRadix22.scala 164:54]
  wire  enableInit = _T_41 | _T_103; // @[SDFChainRadix22.scala 164:33]
  wire [7:0] _T_106 = cnt + 8'h1; // @[SDFChainRadix22.scala 170:16]
  reg  _T_108; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_9;
  reg  _T_109; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_10;
  reg  _T_110; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_11;
  reg  enableVector_1; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_12;
  reg [7:0] _T_113; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_13;
  reg [7:0] _T_114; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_14;
  reg [7:0] _T_115; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_15;
  reg [7:0] _T_116; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_16;
  reg  _T_118; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_17;
  reg  _T_119; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_18;
  reg  _T_120; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_19;
  reg  enableVector_2; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_20;
  reg [7:0] _T_123; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_21;
  reg [7:0] _T_124; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_22;
  reg [7:0] _T_125; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_23;
  reg [7:0] _T_126; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_24;
  reg  _T_128; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_25;
  reg  _T_129; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_26;
  reg  _T_130; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_27;
  reg  enableVector_3; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_28;
  reg [7:0] _T_133; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_29;
  reg [7:0] _T_134; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_30;
  reg [7:0] _T_135; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_31;
  reg [7:0] _T_136; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_32;
  reg  _T_138; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_33;
  reg  _T_139; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_34;
  reg  _T_140; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_35;
  reg  enableVector_4; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_36;
  reg [7:0] _T_143; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_37;
  reg [7:0] _T_144; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_38;
  reg [7:0] _T_145; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_39;
  reg [7:0] _T_146; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_40;
  reg  _T_148; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_41;
  reg  _T_149; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_42;
  reg  _T_150; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_43;
  reg  enableVector_5; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_44;
  reg [7:0] _T_153; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_45;
  reg [7:0] _T_154; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_46;
  reg [7:0] _T_155; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_47;
  reg [7:0] _T_156; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_48;
  reg  _T_158; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_49;
  reg  _T_159; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_50;
  reg  _T_160; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_51;
  reg  enableVector_6; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_52;
  reg [7:0] _T_163; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_53;
  reg [7:0] _T_164; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_54;
  reg [7:0] _T_165; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_55;
  reg [7:0] _T_166; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_56;
  wire [7:0] _T_184 = numPoints - 8'h2; // @[SDFChainRadix22.scala 186:37]
  wire [6:0] cntr_wires_0 = cnt[6:0]; // @[SDFChainRadix22.scala 48:24 SDFChainRadix22.scala 176:29]
  wire [6:0] cntr_wires_1 = _T_116[6:0]; // @[SDFChainRadix22.scala 48:24 SDFChainRadix22.scala 176:29]
  wire [6:0] _GEN_146 = 3'h1 == _T_39[2:0] ? cntr_wires_1 : cntr_wires_0; // @[SDFChainRadix22.scala 186:22]
  wire [6:0] cntr_wires_2 = _T_126[6:0]; // @[SDFChainRadix22.scala 48:24 SDFChainRadix22.scala 176:29]
  wire [6:0] _GEN_147 = 3'h2 == _T_39[2:0] ? cntr_wires_2 : _GEN_146; // @[SDFChainRadix22.scala 186:22]
  wire [6:0] cntr_wires_3 = _T_136[6:0]; // @[SDFChainRadix22.scala 48:24 SDFChainRadix22.scala 176:29]
  wire [6:0] _GEN_148 = 3'h3 == _T_39[2:0] ? cntr_wires_3 : _GEN_147; // @[SDFChainRadix22.scala 186:22]
  wire [6:0] cntr_wires_4 = _T_146[6:0]; // @[SDFChainRadix22.scala 48:24 SDFChainRadix22.scala 176:29]
  wire [6:0] _GEN_149 = 3'h4 == _T_39[2:0] ? cntr_wires_4 : _GEN_148; // @[SDFChainRadix22.scala 186:22]
  wire [6:0] cntr_wires_5 = _T_156[6:0]; // @[SDFChainRadix22.scala 48:24 SDFChainRadix22.scala 176:29]
  wire [6:0] _GEN_150 = 3'h5 == _T_39[2:0] ? cntr_wires_5 : _GEN_149; // @[SDFChainRadix22.scala 186:22]
  wire [6:0] cntr_wires_6 = _T_166[6:0]; // @[SDFChainRadix22.scala 48:24 SDFChainRadix22.scala 176:29]
  wire [6:0] _GEN_151 = 3'h6 == _T_39[2:0] ? cntr_wires_6 : _GEN_150; // @[SDFChainRadix22.scala 186:22]
  wire [7:0] _GEN_940 = {{1'd0}, _GEN_151}; // @[SDFChainRadix22.scala 186:22]
  wire  _T_185 = _GEN_940 == _T_184; // @[SDFChainRadix22.scala 186:22]
  wire  _GEN_153 = 3'h1 == _T_39[2:0] ? enableVector_1 : enableInit; // @[SDFChainRadix22.scala 186:44]
  wire  _GEN_154 = 3'h2 == _T_39[2:0] ? enableVector_2 : _GEN_153; // @[SDFChainRadix22.scala 186:44]
  wire  _GEN_155 = 3'h3 == _T_39[2:0] ? enableVector_3 : _GEN_154; // @[SDFChainRadix22.scala 186:44]
  wire  _GEN_156 = 3'h4 == _T_39[2:0] ? enableVector_4 : _GEN_155; // @[SDFChainRadix22.scala 186:44]
  wire  _GEN_157 = 3'h5 == _T_39[2:0] ? enableVector_5 : _GEN_156; // @[SDFChainRadix22.scala 186:44]
  wire  _GEN_158 = 3'h6 == _T_39[2:0] ? enableVector_6 : _GEN_157; // @[SDFChainRadix22.scala 186:44]
  wire  _T_186 = _T_185 & _GEN_158; // @[SDFChainRadix22.scala 186:44]
  wire  _GEN_159 = _T_51 ? 1'h0 : initialOutDone; // @[SDFChainRadix22.scala 189:36]
  wire  _GEN_160 = _T_186 | _GEN_159; // @[SDFChainRadix22.scala 186:60]
  wire  _T_188 = numPoints == 8'h2; // @[SDFChainRadix22.scala 193:43]
  reg  _T_189; // @[SDFChainRadix22.scala 193:59]
  reg [31:0] _RAND_57;
  wire  _T_191 = _T_189 & _T_41; // @[SDFChainRadix22.scala 193:72]
  wire  _T_192 = _GEN_158 & initialOutDone; // @[SDFChainRadix22.scala 193:101]
  wire [15:0] input_data_real = activeStages_0 ? $signed(io_in_bits_real) : $signed(16'sh0); // @[SDFChainRadix22.scala 211:23]
  wire [15:0] input_data_imag = activeStages_0 ? $signed(io_in_bits_imag) : $signed(16'sh0); // @[SDFChainRadix22.scala 211:23]
  wire  _T_202 = 7'h0 < _T_71; // @[SDFChainRadix22.scala 214:67]
  wire [6:0] _T_206 = 7'h0 - _T_71; // @[SDFChainRadix22.scala 215:63]
  wire  _GEN_164 = 3'h1 == _T_206[2:0] ? enableVector_1 : enableInit; // @[SDFChainRadix22.scala 216:20]
  wire  _GEN_165 = 3'h2 == _T_206[2:0] ? enableVector_2 : _GEN_164; // @[SDFChainRadix22.scala 216:20]
  wire  _GEN_166 = 3'h3 == _T_206[2:0] ? enableVector_3 : _GEN_165; // @[SDFChainRadix22.scala 216:20]
  wire  _GEN_167 = 3'h4 == _T_206[2:0] ? enableVector_4 : _GEN_166; // @[SDFChainRadix22.scala 216:20]
  wire  _GEN_168 = 3'h5 == _T_206[2:0] ? enableVector_5 : _GEN_167; // @[SDFChainRadix22.scala 216:20]
  wire  _GEN_169 = 3'h6 == _T_206[2:0] ? enableVector_6 : _GEN_168; // @[SDFChainRadix22.scala 216:20]
  wire [6:0] _T_211 = 7'h0 - cumulativeDelayWire; // @[SDFChainRadix22.scala 217:68]
  wire [6:0] _GEN_171 = 3'h1 == _T_206[2:0] ? cntr_wires_1 : cntr_wires_0; // @[SDFChainRadix22.scala 217:38]
  wire [6:0] _GEN_172 = 3'h2 == _T_206[2:0] ? cntr_wires_2 : _GEN_171; // @[SDFChainRadix22.scala 217:38]
  wire [6:0] _GEN_173 = 3'h3 == _T_206[2:0] ? cntr_wires_3 : _GEN_172; // @[SDFChainRadix22.scala 217:38]
  wire [6:0] _GEN_174 = 3'h4 == _T_206[2:0] ? cntr_wires_4 : _GEN_173; // @[SDFChainRadix22.scala 217:38]
  wire [6:0] _GEN_175 = 3'h5 == _T_206[2:0] ? cntr_wires_5 : _GEN_174; // @[SDFChainRadix22.scala 217:38]
  wire [6:0] _GEN_176 = 3'h6 == _T_206[2:0] ? cntr_wires_6 : _GEN_175; // @[SDFChainRadix22.scala 217:38]
  wire  _T_217 = 7'h1 < _T_71; // @[SDFChainRadix22.scala 214:67]
  wire [6:0] _T_221 = 7'h1 - _T_71; // @[SDFChainRadix22.scala 215:63]
  wire  _GEN_178 = 3'h1 == _T_221[2:0] ? enableVector_1 : enableInit; // @[SDFChainRadix22.scala 216:20]
  wire  _GEN_179 = 3'h2 == _T_221[2:0] ? enableVector_2 : _GEN_178; // @[SDFChainRadix22.scala 216:20]
  wire  _GEN_180 = 3'h3 == _T_221[2:0] ? enableVector_3 : _GEN_179; // @[SDFChainRadix22.scala 216:20]
  wire  _GEN_181 = 3'h4 == _T_221[2:0] ? enableVector_4 : _GEN_180; // @[SDFChainRadix22.scala 216:20]
  wire  _GEN_182 = 3'h5 == _T_221[2:0] ? enableVector_5 : _GEN_181; // @[SDFChainRadix22.scala 216:20]
  wire  _GEN_183 = 3'h6 == _T_221[2:0] ? enableVector_6 : _GEN_182; // @[SDFChainRadix22.scala 216:20]
  wire [6:0] _T_226 = 7'h40 - cumulativeDelayWire; // @[SDFChainRadix22.scala 217:68]
  wire [6:0] _GEN_185 = 3'h1 == _T_221[2:0] ? cntr_wires_1 : cntr_wires_0; // @[SDFChainRadix22.scala 217:38]
  wire [6:0] _GEN_186 = 3'h2 == _T_221[2:0] ? cntr_wires_2 : _GEN_185; // @[SDFChainRadix22.scala 217:38]
  wire [6:0] _GEN_187 = 3'h3 == _T_221[2:0] ? cntr_wires_3 : _GEN_186; // @[SDFChainRadix22.scala 217:38]
  wire [6:0] _GEN_188 = 3'h4 == _T_221[2:0] ? cntr_wires_4 : _GEN_187; // @[SDFChainRadix22.scala 217:38]
  wire [6:0] _GEN_189 = 3'h5 == _T_221[2:0] ? cntr_wires_5 : _GEN_188; // @[SDFChainRadix22.scala 217:38]
  wire [6:0] _GEN_190 = 3'h6 == _T_221[2:0] ? cntr_wires_6 : _GEN_189; // @[SDFChainRadix22.scala 217:38]
  wire [6:0] _T_228 = _GEN_190 - _T_226; // @[SDFChainRadix22.scala 217:38]
  wire  _T_232 = 7'h2 < _T_71; // @[SDFChainRadix22.scala 214:67]
  wire [6:0] _T_236 = 7'h2 - _T_71; // @[SDFChainRadix22.scala 215:63]
  wire  _GEN_192 = 3'h1 == _T_236[2:0] ? enableVector_1 : enableInit; // @[SDFChainRadix22.scala 216:20]
  wire  _GEN_193 = 3'h2 == _T_236[2:0] ? enableVector_2 : _GEN_192; // @[SDFChainRadix22.scala 216:20]
  wire  _GEN_194 = 3'h3 == _T_236[2:0] ? enableVector_3 : _GEN_193; // @[SDFChainRadix22.scala 216:20]
  wire  _GEN_195 = 3'h4 == _T_236[2:0] ? enableVector_4 : _GEN_194; // @[SDFChainRadix22.scala 216:20]
  wire  _GEN_196 = 3'h5 == _T_236[2:0] ? enableVector_5 : _GEN_195; // @[SDFChainRadix22.scala 216:20]
  wire  _GEN_197 = 3'h6 == _T_236[2:0] ? enableVector_6 : _GEN_196; // @[SDFChainRadix22.scala 216:20]
  wire [6:0] _T_241 = 7'h60 - cumulativeDelayWire; // @[SDFChainRadix22.scala 217:68]
  wire [6:0] _GEN_199 = 3'h1 == _T_236[2:0] ? cntr_wires_1 : cntr_wires_0; // @[SDFChainRadix22.scala 217:38]
  wire [6:0] _GEN_200 = 3'h2 == _T_236[2:0] ? cntr_wires_2 : _GEN_199; // @[SDFChainRadix22.scala 217:38]
  wire [6:0] _GEN_201 = 3'h3 == _T_236[2:0] ? cntr_wires_3 : _GEN_200; // @[SDFChainRadix22.scala 217:38]
  wire [6:0] _GEN_202 = 3'h4 == _T_236[2:0] ? cntr_wires_4 : _GEN_201; // @[SDFChainRadix22.scala 217:38]
  wire [6:0] _GEN_203 = 3'h5 == _T_236[2:0] ? cntr_wires_5 : _GEN_202; // @[SDFChainRadix22.scala 217:38]
  wire [6:0] _GEN_204 = 3'h6 == _T_236[2:0] ? cntr_wires_6 : _GEN_203; // @[SDFChainRadix22.scala 217:38]
  wire [6:0] _T_243 = _GEN_204 - _T_241; // @[SDFChainRadix22.scala 217:38]
  wire  _T_247 = 7'h3 < _T_71; // @[SDFChainRadix22.scala 214:67]
  wire [6:0] _T_251 = 7'h3 - _T_71; // @[SDFChainRadix22.scala 215:63]
  wire  _GEN_206 = 3'h1 == _T_251[2:0] ? enableVector_1 : enableInit; // @[SDFChainRadix22.scala 216:20]
  wire  _GEN_207 = 3'h2 == _T_251[2:0] ? enableVector_2 : _GEN_206; // @[SDFChainRadix22.scala 216:20]
  wire  _GEN_208 = 3'h3 == _T_251[2:0] ? enableVector_3 : _GEN_207; // @[SDFChainRadix22.scala 216:20]
  wire  _GEN_209 = 3'h4 == _T_251[2:0] ? enableVector_4 : _GEN_208; // @[SDFChainRadix22.scala 216:20]
  wire  _GEN_210 = 3'h5 == _T_251[2:0] ? enableVector_5 : _GEN_209; // @[SDFChainRadix22.scala 216:20]
  wire  _GEN_211 = 3'h6 == _T_251[2:0] ? enableVector_6 : _GEN_210; // @[SDFChainRadix22.scala 216:20]
  wire [6:0] _T_256 = 7'h70 - cumulativeDelayWire; // @[SDFChainRadix22.scala 217:68]
  wire [6:0] _GEN_213 = 3'h1 == _T_251[2:0] ? cntr_wires_1 : cntr_wires_0; // @[SDFChainRadix22.scala 217:38]
  wire [6:0] _GEN_214 = 3'h2 == _T_251[2:0] ? cntr_wires_2 : _GEN_213; // @[SDFChainRadix22.scala 217:38]
  wire [6:0] _GEN_215 = 3'h3 == _T_251[2:0] ? cntr_wires_3 : _GEN_214; // @[SDFChainRadix22.scala 217:38]
  wire [6:0] _GEN_216 = 3'h4 == _T_251[2:0] ? cntr_wires_4 : _GEN_215; // @[SDFChainRadix22.scala 217:38]
  wire [6:0] _GEN_217 = 3'h5 == _T_251[2:0] ? cntr_wires_5 : _GEN_216; // @[SDFChainRadix22.scala 217:38]
  wire [6:0] _GEN_218 = 3'h6 == _T_251[2:0] ? cntr_wires_6 : _GEN_217; // @[SDFChainRadix22.scala 217:38]
  wire [6:0] _T_258 = _GEN_218 - _T_256; // @[SDFChainRadix22.scala 217:38]
  wire  _T_262 = 7'h4 < _T_71; // @[SDFChainRadix22.scala 214:67]
  wire [6:0] _T_266 = 7'h4 - _T_71; // @[SDFChainRadix22.scala 215:63]
  wire  _GEN_220 = 3'h1 == _T_266[2:0] ? enableVector_1 : enableInit; // @[SDFChainRadix22.scala 216:20]
  wire  _GEN_221 = 3'h2 == _T_266[2:0] ? enableVector_2 : _GEN_220; // @[SDFChainRadix22.scala 216:20]
  wire  _GEN_222 = 3'h3 == _T_266[2:0] ? enableVector_3 : _GEN_221; // @[SDFChainRadix22.scala 216:20]
  wire  _GEN_223 = 3'h4 == _T_266[2:0] ? enableVector_4 : _GEN_222; // @[SDFChainRadix22.scala 216:20]
  wire  _GEN_224 = 3'h5 == _T_266[2:0] ? enableVector_5 : _GEN_223; // @[SDFChainRadix22.scala 216:20]
  wire  _GEN_225 = 3'h6 == _T_266[2:0] ? enableVector_6 : _GEN_224; // @[SDFChainRadix22.scala 216:20]
  wire [6:0] _T_271 = 7'h78 - cumulativeDelayWire; // @[SDFChainRadix22.scala 217:68]
  wire [6:0] _GEN_227 = 3'h1 == _T_266[2:0] ? cntr_wires_1 : cntr_wires_0; // @[SDFChainRadix22.scala 217:38]
  wire [6:0] _GEN_228 = 3'h2 == _T_266[2:0] ? cntr_wires_2 : _GEN_227; // @[SDFChainRadix22.scala 217:38]
  wire [6:0] _GEN_229 = 3'h3 == _T_266[2:0] ? cntr_wires_3 : _GEN_228; // @[SDFChainRadix22.scala 217:38]
  wire [6:0] _GEN_230 = 3'h4 == _T_266[2:0] ? cntr_wires_4 : _GEN_229; // @[SDFChainRadix22.scala 217:38]
  wire [6:0] _GEN_231 = 3'h5 == _T_266[2:0] ? cntr_wires_5 : _GEN_230; // @[SDFChainRadix22.scala 217:38]
  wire [6:0] _GEN_232 = 3'h6 == _T_266[2:0] ? cntr_wires_6 : _GEN_231; // @[SDFChainRadix22.scala 217:38]
  wire [6:0] _T_273 = _GEN_232 - _T_271; // @[SDFChainRadix22.scala 217:38]
  wire  _T_277 = 7'h5 < _T_71; // @[SDFChainRadix22.scala 214:67]
  wire [6:0] _T_281 = 7'h5 - _T_71; // @[SDFChainRadix22.scala 215:63]
  wire  _GEN_234 = 3'h1 == _T_281[2:0] ? enableVector_1 : enableInit; // @[SDFChainRadix22.scala 216:20]
  wire  _GEN_235 = 3'h2 == _T_281[2:0] ? enableVector_2 : _GEN_234; // @[SDFChainRadix22.scala 216:20]
  wire  _GEN_236 = 3'h3 == _T_281[2:0] ? enableVector_3 : _GEN_235; // @[SDFChainRadix22.scala 216:20]
  wire  _GEN_237 = 3'h4 == _T_281[2:0] ? enableVector_4 : _GEN_236; // @[SDFChainRadix22.scala 216:20]
  wire  _GEN_238 = 3'h5 == _T_281[2:0] ? enableVector_5 : _GEN_237; // @[SDFChainRadix22.scala 216:20]
  wire  _GEN_239 = 3'h6 == _T_281[2:0] ? enableVector_6 : _GEN_238; // @[SDFChainRadix22.scala 216:20]
  wire [6:0] _T_286 = 7'h7c - cumulativeDelayWire; // @[SDFChainRadix22.scala 217:68]
  wire [6:0] _GEN_241 = 3'h1 == _T_281[2:0] ? cntr_wires_1 : cntr_wires_0; // @[SDFChainRadix22.scala 217:38]
  wire [6:0] _GEN_242 = 3'h2 == _T_281[2:0] ? cntr_wires_2 : _GEN_241; // @[SDFChainRadix22.scala 217:38]
  wire [6:0] _GEN_243 = 3'h3 == _T_281[2:0] ? cntr_wires_3 : _GEN_242; // @[SDFChainRadix22.scala 217:38]
  wire [6:0] _GEN_244 = 3'h4 == _T_281[2:0] ? cntr_wires_4 : _GEN_243; // @[SDFChainRadix22.scala 217:38]
  wire [6:0] _GEN_245 = 3'h5 == _T_281[2:0] ? cntr_wires_5 : _GEN_244; // @[SDFChainRadix22.scala 217:38]
  wire [6:0] _GEN_246 = 3'h6 == _T_281[2:0] ? cntr_wires_6 : _GEN_245; // @[SDFChainRadix22.scala 217:38]
  wire [6:0] _T_288 = _GEN_246 - _T_286; // @[SDFChainRadix22.scala 217:38]
  wire  _T_292 = 7'h6 < _T_71; // @[SDFChainRadix22.scala 214:67]
  wire [6:0] _T_296 = 7'h6 - _T_71; // @[SDFChainRadix22.scala 215:63]
  wire  _GEN_248 = 3'h1 == _T_296[2:0] ? enableVector_1 : enableInit; // @[SDFChainRadix22.scala 216:20]
  wire  _GEN_249 = 3'h2 == _T_296[2:0] ? enableVector_2 : _GEN_248; // @[SDFChainRadix22.scala 216:20]
  wire  _GEN_250 = 3'h3 == _T_296[2:0] ? enableVector_3 : _GEN_249; // @[SDFChainRadix22.scala 216:20]
  wire  _GEN_251 = 3'h4 == _T_296[2:0] ? enableVector_4 : _GEN_250; // @[SDFChainRadix22.scala 216:20]
  wire  _GEN_252 = 3'h5 == _T_296[2:0] ? enableVector_5 : _GEN_251; // @[SDFChainRadix22.scala 216:20]
  wire  _GEN_253 = 3'h6 == _T_296[2:0] ? enableVector_6 : _GEN_252; // @[SDFChainRadix22.scala 216:20]
  wire [6:0] _T_301 = 7'h7e - cumulativeDelayWire; // @[SDFChainRadix22.scala 217:68]
  wire [6:0] _GEN_255 = 3'h1 == _T_296[2:0] ? cntr_wires_1 : cntr_wires_0; // @[SDFChainRadix22.scala 217:38]
  wire [6:0] _GEN_256 = 3'h2 == _T_296[2:0] ? cntr_wires_2 : _GEN_255; // @[SDFChainRadix22.scala 217:38]
  wire [6:0] _GEN_257 = 3'h3 == _T_296[2:0] ? cntr_wires_3 : _GEN_256; // @[SDFChainRadix22.scala 217:38]
  wire [6:0] _GEN_258 = 3'h4 == _T_296[2:0] ? cntr_wires_4 : _GEN_257; // @[SDFChainRadix22.scala 217:38]
  wire [6:0] _GEN_259 = 3'h5 == _T_296[2:0] ? cntr_wires_5 : _GEN_258; // @[SDFChainRadix22.scala 217:38]
  wire [6:0] _GEN_260 = 3'h6 == _T_296[2:0] ? cntr_wires_6 : _GEN_259; // @[SDFChainRadix22.scala 217:38]
  wire [6:0] _T_303 = _GEN_260 - _T_301; // @[SDFChainRadix22.scala 217:38]
  wire  _T_310 = 7'h0 == _T_71; // @[SDFChainRadix22.scala 234:23]
  wire [15:0] _GEN_261 = _T_310 ? $signed(io_in_bits_imag) : $signed(input_data_imag); // @[SDFChainRadix22.scala 234:55]
  wire [15:0] _GEN_262 = _T_310 ? $signed(io_in_bits_real) : $signed(input_data_real); // @[SDFChainRadix22.scala 234:55]
  wire  _T_311 = sdf_stages_0_io_cntr < 7'h40; // @[SDFChainRadix22.scala 320:98]
  wire  _T_313 = sdf_stages_0_io_cntr < 7'h20; // @[SDFChainRadix22.scala 320:135]
  wire  _T_314 = _T_313 ? 1'h0 : 1'h1; // @[SDFChainRadix22.scala 320:122]
  reg  _T_316; // @[Reg.scala 15:16]
  reg [31:0] _RAND_58;
  wire [15:0] _T_322 = 16'sh0 - $signed(sdf_stages_0_io_out_real); // @[FixedPointTypeClass.scala 39:43]
  wire [15:0] _T_319_real = sdf_stages_0_io_out_imag; // @[SDFChainRadix22.scala 322:32 SDFChainRadix22.scala 325:29]
  reg [15:0] _T_328_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_59;
  reg [15:0] _T_328_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_60;
  reg [15:0] _T_331_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_61;
  reg [15:0] _T_331_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_62;
  reg [15:0] outputWires_0_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_63;
  reg [15:0] outputWires_0_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_64;
  wire  _T_340 = 7'h1 == _T_71; // @[SDFChainRadix22.scala 234:23]
  wire [15:0] _GEN_272 = _T_340 ? $signed(io_in_bits_imag) : $signed(outputWires_0_imag); // @[SDFChainRadix22.scala 234:55]
  wire [15:0] _GEN_273 = _T_340 ? $signed(io_in_bits_real) : $signed(outputWires_0_real); // @[SDFChainRadix22.scala 234:55]
  wire [6:0] _T_673 = _GEN_190 + 7'h1; // @[SDFChainRadix22.scala 276:83]
  wire [6:0] _T_677 = _T_673 - _T_241; // @[SDFChainRadix22.scala 276:89]
  reg [6:0] _T_679; // @[Reg.scala 15:16]
  reg [31:0] _RAND_65;
  reg [15:0] twiddles_1_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_66;
  reg [15:0] twiddles_1_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_67;
  wire [5:0] _GEN_331 = 7'h21 == _T_679 ? 6'h2 : 6'h0; // @[Reg.scala 16:23]
  wire [5:0] _GEN_332 = 7'h22 == _T_679 ? 6'h4 : _GEN_331; // @[Reg.scala 16:23]
  wire [5:0] _GEN_333 = 7'h23 == _T_679 ? 6'h6 : _GEN_332; // @[Reg.scala 16:23]
  wire [5:0] _GEN_334 = 7'h24 == _T_679 ? 6'h8 : _GEN_333; // @[Reg.scala 16:23]
  wire [5:0] _GEN_335 = 7'h25 == _T_679 ? 6'ha : _GEN_334; // @[Reg.scala 16:23]
  wire [5:0] _GEN_336 = 7'h26 == _T_679 ? 6'hc : _GEN_335; // @[Reg.scala 16:23]
  wire [5:0] _GEN_337 = 7'h27 == _T_679 ? 6'he : _GEN_336; // @[Reg.scala 16:23]
  wire [5:0] _GEN_338 = 7'h28 == _T_679 ? 6'h10 : _GEN_337; // @[Reg.scala 16:23]
  wire [5:0] _GEN_339 = 7'h29 == _T_679 ? 6'h12 : _GEN_338; // @[Reg.scala 16:23]
  wire [5:0] _GEN_340 = 7'h2a == _T_679 ? 6'h14 : _GEN_339; // @[Reg.scala 16:23]
  wire [5:0] _GEN_341 = 7'h2b == _T_679 ? 6'h16 : _GEN_340; // @[Reg.scala 16:23]
  wire [5:0] _GEN_342 = 7'h2c == _T_679 ? 6'h18 : _GEN_341; // @[Reg.scala 16:23]
  wire [5:0] _GEN_343 = 7'h2d == _T_679 ? 6'h1a : _GEN_342; // @[Reg.scala 16:23]
  wire [5:0] _GEN_344 = 7'h2e == _T_679 ? 6'h1c : _GEN_343; // @[Reg.scala 16:23]
  wire [5:0] _GEN_345 = 7'h2f == _T_679 ? 6'h1e : _GEN_344; // @[Reg.scala 16:23]
  wire [5:0] _GEN_346 = 7'h30 == _T_679 ? 6'h20 : _GEN_345; // @[Reg.scala 16:23]
  wire [5:0] _GEN_347 = 7'h31 == _T_679 ? 6'h22 : _GEN_346; // @[Reg.scala 16:23]
  wire [5:0] _GEN_348 = 7'h32 == _T_679 ? 6'h23 : _GEN_347; // @[Reg.scala 16:23]
  wire [5:0] _GEN_349 = 7'h33 == _T_679 ? 6'h24 : _GEN_348; // @[Reg.scala 16:23]
  wire [5:0] _GEN_350 = 7'h34 == _T_679 ? 6'h26 : _GEN_349; // @[Reg.scala 16:23]
  wire [5:0] _GEN_351 = 7'h35 == _T_679 ? 6'h27 : _GEN_350; // @[Reg.scala 16:23]
  wire [5:0] _GEN_352 = 7'h36 == _T_679 ? 6'h28 : _GEN_351; // @[Reg.scala 16:23]
  wire [5:0] _GEN_353 = 7'h37 == _T_679 ? 6'h2a : _GEN_352; // @[Reg.scala 16:23]
  wire [5:0] _GEN_354 = 7'h38 == _T_679 ? 6'h2b : _GEN_353; // @[Reg.scala 16:23]
  wire [5:0] _GEN_355 = 7'h39 == _T_679 ? 6'h2c : _GEN_354; // @[Reg.scala 16:23]
  wire [5:0] _GEN_356 = 7'h3a == _T_679 ? 6'h2e : _GEN_355; // @[Reg.scala 16:23]
  wire [5:0] _GEN_357 = 7'h3b == _T_679 ? 6'h2f : _GEN_356; // @[Reg.scala 16:23]
  wire [5:0] _GEN_358 = 7'h3c == _T_679 ? 6'h30 : _GEN_357; // @[Reg.scala 16:23]
  wire [5:0] _GEN_359 = 7'h3d == _T_679 ? 6'h32 : _GEN_358; // @[Reg.scala 16:23]
  wire [5:0] _GEN_360 = 7'h3e == _T_679 ? 6'h33 : _GEN_359; // @[Reg.scala 16:23]
  wire [5:0] _GEN_361 = 7'h3f == _T_679 ? 6'h34 : _GEN_360; // @[Reg.scala 16:23]
  wire [5:0] _GEN_362 = 7'h40 == _T_679 ? 6'h0 : _GEN_361; // @[Reg.scala 16:23]
  wire [5:0] _GEN_363 = 7'h41 == _T_679 ? 6'h1 : _GEN_362; // @[Reg.scala 16:23]
  wire [5:0] _GEN_364 = 7'h42 == _T_679 ? 6'h2 : _GEN_363; // @[Reg.scala 16:23]
  wire [5:0] _GEN_365 = 7'h43 == _T_679 ? 6'h3 : _GEN_364; // @[Reg.scala 16:23]
  wire [5:0] _GEN_366 = 7'h44 == _T_679 ? 6'h4 : _GEN_365; // @[Reg.scala 16:23]
  wire [5:0] _GEN_367 = 7'h45 == _T_679 ? 6'h5 : _GEN_366; // @[Reg.scala 16:23]
  wire [5:0] _GEN_368 = 7'h46 == _T_679 ? 6'h6 : _GEN_367; // @[Reg.scala 16:23]
  wire [5:0] _GEN_369 = 7'h47 == _T_679 ? 6'h7 : _GEN_368; // @[Reg.scala 16:23]
  wire [5:0] _GEN_370 = 7'h48 == _T_679 ? 6'h8 : _GEN_369; // @[Reg.scala 16:23]
  wire [5:0] _GEN_371 = 7'h49 == _T_679 ? 6'h9 : _GEN_370; // @[Reg.scala 16:23]
  wire [5:0] _GEN_372 = 7'h4a == _T_679 ? 6'ha : _GEN_371; // @[Reg.scala 16:23]
  wire [5:0] _GEN_373 = 7'h4b == _T_679 ? 6'hb : _GEN_372; // @[Reg.scala 16:23]
  wire [5:0] _GEN_374 = 7'h4c == _T_679 ? 6'hc : _GEN_373; // @[Reg.scala 16:23]
  wire [5:0] _GEN_375 = 7'h4d == _T_679 ? 6'hd : _GEN_374; // @[Reg.scala 16:23]
  wire [5:0] _GEN_376 = 7'h4e == _T_679 ? 6'he : _GEN_375; // @[Reg.scala 16:23]
  wire [5:0] _GEN_377 = 7'h4f == _T_679 ? 6'hf : _GEN_376; // @[Reg.scala 16:23]
  wire [5:0] _GEN_378 = 7'h50 == _T_679 ? 6'h10 : _GEN_377; // @[Reg.scala 16:23]
  wire [5:0] _GEN_379 = 7'h51 == _T_679 ? 6'h11 : _GEN_378; // @[Reg.scala 16:23]
  wire [5:0] _GEN_380 = 7'h52 == _T_679 ? 6'h12 : _GEN_379; // @[Reg.scala 16:23]
  wire [5:0] _GEN_381 = 7'h53 == _T_679 ? 6'h13 : _GEN_380; // @[Reg.scala 16:23]
  wire [5:0] _GEN_382 = 7'h54 == _T_679 ? 6'h14 : _GEN_381; // @[Reg.scala 16:23]
  wire [5:0] _GEN_383 = 7'h55 == _T_679 ? 6'h15 : _GEN_382; // @[Reg.scala 16:23]
  wire [5:0] _GEN_384 = 7'h56 == _T_679 ? 6'h16 : _GEN_383; // @[Reg.scala 16:23]
  wire [5:0] _GEN_385 = 7'h57 == _T_679 ? 6'h17 : _GEN_384; // @[Reg.scala 16:23]
  wire [5:0] _GEN_386 = 7'h58 == _T_679 ? 6'h18 : _GEN_385; // @[Reg.scala 16:23]
  wire [5:0] _GEN_387 = 7'h59 == _T_679 ? 6'h19 : _GEN_386; // @[Reg.scala 16:23]
  wire [5:0] _GEN_388 = 7'h5a == _T_679 ? 6'h1a : _GEN_387; // @[Reg.scala 16:23]
  wire [5:0] _GEN_389 = 7'h5b == _T_679 ? 6'h1b : _GEN_388; // @[Reg.scala 16:23]
  wire [5:0] _GEN_390 = 7'h5c == _T_679 ? 6'h1c : _GEN_389; // @[Reg.scala 16:23]
  wire [5:0] _GEN_391 = 7'h5d == _T_679 ? 6'h1d : _GEN_390; // @[Reg.scala 16:23]
  wire [5:0] _GEN_392 = 7'h5e == _T_679 ? 6'h1e : _GEN_391; // @[Reg.scala 16:23]
  wire [5:0] _GEN_393 = 7'h5f == _T_679 ? 6'h1f : _GEN_392; // @[Reg.scala 16:23]
  wire [5:0] _GEN_394 = 7'h60 == _T_679 ? 6'h0 : _GEN_393; // @[Reg.scala 16:23]
  wire [5:0] _GEN_395 = 7'h61 == _T_679 ? 6'h3 : _GEN_394; // @[Reg.scala 16:23]
  wire [5:0] _GEN_396 = 7'h62 == _T_679 ? 6'h6 : _GEN_395; // @[Reg.scala 16:23]
  wire [5:0] _GEN_397 = 7'h63 == _T_679 ? 6'h9 : _GEN_396; // @[Reg.scala 16:23]
  wire [5:0] _GEN_398 = 7'h64 == _T_679 ? 6'hc : _GEN_397; // @[Reg.scala 16:23]
  wire [5:0] _GEN_399 = 7'h65 == _T_679 ? 6'hf : _GEN_398; // @[Reg.scala 16:23]
  wire [5:0] _GEN_400 = 7'h66 == _T_679 ? 6'h12 : _GEN_399; // @[Reg.scala 16:23]
  wire [5:0] _GEN_401 = 7'h67 == _T_679 ? 6'h15 : _GEN_400; // @[Reg.scala 16:23]
  wire [5:0] _GEN_402 = 7'h68 == _T_679 ? 6'h18 : _GEN_401; // @[Reg.scala 16:23]
  wire [5:0] _GEN_403 = 7'h69 == _T_679 ? 6'h1b : _GEN_402; // @[Reg.scala 16:23]
  wire [5:0] _GEN_404 = 7'h6a == _T_679 ? 6'h1e : _GEN_403; // @[Reg.scala 16:23]
  wire [5:0] _GEN_405 = 7'h6b == _T_679 ? 6'h21 : _GEN_404; // @[Reg.scala 16:23]
  wire [5:0] _GEN_406 = 7'h6c == _T_679 ? 6'h23 : _GEN_405; // @[Reg.scala 16:23]
  wire [5:0] _GEN_407 = 7'h6d == _T_679 ? 6'h25 : _GEN_406; // @[Reg.scala 16:23]
  wire [5:0] _GEN_408 = 7'h6e == _T_679 ? 6'h27 : _GEN_407; // @[Reg.scala 16:23]
  wire [5:0] _GEN_409 = 7'h6f == _T_679 ? 6'h29 : _GEN_408; // @[Reg.scala 16:23]
  wire [5:0] _GEN_410 = 7'h70 == _T_679 ? 6'h2b : _GEN_409; // @[Reg.scala 16:23]
  wire [5:0] _GEN_411 = 7'h71 == _T_679 ? 6'h2d : _GEN_410; // @[Reg.scala 16:23]
  wire [5:0] _GEN_412 = 7'h72 == _T_679 ? 6'h2f : _GEN_411; // @[Reg.scala 16:23]
  wire [5:0] _GEN_413 = 7'h73 == _T_679 ? 6'h31 : _GEN_412; // @[Reg.scala 16:23]
  wire [5:0] _GEN_414 = 7'h74 == _T_679 ? 6'h33 : _GEN_413; // @[Reg.scala 16:23]
  wire [5:0] _GEN_415 = 7'h75 == _T_679 ? 6'h35 : _GEN_414; // @[Reg.scala 16:23]
  wire [5:0] _GEN_416 = 7'h76 == _T_679 ? 6'h36 : _GEN_415; // @[Reg.scala 16:23]
  wire [5:0] _GEN_417 = 7'h77 == _T_679 ? 6'h37 : _GEN_416; // @[Reg.scala 16:23]
  wire [5:0] _GEN_418 = 7'h78 == _T_679 ? 6'h38 : _GEN_417; // @[Reg.scala 16:23]
  wire [5:0] _GEN_419 = 7'h79 == _T_679 ? 6'h39 : _GEN_418; // @[Reg.scala 16:23]
  wire [5:0] _GEN_420 = 7'h7a == _T_679 ? 6'h3a : _GEN_419; // @[Reg.scala 16:23]
  wire [5:0] _GEN_421 = 7'h7b == _T_679 ? 6'h3b : _GEN_420; // @[Reg.scala 16:23]
  wire [5:0] _GEN_422 = 7'h7c == _T_679 ? 6'h3c : _GEN_421; // @[Reg.scala 16:23]
  wire [5:0] _GEN_423 = 7'h7d == _T_679 ? 6'h3d : _GEN_422; // @[Reg.scala 16:23]
  wire [5:0] _GEN_424 = 7'h7e == _T_679 ? 6'h3e : _GEN_423; // @[Reg.scala 16:23]
  wire [5:0] _GEN_425 = 7'h7f == _T_679 ? 6'h3f : _GEN_424; // @[Reg.scala 16:23]
  reg [15:0] _T_688; // @[Reg.scala 15:16]
  reg [31:0] _RAND_68;
  reg [15:0] _T_689; // @[Reg.scala 15:16]
  reg [31:0] _RAND_69;
  reg [15:0] _T_690; // @[Reg.scala 15:16]
  reg [31:0] _RAND_70;
  reg [16:0] _T_692; // @[Reg.scala 15:16]
  reg [31:0] _RAND_71;
  reg [16:0] _T_694; // @[Reg.scala 15:16]
  reg [31:0] _RAND_72;
  reg [16:0] _T_696; // @[Reg.scala 15:16]
  reg [31:0] _RAND_73;
  wire [16:0] _GEN_941 = {{1{_T_688[15]}},_T_688}; // @[FixedPointTypeClass.scala 211:35]
  reg [32:0] _T_698; // @[Reg.scala 15:16]
  reg [63:0] _RAND_74;
  wire [34:0] _GEN_942 = {$signed(_T_698), 2'h0}; // @[FixedPointTypeClass.scala 20:58]
  wire [34:0] _T_701 = $signed(_GEN_942) + 35'sh1; // @[FixedPointTypeClass.scala 20:58]
  wire [33:0] _T_702 = _T_701[34:1]; // @[FixedPointTypeClass.scala 176:41]
  wire [16:0] _GEN_943 = {{1{_T_690[15]}},_T_690}; // @[FixedPointTypeClass.scala 211:35]
  reg [32:0] _T_704; // @[Reg.scala 15:16]
  reg [63:0] _RAND_75;
  wire [34:0] _GEN_944 = {$signed(_T_704), 2'h0}; // @[FixedPointTypeClass.scala 20:58]
  wire [34:0] _T_707 = $signed(_GEN_944) + 35'sh1; // @[FixedPointTypeClass.scala 20:58]
  wire [33:0] _T_708 = _T_707[34:1]; // @[FixedPointTypeClass.scala 176:41]
  wire [16:0] _GEN_945 = {{1{_T_689[15]}},_T_689}; // @[FixedPointTypeClass.scala 211:35]
  reg [32:0] _T_710; // @[Reg.scala 15:16]
  reg [63:0] _RAND_76;
  wire [34:0] _GEN_946 = {$signed(_T_710), 2'h0}; // @[FixedPointTypeClass.scala 20:58]
  wire [34:0] _T_713 = $signed(_GEN_946) + 35'sh1; // @[FixedPointTypeClass.scala 20:58]
  wire [33:0] _T_714 = _T_713[34:1]; // @[FixedPointTypeClass.scala 176:41]
  reg [34:0] _T_716; // @[Reg.scala 15:16]
  reg [63:0] _RAND_77;
  reg [34:0] _T_718; // @[Reg.scala 15:16]
  reg [63:0] _RAND_78;
  wire [34:0] _T_724 = $signed(_T_716) + 35'sh4000; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] _T_725 = _T_724[34:15]; // @[FixedPointTypeClass.scala 176:41]
  wire [34:0] _T_728 = $signed(_T_718) + 35'sh4000; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] _T_729 = _T_728[34:15]; // @[FixedPointTypeClass.scala 176:41]
  wire  _T_738 = 7'h2 == _T_71; // @[SDFChainRadix22.scala 234:23]
  wire [15:0] outputWires_1_imag = _T_729[15:0]; // @[SDFChainRadix22.scala 286:27 SDFChainRadix22.scala 306:19]
  wire [15:0] _GEN_695 = _T_738 ? $signed(io_in_bits_imag) : $signed(outputWires_1_imag); // @[SDFChainRadix22.scala 234:55]
  wire [15:0] outputWires_1_real = _T_725[15:0]; // @[SDFChainRadix22.scala 286:27 SDFChainRadix22.scala 306:19]
  wire [15:0] _GEN_696 = _T_738 ? $signed(io_in_bits_real) : $signed(outputWires_1_real); // @[SDFChainRadix22.scala 234:55]
  wire  _T_739 = sdf_stages_2_io_cntr < 7'h10; // @[SDFChainRadix22.scala 320:98]
  wire  _T_741 = sdf_stages_2_io_cntr < 7'h8; // @[SDFChainRadix22.scala 320:135]
  wire  _T_742 = _T_741 ? 1'h0 : 1'h1; // @[SDFChainRadix22.scala 320:122]
  reg  _T_744; // @[Reg.scala 15:16]
  reg [31:0] _RAND_79;
  wire [15:0] _T_750 = 16'sh0 - $signed(sdf_stages_2_io_out_real); // @[FixedPointTypeClass.scala 39:43]
  wire [15:0] _T_747_real = sdf_stages_2_io_out_imag; // @[SDFChainRadix22.scala 322:32 SDFChainRadix22.scala 325:29]
  reg [15:0] _T_756_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_80;
  reg [15:0] _T_756_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_81;
  reg [15:0] _T_759_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_82;
  reg [15:0] _T_759_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_83;
  reg [15:0] outputWires_2_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_84;
  reg [15:0] outputWires_2_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_85;
  wire  _T_768 = 7'h3 == _T_71; // @[SDFChainRadix22.scala 234:23]
  wire [15:0] _GEN_706 = _T_768 ? $signed(io_in_bits_imag) : $signed(outputWires_2_imag); // @[SDFChainRadix22.scala 234:55]
  wire [15:0] _GEN_707 = _T_768 ? $signed(io_in_bits_real) : $signed(outputWires_2_real); // @[SDFChainRadix22.scala 234:55]
  wire [6:0] _T_861 = _GEN_218 + 7'h1; // @[SDFChainRadix22.scala 276:83]
  wire [6:0] _T_865 = _T_861 - _T_271; // @[SDFChainRadix22.scala 276:89]
  reg [6:0] _T_867; // @[Reg.scala 15:16]
  reg [31:0] _RAND_86;
  reg [15:0] twiddles_3_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_87;
  reg [15:0] twiddles_3_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_88;
  wire [3:0] _GEN_741 = 5'h9 == _T_867[4:0] ? 4'h2 : 4'h0; // @[Reg.scala 16:23]
  wire [3:0] _GEN_742 = 5'ha == _T_867[4:0] ? 4'h4 : _GEN_741; // @[Reg.scala 16:23]
  wire [3:0] _GEN_743 = 5'hb == _T_867[4:0] ? 4'h6 : _GEN_742; // @[Reg.scala 16:23]
  wire [3:0] _GEN_744 = 5'hc == _T_867[4:0] ? 4'h8 : _GEN_743; // @[Reg.scala 16:23]
  wire [3:0] _GEN_745 = 5'hd == _T_867[4:0] ? 4'ha : _GEN_744; // @[Reg.scala 16:23]
  wire [3:0] _GEN_746 = 5'he == _T_867[4:0] ? 4'hb : _GEN_745; // @[Reg.scala 16:23]
  wire [3:0] _GEN_747 = 5'hf == _T_867[4:0] ? 4'hc : _GEN_746; // @[Reg.scala 16:23]
  wire [3:0] _GEN_748 = 5'h10 == _T_867[4:0] ? 4'h0 : _GEN_747; // @[Reg.scala 16:23]
  wire [3:0] _GEN_749 = 5'h11 == _T_867[4:0] ? 4'h1 : _GEN_748; // @[Reg.scala 16:23]
  wire [3:0] _GEN_750 = 5'h12 == _T_867[4:0] ? 4'h2 : _GEN_749; // @[Reg.scala 16:23]
  wire [3:0] _GEN_751 = 5'h13 == _T_867[4:0] ? 4'h3 : _GEN_750; // @[Reg.scala 16:23]
  wire [3:0] _GEN_752 = 5'h14 == _T_867[4:0] ? 4'h4 : _GEN_751; // @[Reg.scala 16:23]
  wire [3:0] _GEN_753 = 5'h15 == _T_867[4:0] ? 4'h5 : _GEN_752; // @[Reg.scala 16:23]
  wire [3:0] _GEN_754 = 5'h16 == _T_867[4:0] ? 4'h6 : _GEN_753; // @[Reg.scala 16:23]
  wire [3:0] _GEN_755 = 5'h17 == _T_867[4:0] ? 4'h7 : _GEN_754; // @[Reg.scala 16:23]
  wire [3:0] _GEN_756 = 5'h18 == _T_867[4:0] ? 4'h0 : _GEN_755; // @[Reg.scala 16:23]
  wire [3:0] _GEN_757 = 5'h19 == _T_867[4:0] ? 4'h3 : _GEN_756; // @[Reg.scala 16:23]
  wire [3:0] _GEN_758 = 5'h1a == _T_867[4:0] ? 4'h6 : _GEN_757; // @[Reg.scala 16:23]
  wire [3:0] _GEN_759 = 5'h1b == _T_867[4:0] ? 4'h9 : _GEN_758; // @[Reg.scala 16:23]
  wire [3:0] _GEN_760 = 5'h1c == _T_867[4:0] ? 4'hb : _GEN_759; // @[Reg.scala 16:23]
  wire [3:0] _GEN_761 = 5'h1d == _T_867[4:0] ? 4'hd : _GEN_760; // @[Reg.scala 16:23]
  wire [3:0] _GEN_762 = 5'h1e == _T_867[4:0] ? 4'he : _GEN_761; // @[Reg.scala 16:23]
  wire [3:0] _GEN_763 = 5'h1f == _T_867[4:0] ? 4'hf : _GEN_762; // @[Reg.scala 16:23]
  reg [15:0] _T_877; // @[Reg.scala 15:16]
  reg [31:0] _RAND_89;
  reg [15:0] _T_878; // @[Reg.scala 15:16]
  reg [31:0] _RAND_90;
  reg [15:0] _T_879; // @[Reg.scala 15:16]
  reg [31:0] _RAND_91;
  reg [16:0] _T_881; // @[Reg.scala 15:16]
  reg [31:0] _RAND_92;
  reg [16:0] _T_883; // @[Reg.scala 15:16]
  reg [31:0] _RAND_93;
  reg [16:0] _T_885; // @[Reg.scala 15:16]
  reg [31:0] _RAND_94;
  wire [16:0] _GEN_949 = {{1{_T_877[15]}},_T_877}; // @[FixedPointTypeClass.scala 211:35]
  reg [32:0] _T_887; // @[Reg.scala 15:16]
  reg [63:0] _RAND_95;
  wire [34:0] _GEN_950 = {$signed(_T_887), 2'h0}; // @[FixedPointTypeClass.scala 20:58]
  wire [34:0] _T_890 = $signed(_GEN_950) + 35'sh1; // @[FixedPointTypeClass.scala 20:58]
  wire [33:0] _T_891 = _T_890[34:1]; // @[FixedPointTypeClass.scala 176:41]
  wire [16:0] _GEN_951 = {{1{_T_879[15]}},_T_879}; // @[FixedPointTypeClass.scala 211:35]
  reg [32:0] _T_893; // @[Reg.scala 15:16]
  reg [63:0] _RAND_96;
  wire [34:0] _GEN_952 = {$signed(_T_893), 2'h0}; // @[FixedPointTypeClass.scala 20:58]
  wire [34:0] _T_896 = $signed(_GEN_952) + 35'sh1; // @[FixedPointTypeClass.scala 20:58]
  wire [33:0] _T_897 = _T_896[34:1]; // @[FixedPointTypeClass.scala 176:41]
  wire [16:0] _GEN_953 = {{1{_T_878[15]}},_T_878}; // @[FixedPointTypeClass.scala 211:35]
  reg [32:0] _T_899; // @[Reg.scala 15:16]
  reg [63:0] _RAND_97;
  wire [34:0] _GEN_954 = {$signed(_T_899), 2'h0}; // @[FixedPointTypeClass.scala 20:58]
  wire [34:0] _T_902 = $signed(_GEN_954) + 35'sh1; // @[FixedPointTypeClass.scala 20:58]
  wire [33:0] _T_903 = _T_902[34:1]; // @[FixedPointTypeClass.scala 176:41]
  reg [34:0] _T_905; // @[Reg.scala 15:16]
  reg [63:0] _RAND_98;
  reg [34:0] _T_907; // @[Reg.scala 15:16]
  reg [63:0] _RAND_99;
  wire [34:0] _T_913 = $signed(_T_905) + 35'sh4000; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] _T_914 = _T_913[34:15]; // @[FixedPointTypeClass.scala 176:41]
  wire [34:0] _T_917 = $signed(_T_907) + 35'sh4000; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] _T_918 = _T_917[34:15]; // @[FixedPointTypeClass.scala 176:41]
  wire  _T_927 = 7'h4 == _T_71; // @[SDFChainRadix22.scala 234:23]
  wire [15:0] outputWires_3_imag = _T_918[15:0]; // @[SDFChainRadix22.scala 286:27 SDFChainRadix22.scala 306:19]
  wire [15:0] _GEN_841 = _T_927 ? $signed(io_in_bits_imag) : $signed(outputWires_3_imag); // @[SDFChainRadix22.scala 234:55]
  wire [15:0] outputWires_3_real = _T_914[15:0]; // @[SDFChainRadix22.scala 286:27 SDFChainRadix22.scala 306:19]
  wire [15:0] _GEN_842 = _T_927 ? $signed(io_in_bits_real) : $signed(outputWires_3_real); // @[SDFChainRadix22.scala 234:55]
  wire  _T_928 = sdf_stages_4_io_cntr < 7'h4; // @[SDFChainRadix22.scala 320:98]
  wire  _T_930 = sdf_stages_4_io_cntr < 7'h2; // @[SDFChainRadix22.scala 320:135]
  wire  _T_931 = _T_930 ? 1'h0 : 1'h1; // @[SDFChainRadix22.scala 320:122]
  reg  _T_933; // @[Reg.scala 15:16]
  reg [31:0] _RAND_100;
  wire [15:0] _T_939 = 16'sh0 - $signed(sdf_stages_4_io_out_real); // @[FixedPointTypeClass.scala 39:43]
  wire [15:0] _T_936_real = sdf_stages_4_io_out_imag; // @[SDFChainRadix22.scala 322:32 SDFChainRadix22.scala 325:29]
  reg [15:0] _T_945_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_101;
  reg [15:0] _T_945_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_102;
  reg [15:0] _T_948_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_103;
  reg [15:0] _T_948_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_104;
  reg [15:0] outputWires_4_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_105;
  reg [15:0] outputWires_4_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_106;
  wire  _T_957 = 7'h5 == _T_71; // @[SDFChainRadix22.scala 234:23]
  wire [15:0] _GEN_852 = _T_957 ? $signed(io_in_bits_imag) : $signed(outputWires_4_imag); // @[SDFChainRadix22.scala 234:55]
  wire [15:0] _GEN_853 = _T_957 ? $signed(io_in_bits_real) : $signed(outputWires_4_real); // @[SDFChainRadix22.scala 234:55]
  wire [6:0] _T_990 = _GEN_246 + 7'h1; // @[SDFChainRadix22.scala 276:83]
  wire [6:0] _T_994 = _T_990 - _T_301; // @[SDFChainRadix22.scala 276:89]
  reg [6:0] _T_996; // @[Reg.scala 15:16]
  reg [31:0] _RAND_107;
  reg [15:0] twiddles_5_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_108;
  reg [15:0] twiddles_5_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_109;
  wire [1:0] _GEN_881 = 3'h3 == _T_996[2:0] ? 2'h2 : 2'h0; // @[Reg.scala 16:23]
  wire [1:0] _GEN_882 = 3'h4 == _T_996[2:0] ? 2'h0 : _GEN_881; // @[Reg.scala 16:23]
  wire [1:0] _GEN_883 = 3'h5 == _T_996[2:0] ? 2'h1 : _GEN_882; // @[Reg.scala 16:23]
  wire [1:0] _GEN_884 = 3'h6 == _T_996[2:0] ? 2'h0 : _GEN_883; // @[Reg.scala 16:23]
  wire [1:0] _GEN_885 = 3'h7 == _T_996[2:0] ? 2'h3 : _GEN_884; // @[Reg.scala 16:23]
  reg [15:0] _T_1006; // @[Reg.scala 15:16]
  reg [31:0] _RAND_110;
  reg [15:0] _T_1007; // @[Reg.scala 15:16]
  reg [31:0] _RAND_111;
  reg [15:0] _T_1008; // @[Reg.scala 15:16]
  reg [31:0] _RAND_112;
  reg [16:0] _T_1010; // @[Reg.scala 15:16]
  reg [31:0] _RAND_113;
  reg [16:0] _T_1012; // @[Reg.scala 15:16]
  reg [31:0] _RAND_114;
  reg [16:0] _T_1014; // @[Reg.scala 15:16]
  reg [31:0] _RAND_115;
  wire [16:0] _GEN_957 = {{1{_T_1006[15]}},_T_1006}; // @[FixedPointTypeClass.scala 211:35]
  reg [32:0] _T_1016; // @[Reg.scala 15:16]
  reg [63:0] _RAND_116;
  wire [34:0] _GEN_958 = {$signed(_T_1016), 2'h0}; // @[FixedPointTypeClass.scala 20:58]
  wire [34:0] _T_1019 = $signed(_GEN_958) + 35'sh1; // @[FixedPointTypeClass.scala 20:58]
  wire [33:0] _T_1020 = _T_1019[34:1]; // @[FixedPointTypeClass.scala 176:41]
  wire [16:0] _GEN_959 = {{1{_T_1008[15]}},_T_1008}; // @[FixedPointTypeClass.scala 211:35]
  reg [32:0] _T_1022; // @[Reg.scala 15:16]
  reg [63:0] _RAND_117;
  wire [34:0] _GEN_960 = {$signed(_T_1022), 2'h0}; // @[FixedPointTypeClass.scala 20:58]
  wire [34:0] _T_1025 = $signed(_GEN_960) + 35'sh1; // @[FixedPointTypeClass.scala 20:58]
  wire [33:0] _T_1026 = _T_1025[34:1]; // @[FixedPointTypeClass.scala 176:41]
  wire [16:0] _GEN_961 = {{1{_T_1007[15]}},_T_1007}; // @[FixedPointTypeClass.scala 211:35]
  reg [32:0] _T_1028; // @[Reg.scala 15:16]
  reg [63:0] _RAND_118;
  wire [34:0] _GEN_962 = {$signed(_T_1028), 2'h0}; // @[FixedPointTypeClass.scala 20:58]
  wire [34:0] _T_1031 = $signed(_GEN_962) + 35'sh1; // @[FixedPointTypeClass.scala 20:58]
  wire [33:0] _T_1032 = _T_1031[34:1]; // @[FixedPointTypeClass.scala 176:41]
  reg [34:0] _T_1034; // @[Reg.scala 15:16]
  reg [63:0] _RAND_119;
  reg [34:0] _T_1036; // @[Reg.scala 15:16]
  reg [63:0] _RAND_120;
  wire [34:0] _T_1042 = $signed(_T_1034) + 35'sh4000; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] _T_1043 = _T_1042[34:15]; // @[FixedPointTypeClass.scala 176:41]
  wire [34:0] _T_1046 = $signed(_T_1036) + 35'sh4000; // @[FixedPointTypeClass.scala 20:58]
  wire [19:0] _T_1047 = _T_1046[34:15]; // @[FixedPointTypeClass.scala 176:41]
  wire  _T_1056 = 7'h6 == _T_71; // @[SDFChainRadix22.scala 234:23]
  wire [15:0] outputWires_5_imag = _T_1047[15:0]; // @[SDFChainRadix22.scala 286:27 SDFChainRadix22.scala 306:19]
  wire [15:0] _GEN_915 = _T_1056 ? $signed(io_in_bits_imag) : $signed(outputWires_5_imag); // @[SDFChainRadix22.scala 234:55]
  wire [15:0] outputWires_5_real = _T_1043[15:0]; // @[SDFChainRadix22.scala 286:27 SDFChainRadix22.scala 306:19]
  wire [15:0] _GEN_916 = _T_1056 ? $signed(io_in_bits_real) : $signed(outputWires_5_real); // @[SDFChainRadix22.scala 234:55]
  reg [15:0] _T_1059_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_121;
  reg [15:0] _T_1059_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_122;
  reg [15:0] _T_1062_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_123;
  reg [15:0] _T_1062_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_124;
  reg [15:0] outputWires_6_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_125;
  reg [15:0] outputWires_6_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_126;
  reg  _T_1067; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_127;
  reg  _T_1068; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_128;
  reg  _T_1069; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_129;
  reg  outValid; // @[SDFFFTUtil.scala 14:20]
  reg [31:0] _RAND_130;
  wire  _T_1070 = ~initialOutDone; // @[SDFChainRadix22.scala 361:33]
  reg  _T_1071; // @[Reg.scala 27:20]
  reg [31:0] _RAND_131;
  reg  _T_1072; // @[Reg.scala 27:20]
  reg [31:0] _RAND_132;
  reg  _T_1073; // @[Reg.scala 27:20]
  reg [31:0] _RAND_133;
  reg  _T_1074; // @[Reg.scala 27:20]
  reg [31:0] _RAND_134;
  wire  _T_1075 = state != 2'h2; // @[SDFChainRadix22.scala 361:127]
  wire  _T_1076 = io_out_ready & _T_1075; // @[SDFChainRadix22.scala 361:117]
  wire [29:0] _GEN_965 = {$signed(outQueue_io_deq_bits_imag), 14'h0}; // @[SDFChainRadix22.scala 375:33]
  wire [31:0] _GEN_937 = {{2{_GEN_965[29]}},_GEN_965}; // @[SDFChainRadix22.scala 375:33]
  wire [29:0] _GEN_966 = {$signed(outQueue_io_deq_bits_real), 14'h0}; // @[SDFChainRadix22.scala 375:33]
  wire [31:0] _GEN_938 = {{2{_GEN_966[29]}},_GEN_966}; // @[SDFChainRadix22.scala 375:33]
  wire [17:0] _GEN_967 = _GEN_938[31:14]; // @[SDFChainRadix22.scala 59:26 SDFChainRadix22.scala 376:20 SDFChainRadix22.scala 379:25]
  wire [17:0] _GEN_969 = _GEN_937[31:14]; // @[SDFChainRadix22.scala 59:26 SDFChainRadix22.scala 376:20 SDFChainRadix22.scala 380:25]
  SDFStageRadix22 sdf_stages_0 ( // @[SDFChainRadix22.scala 155:25]
    .clock(sdf_stages_0_clock),
    .reset(sdf_stages_0_reset),
    .io_in_real(sdf_stages_0_io_in_real),
    .io_in_imag(sdf_stages_0_io_in_imag),
    .io_out_real(sdf_stages_0_io_out_real),
    .io_out_imag(sdf_stages_0_io_out_imag),
    .io_cntr(sdf_stages_0_io_cntr),
    .io_en(sdf_stages_0_io_en)
  );
  SDFStageRadix22_1 sdf_stages_1 ( // @[SDFChainRadix22.scala 155:25]
    .clock(sdf_stages_1_clock),
    .reset(sdf_stages_1_reset),
    .io_in_real(sdf_stages_1_io_in_real),
    .io_in_imag(sdf_stages_1_io_in_imag),
    .io_out_real(sdf_stages_1_io_out_real),
    .io_out_imag(sdf_stages_1_io_out_imag),
    .io_cntr(sdf_stages_1_io_cntr),
    .io_en(sdf_stages_1_io_en)
  );
  SDFStageRadix22_2 sdf_stages_2 ( // @[SDFChainRadix22.scala 155:25]
    .clock(sdf_stages_2_clock),
    .reset(sdf_stages_2_reset),
    .io_in_real(sdf_stages_2_io_in_real),
    .io_in_imag(sdf_stages_2_io_in_imag),
    .io_out_real(sdf_stages_2_io_out_real),
    .io_out_imag(sdf_stages_2_io_out_imag),
    .io_cntr(sdf_stages_2_io_cntr),
    .io_en(sdf_stages_2_io_en)
  );
  SDFStageRadix22_3 sdf_stages_3 ( // @[SDFChainRadix22.scala 155:25]
    .clock(sdf_stages_3_clock),
    .reset(sdf_stages_3_reset),
    .io_in_real(sdf_stages_3_io_in_real),
    .io_in_imag(sdf_stages_3_io_in_imag),
    .io_out_real(sdf_stages_3_io_out_real),
    .io_out_imag(sdf_stages_3_io_out_imag),
    .io_cntr(sdf_stages_3_io_cntr),
    .io_en(sdf_stages_3_io_en)
  );
  SDFStageRadix22_4 sdf_stages_4 ( // @[SDFChainRadix22.scala 155:25]
    .clock(sdf_stages_4_clock),
    .reset(sdf_stages_4_reset),
    .io_in_real(sdf_stages_4_io_in_real),
    .io_in_imag(sdf_stages_4_io_in_imag),
    .io_out_real(sdf_stages_4_io_out_real),
    .io_out_imag(sdf_stages_4_io_out_imag),
    .io_cntr(sdf_stages_4_io_cntr),
    .io_en(sdf_stages_4_io_en)
  );
  SDFStageRadix22_5 sdf_stages_5 ( // @[SDFChainRadix22.scala 155:25]
    .clock(sdf_stages_5_clock),
    .reset(sdf_stages_5_reset),
    .io_in_real(sdf_stages_5_io_in_real),
    .io_in_imag(sdf_stages_5_io_in_imag),
    .io_out_real(sdf_stages_5_io_out_real),
    .io_out_imag(sdf_stages_5_io_out_imag),
    .io_cntr(sdf_stages_5_io_cntr),
    .io_en(sdf_stages_5_io_en)
  );
  SDFStageRadix22_6 sdf_stages_6 ( // @[SDFChainRadix22.scala 155:25]
    .clock(sdf_stages_6_clock),
    .reset(sdf_stages_6_reset),
    .io_in_real(sdf_stages_6_io_in_real),
    .io_in_imag(sdf_stages_6_io_in_imag),
    .io_out_real(sdf_stages_6_io_out_real),
    .io_out_imag(sdf_stages_6_io_out_imag),
    .io_cntr(sdf_stages_6_io_cntr),
    .io_en(sdf_stages_6_io_en)
  );
  Queue_10 outQueue ( // @[SDFChainRadix22.scala 356:25]
    .clock(outQueue_clock),
    .reset(outQueue_reset),
    .io_enq_ready(outQueue_io_enq_ready),
    .io_enq_valid(outQueue_io_enq_valid),
    .io_enq_bits_real(outQueue_io_enq_bits_real),
    .io_enq_bits_imag(outQueue_io_enq_bits_imag),
    .io_deq_ready(outQueue_io_deq_ready),
    .io_deq_valid(outQueue_io_deq_valid),
    .io_deq_bits_real(outQueue_io_deq_bits_real),
    .io_deq_bits_imag(outQueue_io_deq_bits_imag)
  );
  assign io_in_ready = _T_1074 | _T_1076; // @[SDFChainRadix22.scala 361:15]
  assign io_out_valid = outQueue_io_deq_valid; // @[SDFChainRadix22.scala 383:18]
  assign io_out_bits_real = _GEN_967[15:0]; // @[SDFChainRadix22.scala 382:17]
  assign io_out_bits_imag = _GEN_969[15:0]; // @[SDFChainRadix22.scala 382:17]
  assign io_lastOut = lastWait ? _T_67 : _T_69; // @[SDFChainRadix22.scala 389:14]
  assign io_busy = state == 2'h2; // @[SDFChainRadix22.scala 390:11]
  assign sdf_stages_0_clock = clock;
  assign sdf_stages_0_reset = reset;
  assign sdf_stages_0_io_in_real = activeStages_0 ? $signed(_GEN_262) : $signed(16'sh0); // @[SDFChainRadix22.scala 245:21 SDFChainRadix22.scala 248:21]
  assign sdf_stages_0_io_in_imag = activeStages_0 ? $signed(_GEN_261) : $signed(16'sh0); // @[SDFChainRadix22.scala 245:21 SDFChainRadix22.scala 248:21]
  assign sdf_stages_0_io_cntr = _GEN_176 - _T_211; // @[SDFChainRadix22.scala 217:16]
  assign sdf_stages_0_io_en = _T_202 ? 1'h0 : _GEN_169; // @[SDFChainRadix22.scala 216:14]
  assign sdf_stages_1_clock = clock;
  assign sdf_stages_1_reset = reset;
  assign sdf_stages_1_io_in_real = activeStages_1 ? $signed(_GEN_273) : $signed(16'sh0); // @[SDFChainRadix22.scala 245:21 SDFChainRadix22.scala 248:21]
  assign sdf_stages_1_io_in_imag = activeStages_1 ? $signed(_GEN_272) : $signed(16'sh0); // @[SDFChainRadix22.scala 245:21 SDFChainRadix22.scala 248:21]
  assign sdf_stages_1_io_cntr = {{1'd0}, _T_228[5:0]}; // @[SDFChainRadix22.scala 217:16]
  assign sdf_stages_1_io_en = _T_217 ? 1'h0 : _GEN_183; // @[SDFChainRadix22.scala 216:14]
  assign sdf_stages_2_clock = clock;
  assign sdf_stages_2_reset = reset;
  assign sdf_stages_2_io_in_real = activeStages_2 ? $signed(_GEN_696) : $signed(16'sh0); // @[SDFChainRadix22.scala 245:21 SDFChainRadix22.scala 248:21]
  assign sdf_stages_2_io_in_imag = activeStages_2 ? $signed(_GEN_695) : $signed(16'sh0); // @[SDFChainRadix22.scala 245:21 SDFChainRadix22.scala 248:21]
  assign sdf_stages_2_io_cntr = {{2'd0}, _T_243[4:0]}; // @[SDFChainRadix22.scala 217:16]
  assign sdf_stages_2_io_en = _T_232 ? 1'h0 : _GEN_197; // @[SDFChainRadix22.scala 216:14]
  assign sdf_stages_3_clock = clock;
  assign sdf_stages_3_reset = reset;
  assign sdf_stages_3_io_in_real = activeStages_3 ? $signed(_GEN_707) : $signed(16'sh0); // @[SDFChainRadix22.scala 245:21 SDFChainRadix22.scala 248:21]
  assign sdf_stages_3_io_in_imag = activeStages_3 ? $signed(_GEN_706) : $signed(16'sh0); // @[SDFChainRadix22.scala 245:21 SDFChainRadix22.scala 248:21]
  assign sdf_stages_3_io_cntr = {{3'd0}, _T_258[3:0]}; // @[SDFChainRadix22.scala 217:16]
  assign sdf_stages_3_io_en = _T_247 ? 1'h0 : _GEN_211; // @[SDFChainRadix22.scala 216:14]
  assign sdf_stages_4_clock = clock;
  assign sdf_stages_4_reset = reset;
  assign sdf_stages_4_io_in_real = activeStages_4 ? $signed(_GEN_842) : $signed(16'sh0); // @[SDFChainRadix22.scala 245:21 SDFChainRadix22.scala 248:21]
  assign sdf_stages_4_io_in_imag = activeStages_4 ? $signed(_GEN_841) : $signed(16'sh0); // @[SDFChainRadix22.scala 245:21 SDFChainRadix22.scala 248:21]
  assign sdf_stages_4_io_cntr = {{4'd0}, _T_273[2:0]}; // @[SDFChainRadix22.scala 217:16]
  assign sdf_stages_4_io_en = _T_262 ? 1'h0 : _GEN_225; // @[SDFChainRadix22.scala 216:14]
  assign sdf_stages_5_clock = clock;
  assign sdf_stages_5_reset = reset;
  assign sdf_stages_5_io_in_real = activeStages_5 ? $signed(_GEN_853) : $signed(16'sh0); // @[SDFChainRadix22.scala 245:21 SDFChainRadix22.scala 248:21]
  assign sdf_stages_5_io_in_imag = activeStages_5 ? $signed(_GEN_852) : $signed(16'sh0); // @[SDFChainRadix22.scala 245:21 SDFChainRadix22.scala 248:21]
  assign sdf_stages_5_io_cntr = {{5'd0}, _T_288[1:0]}; // @[SDFChainRadix22.scala 217:16]
  assign sdf_stages_5_io_en = _T_277 ? 1'h0 : _GEN_239; // @[SDFChainRadix22.scala 216:14]
  assign sdf_stages_6_clock = clock;
  assign sdf_stages_6_reset = reset;
  assign sdf_stages_6_io_in_real = activeStages_6 ? $signed(_GEN_916) : $signed(16'sh0); // @[SDFChainRadix22.scala 245:21 SDFChainRadix22.scala 248:21]
  assign sdf_stages_6_io_in_imag = activeStages_6 ? $signed(_GEN_915) : $signed(16'sh0); // @[SDFChainRadix22.scala 245:21 SDFChainRadix22.scala 248:21]
  assign sdf_stages_6_io_cntr = {{6'd0}, _T_303[0]}; // @[SDFChainRadix22.scala 217:16]
  assign sdf_stages_6_io_en = _T_292 ? 1'h0 : _GEN_253; // @[SDFChainRadix22.scala 216:14]
  assign outQueue_clock = clock;
  assign outQueue_reset = reset;
  assign outQueue_io_enq_valid = outValid; // @[SDFChainRadix22.scala 358:25]
  assign outQueue_io_enq_bits_real = outputWires_6_real; // @[SDFChainRadix22.scala 357:24]
  assign outQueue_io_enq_bits_imag = outputWires_6_imag; // @[SDFChainRadix22.scala 357:24]
  assign outQueue_io_deq_ready = io_out_ready; // @[SDFChainRadix22.scala 359:25]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regNumStages = _RAND_0[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  state = _RAND_1[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  initialOutDone = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  cnt = _RAND_3[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  cntValidOut = _RAND_4[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  lastWait = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  lastIndeed = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  initialInDone = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  initialInDonePrev = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_108 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_109 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_110 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  enableVector_1 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_113 = _RAND_13[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_114 = _RAND_14[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_115 = _RAND_15[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_116 = _RAND_16[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_118 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_119 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_120 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  enableVector_2 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_123 = _RAND_21[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_124 = _RAND_22[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_125 = _RAND_23[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_126 = _RAND_24[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_128 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_129 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T_130 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  enableVector_3 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_133 = _RAND_29[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_134 = _RAND_30[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T_135 = _RAND_31[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _T_136 = _RAND_32[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _T_138 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _T_139 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _T_140 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  enableVector_4 = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _T_143 = _RAND_37[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _T_144 = _RAND_38[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _T_145 = _RAND_39[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _T_146 = _RAND_40[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  _T_148 = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  _T_149 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  _T_150 = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  enableVector_5 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  _T_153 = _RAND_45[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  _T_154 = _RAND_46[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  _T_155 = _RAND_47[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  _T_156 = _RAND_48[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  _T_158 = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  _T_159 = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  _T_160 = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  enableVector_6 = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  _T_163 = _RAND_53[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  _T_164 = _RAND_54[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  _T_165 = _RAND_55[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  _T_166 = _RAND_56[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  _T_189 = _RAND_57[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  _T_316 = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  _T_328_real = _RAND_59[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  _T_328_imag = _RAND_60[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  _T_331_real = _RAND_61[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  _T_331_imag = _RAND_62[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  outputWires_0_real = _RAND_63[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  outputWires_0_imag = _RAND_64[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  _T_679 = _RAND_65[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  twiddles_1_real = _RAND_66[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  twiddles_1_imag = _RAND_67[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  _T_688 = _RAND_68[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  _T_689 = _RAND_69[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  _T_690 = _RAND_70[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  _T_692 = _RAND_71[16:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  _T_694 = _RAND_72[16:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  _T_696 = _RAND_73[16:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {2{`RANDOM}};
  _T_698 = _RAND_74[32:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {2{`RANDOM}};
  _T_704 = _RAND_75[32:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {2{`RANDOM}};
  _T_710 = _RAND_76[32:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {2{`RANDOM}};
  _T_716 = _RAND_77[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {2{`RANDOM}};
  _T_718 = _RAND_78[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  _T_744 = _RAND_79[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  _T_756_real = _RAND_80[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  _T_756_imag = _RAND_81[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  _T_759_real = _RAND_82[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  _T_759_imag = _RAND_83[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  outputWires_2_real = _RAND_84[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  outputWires_2_imag = _RAND_85[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  _T_867 = _RAND_86[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  twiddles_3_real = _RAND_87[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  twiddles_3_imag = _RAND_88[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  _T_877 = _RAND_89[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  _T_878 = _RAND_90[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  _T_879 = _RAND_91[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  _T_881 = _RAND_92[16:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  _T_883 = _RAND_93[16:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  _T_885 = _RAND_94[16:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {2{`RANDOM}};
  _T_887 = _RAND_95[32:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {2{`RANDOM}};
  _T_893 = _RAND_96[32:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {2{`RANDOM}};
  _T_899 = _RAND_97[32:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {2{`RANDOM}};
  _T_905 = _RAND_98[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {2{`RANDOM}};
  _T_907 = _RAND_99[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  _T_933 = _RAND_100[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  _T_945_real = _RAND_101[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  _T_945_imag = _RAND_102[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  _T_948_real = _RAND_103[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  _T_948_imag = _RAND_104[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  outputWires_4_real = _RAND_105[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  outputWires_4_imag = _RAND_106[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  _T_996 = _RAND_107[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  twiddles_5_real = _RAND_108[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  twiddles_5_imag = _RAND_109[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  _T_1006 = _RAND_110[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  _T_1007 = _RAND_111[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  _T_1008 = _RAND_112[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  _T_1010 = _RAND_113[16:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  _T_1012 = _RAND_114[16:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  _T_1014 = _RAND_115[16:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {2{`RANDOM}};
  _T_1016 = _RAND_116[32:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {2{`RANDOM}};
  _T_1022 = _RAND_117[32:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {2{`RANDOM}};
  _T_1028 = _RAND_118[32:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {2{`RANDOM}};
  _T_1034 = _RAND_119[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {2{`RANDOM}};
  _T_1036 = _RAND_120[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  _T_1059_real = _RAND_121[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  _T_1059_imag = _RAND_122[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  _T_1062_real = _RAND_123[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  _T_1062_imag = _RAND_124[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  outputWires_6_real = _RAND_125[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  outputWires_6_imag = _RAND_126[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  _T_1067 = _RAND_127[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  _T_1068 = _RAND_128[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{`RANDOM}};
  _T_1069 = _RAND_129[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{`RANDOM}};
  outValid = _RAND_130[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{`RANDOM}};
  _T_1071 = _RAND_131[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{`RANDOM}};
  _T_1072 = _RAND_132[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{`RANDOM}};
  _T_1073 = _RAND_133[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{`RANDOM}};
  _T_1074 = _RAND_134[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      regNumStages <= 7'h7;
    end else if (_T_42) begin
      regNumStages <= io_fftSize;
    end
    if (reset) begin
      state <= 2'h0;
    end else if (_T_42) begin
      if (_T_41) begin
        state <= 2'h1;
      end
    end else if (_T_45) begin
      if (fireLast) begin
        state <= 2'h2;
      end
    end else if (_T_46) begin
      if (io_lastOut) begin
        state <= 2'h0;
      end
    end
    if (reset) begin
      initialOutDone <= 1'h0;
    end else begin
      initialOutDone <= _GEN_160;
    end
    if (reset) begin
      cnt <= 8'h0;
    end else if (_T_51) begin
      cnt <= 8'h0;
    end else if (enableInit) begin
      cnt <= _T_106;
    end
    if (reset) begin
      cntValidOut <= 7'h0;
    end else if (_T_61) begin
      cntValidOut <= 7'h0;
    end else if (_T_50) begin
      cntValidOut <= _T_64;
    end
    if (reset) begin
      lastWait <= 1'h0;
    end else if (_T_51) begin
      lastWait <= 1'h0;
    end else begin
      lastWait <= _GEN_17;
    end
    if (reset) begin
      lastIndeed <= 1'h0;
    end else if (_T_51) begin
      lastIndeed <= 1'h0;
    end else begin
      lastIndeed <= _GEN_21;
    end
    if (reset) begin
      initialInDone <= 1'h0;
    end else if (_T_51) begin
      initialInDone <= 1'h0;
    end else begin
      initialInDone <= _GEN_15;
    end
    if (reset) begin
      initialInDonePrev <= 1'h0;
    end else begin
      initialInDonePrev <= initialInDone;
    end
    if (reset) begin
      _T_108 <= 1'h0;
    end else if (_T_51) begin
      _T_108 <= 1'h0;
    end else begin
      _T_108 <= enableInit;
    end
    if (reset) begin
      _T_109 <= 1'h0;
    end else if (_T_51) begin
      _T_109 <= 1'h0;
    end else begin
      _T_109 <= _T_108;
    end
    if (reset) begin
      _T_110 <= 1'h0;
    end else if (_T_51) begin
      _T_110 <= 1'h0;
    end else begin
      _T_110 <= _T_109;
    end
    if (reset) begin
      enableVector_1 <= 1'h0;
    end else if (_T_51) begin
      enableVector_1 <= 1'h0;
    end else begin
      enableVector_1 <= _T_110;
    end
    if (reset) begin
      _T_113 <= 8'h0;
    end else if (_T_51) begin
      _T_113 <= 8'h0;
    end else begin
      _T_113 <= cnt;
    end
    if (reset) begin
      _T_114 <= 8'h0;
    end else if (_T_51) begin
      _T_114 <= 8'h0;
    end else begin
      _T_114 <= _T_113;
    end
    if (reset) begin
      _T_115 <= 8'h0;
    end else if (_T_51) begin
      _T_115 <= 8'h0;
    end else begin
      _T_115 <= _T_114;
    end
    if (reset) begin
      _T_116 <= 8'h0;
    end else if (_T_51) begin
      _T_116 <= 8'h0;
    end else begin
      _T_116 <= _T_115;
    end
    if (reset) begin
      _T_118 <= 1'h0;
    end else if (_T_51) begin
      _T_118 <= 1'h0;
    end else begin
      _T_118 <= enableVector_1;
    end
    if (reset) begin
      _T_119 <= 1'h0;
    end else if (_T_51) begin
      _T_119 <= 1'h0;
    end else begin
      _T_119 <= _T_118;
    end
    if (reset) begin
      _T_120 <= 1'h0;
    end else if (_T_51) begin
      _T_120 <= 1'h0;
    end else begin
      _T_120 <= _T_119;
    end
    if (reset) begin
      enableVector_2 <= 1'h0;
    end else if (_T_51) begin
      enableVector_2 <= 1'h0;
    end else begin
      enableVector_2 <= _T_120;
    end
    if (reset) begin
      _T_123 <= 8'h0;
    end else if (_T_51) begin
      _T_123 <= 8'h0;
    end else begin
      _T_123 <= _T_116;
    end
    if (reset) begin
      _T_124 <= 8'h0;
    end else if (_T_51) begin
      _T_124 <= 8'h0;
    end else begin
      _T_124 <= _T_123;
    end
    if (reset) begin
      _T_125 <= 8'h0;
    end else if (_T_51) begin
      _T_125 <= 8'h0;
    end else begin
      _T_125 <= _T_124;
    end
    if (reset) begin
      _T_126 <= 8'h0;
    end else if (_T_51) begin
      _T_126 <= 8'h0;
    end else begin
      _T_126 <= _T_125;
    end
    if (reset) begin
      _T_128 <= 1'h0;
    end else if (_T_51) begin
      _T_128 <= 1'h0;
    end else begin
      _T_128 <= enableVector_2;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else if (_T_51) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_128;
    end
    if (reset) begin
      _T_130 <= 1'h0;
    end else if (_T_51) begin
      _T_130 <= 1'h0;
    end else begin
      _T_130 <= _T_129;
    end
    if (reset) begin
      enableVector_3 <= 1'h0;
    end else if (_T_51) begin
      enableVector_3 <= 1'h0;
    end else begin
      enableVector_3 <= _T_130;
    end
    if (reset) begin
      _T_133 <= 8'h0;
    end else if (_T_51) begin
      _T_133 <= 8'h0;
    end else begin
      _T_133 <= _T_126;
    end
    if (reset) begin
      _T_134 <= 8'h0;
    end else if (_T_51) begin
      _T_134 <= 8'h0;
    end else begin
      _T_134 <= _T_133;
    end
    if (reset) begin
      _T_135 <= 8'h0;
    end else if (_T_51) begin
      _T_135 <= 8'h0;
    end else begin
      _T_135 <= _T_134;
    end
    if (reset) begin
      _T_136 <= 8'h0;
    end else if (_T_51) begin
      _T_136 <= 8'h0;
    end else begin
      _T_136 <= _T_135;
    end
    if (reset) begin
      _T_138 <= 1'h0;
    end else if (_T_51) begin
      _T_138 <= 1'h0;
    end else begin
      _T_138 <= enableVector_3;
    end
    if (reset) begin
      _T_139 <= 1'h0;
    end else if (_T_51) begin
      _T_139 <= 1'h0;
    end else begin
      _T_139 <= _T_138;
    end
    if (reset) begin
      _T_140 <= 1'h0;
    end else if (_T_51) begin
      _T_140 <= 1'h0;
    end else begin
      _T_140 <= _T_139;
    end
    if (reset) begin
      enableVector_4 <= 1'h0;
    end else if (_T_51) begin
      enableVector_4 <= 1'h0;
    end else begin
      enableVector_4 <= _T_140;
    end
    if (reset) begin
      _T_143 <= 8'h0;
    end else if (_T_51) begin
      _T_143 <= 8'h0;
    end else begin
      _T_143 <= _T_136;
    end
    if (reset) begin
      _T_144 <= 8'h0;
    end else if (_T_51) begin
      _T_144 <= 8'h0;
    end else begin
      _T_144 <= _T_143;
    end
    if (reset) begin
      _T_145 <= 8'h0;
    end else if (_T_51) begin
      _T_145 <= 8'h0;
    end else begin
      _T_145 <= _T_144;
    end
    if (reset) begin
      _T_146 <= 8'h0;
    end else if (_T_51) begin
      _T_146 <= 8'h0;
    end else begin
      _T_146 <= _T_145;
    end
    if (reset) begin
      _T_148 <= 1'h0;
    end else if (_T_51) begin
      _T_148 <= 1'h0;
    end else begin
      _T_148 <= enableVector_4;
    end
    if (reset) begin
      _T_149 <= 1'h0;
    end else if (_T_51) begin
      _T_149 <= 1'h0;
    end else begin
      _T_149 <= _T_148;
    end
    if (reset) begin
      _T_150 <= 1'h0;
    end else if (_T_51) begin
      _T_150 <= 1'h0;
    end else begin
      _T_150 <= _T_149;
    end
    if (reset) begin
      enableVector_5 <= 1'h0;
    end else if (_T_51) begin
      enableVector_5 <= 1'h0;
    end else begin
      enableVector_5 <= _T_150;
    end
    if (reset) begin
      _T_153 <= 8'h0;
    end else if (_T_51) begin
      _T_153 <= 8'h0;
    end else begin
      _T_153 <= _T_146;
    end
    if (reset) begin
      _T_154 <= 8'h0;
    end else if (_T_51) begin
      _T_154 <= 8'h0;
    end else begin
      _T_154 <= _T_153;
    end
    if (reset) begin
      _T_155 <= 8'h0;
    end else if (_T_51) begin
      _T_155 <= 8'h0;
    end else begin
      _T_155 <= _T_154;
    end
    if (reset) begin
      _T_156 <= 8'h0;
    end else if (_T_51) begin
      _T_156 <= 8'h0;
    end else begin
      _T_156 <= _T_155;
    end
    if (reset) begin
      _T_158 <= 1'h0;
    end else if (_T_51) begin
      _T_158 <= 1'h0;
    end else begin
      _T_158 <= enableVector_5;
    end
    if (reset) begin
      _T_159 <= 1'h0;
    end else if (_T_51) begin
      _T_159 <= 1'h0;
    end else begin
      _T_159 <= _T_158;
    end
    if (reset) begin
      _T_160 <= 1'h0;
    end else if (_T_51) begin
      _T_160 <= 1'h0;
    end else begin
      _T_160 <= _T_159;
    end
    if (reset) begin
      enableVector_6 <= 1'h0;
    end else if (_T_51) begin
      enableVector_6 <= 1'h0;
    end else begin
      enableVector_6 <= _T_160;
    end
    if (reset) begin
      _T_163 <= 8'h0;
    end else if (_T_51) begin
      _T_163 <= 8'h0;
    end else begin
      _T_163 <= _T_156;
    end
    if (reset) begin
      _T_164 <= 8'h0;
    end else if (_T_51) begin
      _T_164 <= 8'h0;
    end else begin
      _T_164 <= _T_163;
    end
    if (reset) begin
      _T_165 <= 8'h0;
    end else if (_T_51) begin
      _T_165 <= 8'h0;
    end else begin
      _T_165 <= _T_164;
    end
    if (reset) begin
      _T_166 <= 8'h0;
    end else if (_T_51) begin
      _T_166 <= 8'h0;
    end else begin
      _T_166 <= _T_165;
    end
    _T_189 <= _T_41 | _T_103;
    _T_316 <= _T_311 & _T_314;
    if (_T_316) begin
      _T_328_real <= _T_319_real;
    end else begin
      _T_328_real <= sdf_stages_0_io_out_real;
    end
    if (_T_316) begin
      _T_328_imag <= _T_322;
    end else begin
      _T_328_imag <= sdf_stages_0_io_out_imag;
    end
    _T_331_real <= _T_328_real;
    _T_331_imag <= _T_328_imag;
    outputWires_0_real <= _T_331_real;
    outputWires_0_imag <= _T_331_imag;
    if (_GEN_183) begin
      _T_679 <= _T_677;
    end
    if (6'h3f == _GEN_425) begin
      twiddles_1_real <= -16'sh964;
    end else if (6'h3e == _GEN_425) begin
      twiddles_1_real <= -16'sh1294;
    end else if (6'h3d == _GEN_425) begin
      twiddles_1_real <= -16'sh1b5d;
    end else if (6'h3c == _GEN_425) begin
      twiddles_1_real <= -16'sh238e;
    end else if (6'h3b == _GEN_425) begin
      twiddles_1_real <= -16'sh2afb;
    end else if (6'h3a == _GEN_425) begin
      twiddles_1_real <= -16'sh3179;
    end else if (6'h39 == _GEN_425) begin
      twiddles_1_real <= -16'sh36e5;
    end else if (6'h38 == _GEN_425) begin
      twiddles_1_real <= -16'sh3b21;
    end else if (6'h37 == _GEN_425) begin
      twiddles_1_real <= -16'sh3e15;
    end else if (6'h36 == _GEN_425) begin
      twiddles_1_real <= -16'sh3fb1;
    end else if (6'h35 == _GEN_425) begin
      twiddles_1_real <= -16'sh3fec;
    end else if (6'h34 == _GEN_425) begin
      twiddles_1_real <= -16'sh3fb1;
    end else if (6'h33 == _GEN_425) begin
      twiddles_1_real <= -16'sh3ec5;
    end else if (6'h32 == _GEN_425) begin
      twiddles_1_real <= -16'sh3d3f;
    end else if (6'h31 == _GEN_425) begin
      twiddles_1_real <= -16'sh3c42;
    end else if (6'h30 == _GEN_425) begin
      twiddles_1_real <= -16'sh3b21;
    end else if (6'h2f == _GEN_425) begin
      twiddles_1_real <= -16'sh3871;
    end else if (6'h2e == _GEN_425) begin
      twiddles_1_real <= -16'sh3537;
    end else if (6'h2d == _GEN_425) begin
      twiddles_1_real <= -16'sh3368;
    end else if (6'h2c == _GEN_425) begin
      twiddles_1_real <= -16'sh3179;
    end else if (6'h2b == _GEN_425) begin
      twiddles_1_real <= -16'sh2d41;
    end else if (6'h2a == _GEN_425) begin
      twiddles_1_real <= -16'sh289a;
    end else if (6'h29 == _GEN_425) begin
      twiddles_1_real <= -16'sh2620;
    end else if (6'h28 == _GEN_425) begin
      twiddles_1_real <= -16'sh238e;
    end else if (6'h27 == _GEN_425) begin
      twiddles_1_real <= -16'sh1e2b;
    end else if (6'h26 == _GEN_425) begin
      twiddles_1_real <= -16'sh187e;
    end else if (6'h25 == _GEN_425) begin
      twiddles_1_real <= -16'sh1590;
    end else if (6'h24 == _GEN_425) begin
      twiddles_1_real <= -16'sh1294;
    end else if (6'h23 == _GEN_425) begin
      twiddles_1_real <= -16'shc7c;
    end else if (6'h22 == _GEN_425) begin
      twiddles_1_real <= -16'sh646;
    end else if (6'h21 == _GEN_425) begin
      twiddles_1_real <= -16'sh324;
    end else if (6'h20 == _GEN_425) begin
      twiddles_1_real <= 16'sh0;
    end else if (6'h1f == _GEN_425) begin
      twiddles_1_real <= 16'sh324;
    end else if (6'h1e == _GEN_425) begin
      twiddles_1_real <= 16'sh646;
    end else if (6'h1d == _GEN_425) begin
      twiddles_1_real <= 16'sh964;
    end else if (6'h1c == _GEN_425) begin
      twiddles_1_real <= 16'shc7c;
    end else if (6'h1b == _GEN_425) begin
      twiddles_1_real <= 16'shf8d;
    end else if (6'h1a == _GEN_425) begin
      twiddles_1_real <= 16'sh1294;
    end else if (6'h19 == _GEN_425) begin
      twiddles_1_real <= 16'sh1590;
    end else if (6'h18 == _GEN_425) begin
      twiddles_1_real <= 16'sh187e;
    end else if (6'h17 == _GEN_425) begin
      twiddles_1_real <= 16'sh1b5d;
    end else if (6'h16 == _GEN_425) begin
      twiddles_1_real <= 16'sh1e2b;
    end else if (6'h15 == _GEN_425) begin
      twiddles_1_real <= 16'sh20e7;
    end else if (6'h14 == _GEN_425) begin
      twiddles_1_real <= 16'sh238e;
    end else if (6'h13 == _GEN_425) begin
      twiddles_1_real <= 16'sh2620;
    end else if (6'h12 == _GEN_425) begin
      twiddles_1_real <= 16'sh289a;
    end else if (6'h11 == _GEN_425) begin
      twiddles_1_real <= 16'sh2afb;
    end else if (6'h10 == _GEN_425) begin
      twiddles_1_real <= 16'sh2d41;
    end else if (6'hf == _GEN_425) begin
      twiddles_1_real <= 16'sh2f6c;
    end else if (6'he == _GEN_425) begin
      twiddles_1_real <= 16'sh3179;
    end else if (6'hd == _GEN_425) begin
      twiddles_1_real <= 16'sh3368;
    end else if (6'hc == _GEN_425) begin
      twiddles_1_real <= 16'sh3537;
    end else if (6'hb == _GEN_425) begin
      twiddles_1_real <= 16'sh36e5;
    end else if (6'ha == _GEN_425) begin
      twiddles_1_real <= 16'sh3871;
    end else if (6'h9 == _GEN_425) begin
      twiddles_1_real <= 16'sh39db;
    end else if (6'h8 == _GEN_425) begin
      twiddles_1_real <= 16'sh3b21;
    end else if (6'h7 == _GEN_425) begin
      twiddles_1_real <= 16'sh3c42;
    end else if (6'h6 == _GEN_425) begin
      twiddles_1_real <= 16'sh3d3f;
    end else if (6'h5 == _GEN_425) begin
      twiddles_1_real <= 16'sh3e15;
    end else if (6'h4 == _GEN_425) begin
      twiddles_1_real <= 16'sh3ec5;
    end else if (6'h3 == _GEN_425) begin
      twiddles_1_real <= 16'sh3f4f;
    end else if (6'h2 == _GEN_425) begin
      twiddles_1_real <= 16'sh3fb1;
    end else if (6'h1 == _GEN_425) begin
      twiddles_1_real <= 16'sh3fec;
    end else begin
      twiddles_1_real <= 16'sh4000;
    end
    if (6'h3f == _GEN_425) begin
      twiddles_1_imag <= 16'sh3f4f;
    end else if (6'h3e == _GEN_425) begin
      twiddles_1_imag <= 16'sh3d3f;
    end else if (6'h3d == _GEN_425) begin
      twiddles_1_imag <= 16'sh39db;
    end else if (6'h3c == _GEN_425) begin
      twiddles_1_imag <= 16'sh3537;
    end else if (6'h3b == _GEN_425) begin
      twiddles_1_imag <= 16'sh2f6c;
    end else if (6'h3a == _GEN_425) begin
      twiddles_1_imag <= 16'sh289a;
    end else if (6'h39 == _GEN_425) begin
      twiddles_1_imag <= 16'sh20e7;
    end else if (6'h38 == _GEN_425) begin
      twiddles_1_imag <= 16'sh187e;
    end else if (6'h37 == _GEN_425) begin
      twiddles_1_imag <= 16'shf8d;
    end else if (6'h36 == _GEN_425) begin
      twiddles_1_imag <= 16'sh646;
    end else if (6'h35 == _GEN_425) begin
      twiddles_1_imag <= -16'sh324;
    end else if (6'h34 == _GEN_425) begin
      twiddles_1_imag <= -16'sh646;
    end else if (6'h33 == _GEN_425) begin
      twiddles_1_imag <= -16'shc7c;
    end else if (6'h32 == _GEN_425) begin
      twiddles_1_imag <= -16'sh1294;
    end else if (6'h31 == _GEN_425) begin
      twiddles_1_imag <= -16'sh1590;
    end else if (6'h30 == _GEN_425) begin
      twiddles_1_imag <= -16'sh187e;
    end else if (6'h2f == _GEN_425) begin
      twiddles_1_imag <= -16'sh1e2b;
    end else if (6'h2e == _GEN_425) begin
      twiddles_1_imag <= -16'sh238e;
    end else if (6'h2d == _GEN_425) begin
      twiddles_1_imag <= -16'sh2620;
    end else if (6'h2c == _GEN_425) begin
      twiddles_1_imag <= -16'sh289a;
    end else if (6'h2b == _GEN_425) begin
      twiddles_1_imag <= -16'sh2d41;
    end else if (6'h2a == _GEN_425) begin
      twiddles_1_imag <= -16'sh3179;
    end else if (6'h29 == _GEN_425) begin
      twiddles_1_imag <= -16'sh3368;
    end else if (6'h28 == _GEN_425) begin
      twiddles_1_imag <= -16'sh3537;
    end else if (6'h27 == _GEN_425) begin
      twiddles_1_imag <= -16'sh3871;
    end else if (6'h26 == _GEN_425) begin
      twiddles_1_imag <= -16'sh3b21;
    end else if (6'h25 == _GEN_425) begin
      twiddles_1_imag <= -16'sh3c42;
    end else if (6'h24 == _GEN_425) begin
      twiddles_1_imag <= -16'sh3d3f;
    end else if (6'h23 == _GEN_425) begin
      twiddles_1_imag <= -16'sh3ec5;
    end else if (6'h22 == _GEN_425) begin
      twiddles_1_imag <= -16'sh3fb1;
    end else if (6'h21 == _GEN_425) begin
      twiddles_1_imag <= -16'sh3fec;
    end else if (6'h20 == _GEN_425) begin
      twiddles_1_imag <= -16'sh4000;
    end else if (6'h1f == _GEN_425) begin
      twiddles_1_imag <= -16'sh3fec;
    end else if (6'h1e == _GEN_425) begin
      twiddles_1_imag <= -16'sh3fb1;
    end else if (6'h1d == _GEN_425) begin
      twiddles_1_imag <= -16'sh3f4f;
    end else if (6'h1c == _GEN_425) begin
      twiddles_1_imag <= -16'sh3ec5;
    end else if (6'h1b == _GEN_425) begin
      twiddles_1_imag <= -16'sh3e15;
    end else if (6'h1a == _GEN_425) begin
      twiddles_1_imag <= -16'sh3d3f;
    end else if (6'h19 == _GEN_425) begin
      twiddles_1_imag <= -16'sh3c42;
    end else if (6'h18 == _GEN_425) begin
      twiddles_1_imag <= -16'sh3b21;
    end else if (6'h17 == _GEN_425) begin
      twiddles_1_imag <= -16'sh39db;
    end else if (6'h16 == _GEN_425) begin
      twiddles_1_imag <= -16'sh3871;
    end else if (6'h15 == _GEN_425) begin
      twiddles_1_imag <= -16'sh36e5;
    end else if (6'h14 == _GEN_425) begin
      twiddles_1_imag <= -16'sh3537;
    end else if (6'h13 == _GEN_425) begin
      twiddles_1_imag <= -16'sh3368;
    end else if (6'h12 == _GEN_425) begin
      twiddles_1_imag <= -16'sh3179;
    end else if (6'h11 == _GEN_425) begin
      twiddles_1_imag <= -16'sh2f6c;
    end else if (6'h10 == _GEN_425) begin
      twiddles_1_imag <= -16'sh2d41;
    end else if (6'hf == _GEN_425) begin
      twiddles_1_imag <= -16'sh2afb;
    end else if (6'he == _GEN_425) begin
      twiddles_1_imag <= -16'sh289a;
    end else if (6'hd == _GEN_425) begin
      twiddles_1_imag <= -16'sh2620;
    end else if (6'hc == _GEN_425) begin
      twiddles_1_imag <= -16'sh238e;
    end else if (6'hb == _GEN_425) begin
      twiddles_1_imag <= -16'sh20e7;
    end else if (6'ha == _GEN_425) begin
      twiddles_1_imag <= -16'sh1e2b;
    end else if (6'h9 == _GEN_425) begin
      twiddles_1_imag <= -16'sh1b5d;
    end else if (6'h8 == _GEN_425) begin
      twiddles_1_imag <= -16'sh187e;
    end else if (6'h7 == _GEN_425) begin
      twiddles_1_imag <= -16'sh1590;
    end else if (6'h6 == _GEN_425) begin
      twiddles_1_imag <= -16'sh1294;
    end else if (6'h5 == _GEN_425) begin
      twiddles_1_imag <= -16'shf8d;
    end else if (6'h4 == _GEN_425) begin
      twiddles_1_imag <= -16'shc7c;
    end else if (6'h3 == _GEN_425) begin
      twiddles_1_imag <= -16'sh964;
    end else if (6'h2 == _GEN_425) begin
      twiddles_1_imag <= -16'sh646;
    end else if (6'h1 == _GEN_425) begin
      twiddles_1_imag <= -16'sh324;
    end else begin
      twiddles_1_imag <= 16'sh0;
    end
    _T_688 <= sdf_stages_1_io_out_real;
    _T_689 <= twiddles_1_real;
    _T_690 <= twiddles_1_imag;
    _T_692 <= $signed(twiddles_1_real) + $signed(twiddles_1_imag);
    _T_694 <= $signed(sdf_stages_1_io_out_real) + $signed(sdf_stages_1_io_out_imag);
    _T_696 <= $signed(sdf_stages_1_io_out_imag) - $signed(sdf_stages_1_io_out_real);
    _T_698 <= $signed(_GEN_941) * $signed(_T_692);
    _T_704 <= $signed(_T_694) * $signed(_GEN_943);
    _T_710 <= $signed(_T_696) * $signed(_GEN_945);
    _T_716 <= $signed(_T_702) - $signed(_T_708);
    _T_718 <= $signed(_T_702) + $signed(_T_714);
    _T_744 <= _T_739 & _T_742;
    if (_T_744) begin
      _T_756_real <= _T_747_real;
    end else begin
      _T_756_real <= sdf_stages_2_io_out_real;
    end
    if (_T_744) begin
      _T_756_imag <= _T_750;
    end else begin
      _T_756_imag <= sdf_stages_2_io_out_imag;
    end
    _T_759_real <= _T_756_real;
    _T_759_imag <= _T_756_imag;
    outputWires_2_real <= _T_759_real;
    outputWires_2_imag <= _T_759_imag;
    if (_GEN_211) begin
      _T_867 <= _T_865;
    end
    if (4'hf == _GEN_763) begin
      twiddles_3_real <= -16'sh238e;
    end else if (4'he == _GEN_763) begin
      twiddles_3_real <= -16'sh3b21;
    end else if (4'hd == _GEN_763) begin
      twiddles_3_real <= -16'sh3ec5;
    end else if (4'hc == _GEN_763) begin
      twiddles_3_real <= -16'sh3b21;
    end else if (4'hb == _GEN_763) begin
      twiddles_3_real <= -16'sh2d41;
    end else if (4'ha == _GEN_763) begin
      twiddles_3_real <= -16'sh187e;
    end else if (4'h9 == _GEN_763) begin
      twiddles_3_real <= -16'shc7c;
    end else if (4'h8 == _GEN_763) begin
      twiddles_3_real <= 16'sh0;
    end else if (4'h7 == _GEN_763) begin
      twiddles_3_real <= 16'shc7c;
    end else if (4'h6 == _GEN_763) begin
      twiddles_3_real <= 16'sh187e;
    end else if (4'h5 == _GEN_763) begin
      twiddles_3_real <= 16'sh238e;
    end else if (4'h4 == _GEN_763) begin
      twiddles_3_real <= 16'sh2d41;
    end else if (4'h3 == _GEN_763) begin
      twiddles_3_real <= 16'sh3537;
    end else if (4'h2 == _GEN_763) begin
      twiddles_3_real <= 16'sh3b21;
    end else if (4'h1 == _GEN_763) begin
      twiddles_3_real <= 16'sh3ec5;
    end else begin
      twiddles_3_real <= 16'sh4000;
    end
    if (4'hf == _GEN_763) begin
      twiddles_3_imag <= 16'sh3537;
    end else if (4'he == _GEN_763) begin
      twiddles_3_imag <= 16'sh187e;
    end else if (4'hd == _GEN_763) begin
      twiddles_3_imag <= -16'shc7c;
    end else if (4'hc == _GEN_763) begin
      twiddles_3_imag <= -16'sh187e;
    end else if (4'hb == _GEN_763) begin
      twiddles_3_imag <= -16'sh2d41;
    end else if (4'ha == _GEN_763) begin
      twiddles_3_imag <= -16'sh3b21;
    end else if (4'h9 == _GEN_763) begin
      twiddles_3_imag <= -16'sh3ec5;
    end else if (4'h8 == _GEN_763) begin
      twiddles_3_imag <= -16'sh4000;
    end else if (4'h7 == _GEN_763) begin
      twiddles_3_imag <= -16'sh3ec5;
    end else if (4'h6 == _GEN_763) begin
      twiddles_3_imag <= -16'sh3b21;
    end else if (4'h5 == _GEN_763) begin
      twiddles_3_imag <= -16'sh3537;
    end else if (4'h4 == _GEN_763) begin
      twiddles_3_imag <= -16'sh2d41;
    end else if (4'h3 == _GEN_763) begin
      twiddles_3_imag <= -16'sh238e;
    end else if (4'h2 == _GEN_763) begin
      twiddles_3_imag <= -16'sh187e;
    end else if (4'h1 == _GEN_763) begin
      twiddles_3_imag <= -16'shc7c;
    end else begin
      twiddles_3_imag <= 16'sh0;
    end
    _T_877 <= sdf_stages_3_io_out_real;
    _T_878 <= twiddles_3_real;
    _T_879 <= twiddles_3_imag;
    _T_881 <= $signed(twiddles_3_real) + $signed(twiddles_3_imag);
    _T_883 <= $signed(sdf_stages_3_io_out_real) + $signed(sdf_stages_3_io_out_imag);
    _T_885 <= $signed(sdf_stages_3_io_out_imag) - $signed(sdf_stages_3_io_out_real);
    _T_887 <= $signed(_GEN_949) * $signed(_T_881);
    _T_893 <= $signed(_T_883) * $signed(_GEN_951);
    _T_899 <= $signed(_T_885) * $signed(_GEN_953);
    _T_905 <= $signed(_T_891) - $signed(_T_897);
    _T_907 <= $signed(_T_891) + $signed(_T_903);
    _T_933 <= _T_928 & _T_931;
    if (_T_933) begin
      _T_945_real <= _T_936_real;
    end else begin
      _T_945_real <= sdf_stages_4_io_out_real;
    end
    if (_T_933) begin
      _T_945_imag <= _T_939;
    end else begin
      _T_945_imag <= sdf_stages_4_io_out_imag;
    end
    _T_948_real <= _T_945_real;
    _T_948_imag <= _T_945_imag;
    outputWires_4_real <= _T_948_real;
    outputWires_4_imag <= _T_948_imag;
    if (_GEN_239) begin
      _T_996 <= _T_994;
    end
    if (2'h3 == _GEN_885) begin
      twiddles_5_real <= -16'sh2d41;
    end else if (2'h2 == _GEN_885) begin
      twiddles_5_real <= 16'sh0;
    end else if (2'h1 == _GEN_885) begin
      twiddles_5_real <= 16'sh2d41;
    end else begin
      twiddles_5_real <= 16'sh4000;
    end
    if (2'h3 == _GEN_885) begin
      twiddles_5_imag <= -16'sh2d41;
    end else if (2'h2 == _GEN_885) begin
      twiddles_5_imag <= -16'sh4000;
    end else if (2'h1 == _GEN_885) begin
      twiddles_5_imag <= -16'sh2d41;
    end else begin
      twiddles_5_imag <= 16'sh0;
    end
    _T_1006 <= sdf_stages_5_io_out_real;
    _T_1007 <= twiddles_5_real;
    _T_1008 <= twiddles_5_imag;
    _T_1010 <= $signed(twiddles_5_real) + $signed(twiddles_5_imag);
    _T_1012 <= $signed(sdf_stages_5_io_out_real) + $signed(sdf_stages_5_io_out_imag);
    _T_1014 <= $signed(sdf_stages_5_io_out_imag) - $signed(sdf_stages_5_io_out_real);
    _T_1016 <= $signed(_GEN_957) * $signed(_T_1010);
    _T_1022 <= $signed(_T_1012) * $signed(_GEN_959);
    _T_1028 <= $signed(_T_1014) * $signed(_GEN_961);
    _T_1034 <= $signed(_T_1020) - $signed(_T_1026);
    _T_1036 <= $signed(_T_1020) + $signed(_T_1032);
    _T_1059_real <= sdf_stages_6_io_out_real;
    _T_1059_imag <= sdf_stages_6_io_out_imag;
    _T_1062_real <= _T_1059_real;
    _T_1062_imag <= _T_1059_imag;
    outputWires_6_real <= _T_1062_real;
    outputWires_6_imag <= _T_1062_imag;
    if (reset) begin
      _T_1067 <= 1'h0;
    end else if (_T_51) begin
      _T_1067 <= 1'h0;
    end else if (_T_188) begin
      _T_1067 <= _T_191;
    end else begin
      _T_1067 <= _T_192;
    end
    if (reset) begin
      _T_1068 <= 1'h0;
    end else if (_T_51) begin
      _T_1068 <= 1'h0;
    end else begin
      _T_1068 <= _T_1067;
    end
    if (reset) begin
      _T_1069 <= 1'h0;
    end else if (_T_51) begin
      _T_1069 <= 1'h0;
    end else begin
      _T_1069 <= _T_1068;
    end
    if (reset) begin
      outValid <= 1'h0;
    end else if (_T_51) begin
      outValid <= 1'h0;
    end else begin
      outValid <= _T_1069;
    end
    if (reset) begin
      _T_1071 <= 1'h0;
    end else begin
      _T_1071 <= _T_1070;
    end
    if (reset) begin
      _T_1072 <= 1'h0;
    end else begin
      _T_1072 <= _T_1071;
    end
    if (reset) begin
      _T_1073 <= 1'h0;
    end else begin
      _T_1073 <= _T_1072;
    end
    if (reset) begin
      _T_1074 <= 1'h0;
    end else begin
      _T_1074 <= _T_1073;
    end
  end
endmodule
module SDFFFT_128_16(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [15:0] io_in_bits_real,
  input  [15:0] io_in_bits_imag,
  input         io_out_ready,
  output        io_out_valid,
  output [15:0] io_out_bits_real,
  output [15:0] io_out_bits_imag,
  output        io_lastOut,
  input         io_lastIn,
  input  [6:0]  io_fftSize,
  output        io_busy
);
  wire  SDFChainRadix22_clock; // @[SDFFFT.scala 418:119]
  wire  SDFChainRadix22_reset; // @[SDFFFT.scala 418:119]
  wire  SDFChainRadix22_io_in_ready; // @[SDFFFT.scala 418:119]
  wire  SDFChainRadix22_io_in_valid; // @[SDFFFT.scala 418:119]
  wire [15:0] SDFChainRadix22_io_in_bits_real; // @[SDFFFT.scala 418:119]
  wire [15:0] SDFChainRadix22_io_in_bits_imag; // @[SDFFFT.scala 418:119]
  wire  SDFChainRadix22_io_out_ready; // @[SDFFFT.scala 418:119]
  wire  SDFChainRadix22_io_out_valid; // @[SDFFFT.scala 418:119]
  wire [15:0] SDFChainRadix22_io_out_bits_real; // @[SDFFFT.scala 418:119]
  wire [15:0] SDFChainRadix22_io_out_bits_imag; // @[SDFFFT.scala 418:119]
  wire  SDFChainRadix22_io_lastOut; // @[SDFFFT.scala 418:119]
  wire  SDFChainRadix22_io_lastIn; // @[SDFFFT.scala 418:119]
  wire [6:0] SDFChainRadix22_io_fftSize; // @[SDFFFT.scala 418:119]
  wire  SDFChainRadix22_io_busy; // @[SDFFFT.scala 418:119]
  reg [6:0] cntWin; // @[SDFFFT.scala 265:23]
  reg [31:0] _RAND_0;
  wire [6:0] _T_5 = io_fftSize - 7'h1; // @[SDFFFT.scala 269:41]
  wire [128:0] _T_6 = 129'h2 << _T_5; // @[SDFFFT.scala 269:23]
  wire  _T_7 = io_in_ready & io_in_valid; // @[Decoupled.scala 40:37]
  wire [6:0] _T_9 = cntWin + 7'h1; // @[SDFFFT.scala 274:22]
  wire [6:0] numPoints = _T_6[6:0]; // @[SDFFFT.scala 266:23 SDFFFT.scala 269:15]
  wire [6:0] _T_11 = numPoints - 7'h1; // @[SDFFFT.scala 276:44]
  wire  _T_12 = cntWin == _T_11; // @[SDFFFT.scala 276:29]
  wire  _T_13 = io_lastIn | _T_12; // @[SDFFFT.scala 276:19]
  wire [31:0] _T_84 = $signed(io_in_bits_real) * 16'sh4000; // @[FixedPointTypeClass.scala 42:59]
  wire [31:0] _T_85 = $signed(io_in_bits_imag) * 16'sh4000; // @[FixedPointTypeClass.scala 42:59]
  wire [29:0] _GEN_138 = {$signed(SDFChainRadix22_io_out_bits_imag), 14'h0}; // @[SDFFFT.scala 500:56]
  wire [31:0] _GEN_134 = {{2{_GEN_138[29]}},_GEN_138}; // @[SDFFFT.scala 500:56]
  wire [29:0] _GEN_139 = {$signed(SDFChainRadix22_io_out_bits_real), 14'h0}; // @[SDFFFT.scala 500:56]
  wire [31:0] _GEN_135 = {{2{_GEN_139[29]}},_GEN_139}; // @[SDFFFT.scala 500:56]
  wire [17:0] _GEN_140 = _GEN_135[31:14]; // @[SDFFFT.scala 508:18 SDFFFT.scala 513:28]
  wire [17:0] _GEN_142 = _GEN_134[31:14]; // @[SDFFFT.scala 508:18 SDFFFT.scala 514:28]
  wire [17:0] _GEN_144 = _T_84[31:14]; // @[SDFFFT.scala 503:31 SDFFFT.scala 511:21]
  wire [17:0] _GEN_146 = _T_85[31:14]; // @[SDFFFT.scala 504:31 SDFFFT.scala 511:21]
  SDFChainRadix22 SDFChainRadix22 ( // @[SDFFFT.scala 418:119]
    .clock(SDFChainRadix22_clock),
    .reset(SDFChainRadix22_reset),
    .io_in_ready(SDFChainRadix22_io_in_ready),
    .io_in_valid(SDFChainRadix22_io_in_valid),
    .io_in_bits_real(SDFChainRadix22_io_in_bits_real),
    .io_in_bits_imag(SDFChainRadix22_io_in_bits_imag),
    .io_out_ready(SDFChainRadix22_io_out_ready),
    .io_out_valid(SDFChainRadix22_io_out_valid),
    .io_out_bits_real(SDFChainRadix22_io_out_bits_real),
    .io_out_bits_imag(SDFChainRadix22_io_out_bits_imag),
    .io_lastOut(SDFChainRadix22_io_lastOut),
    .io_lastIn(SDFChainRadix22_io_lastIn),
    .io_fftSize(SDFChainRadix22_io_fftSize),
    .io_busy(SDFChainRadix22_io_busy)
  );
  assign io_in_ready = SDFChainRadix22_io_in_ready; // @[SDFFFT.scala 507:23 SDFFFT.scala 511:21]
  assign io_out_valid = SDFChainRadix22_io_out_valid; // @[SDFFFT.scala 508:18 SDFFFT.scala 516:24]
  assign io_out_bits_real = _GEN_140[15:0]; // @[SDFFFT.scala 508:18 SDFFFT.scala 513:28]
  assign io_out_bits_imag = _GEN_142[15:0]; // @[SDFFFT.scala 508:18 SDFFFT.scala 514:28]
  assign io_lastOut = SDFChainRadix22_io_lastOut; // @[SDFFFT.scala 520:20]
  assign io_busy = SDFChainRadix22_io_busy; // @[SDFFFT.scala 523:15]
  assign SDFChainRadix22_clock = clock;
  assign SDFChainRadix22_reset = reset;
  assign SDFChainRadix22_io_in_valid = io_in_valid; // @[SDFFFT.scala 506:27 SDFFFT.scala 511:21]
  assign SDFChainRadix22_io_in_bits_real = _GEN_144[15:0]; // @[SDFFFT.scala 503:31 SDFFFT.scala 511:21]
  assign SDFChainRadix22_io_in_bits_imag = _GEN_146[15:0]; // @[SDFFFT.scala 504:31 SDFFFT.scala 511:21]
  assign SDFChainRadix22_io_out_ready = io_out_ready; // @[SDFFFT.scala 508:18 SDFFFT.scala 517:28]
  assign SDFChainRadix22_io_lastIn = io_lastIn; // @[SDFFFT.scala 519:23]
  assign SDFChainRadix22_io_fftSize = io_fftSize; // @[SDFFFT.scala 526:28]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cntWin = _RAND_0[6:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      cntWin <= 7'h0;
    end else if (_T_13) begin
      cntWin <= 7'h0;
    end else if (_T_7) begin
      cntWin <= _T_9;
    end
  end
endmodule
module AXI4FFTBlock(
  input         clock,
  input         reset,
  output        auto_mem_in_aw_ready,
  input         auto_mem_in_aw_valid,
  input         auto_mem_in_aw_bits_id,
  input  [29:0] auto_mem_in_aw_bits_addr,
  output        auto_mem_in_w_ready,
  input         auto_mem_in_w_valid,
  input  [31:0] auto_mem_in_w_bits_data,
  input  [3:0]  auto_mem_in_w_bits_strb,
  input         auto_mem_in_b_ready,
  output        auto_mem_in_b_valid,
  output        auto_mem_in_b_bits_id,
  output        auto_mem_in_ar_ready,
  input         auto_mem_in_ar_valid,
  input         auto_mem_in_ar_bits_id,
  input  [29:0] auto_mem_in_ar_bits_addr,
  input  [2:0]  auto_mem_in_ar_bits_size,
  input         auto_mem_in_r_ready,
  output        auto_mem_in_r_valid,
  output        auto_mem_in_r_bits_id,
  output [31:0] auto_mem_in_r_bits_data,
  output        auto_stream_in_ready,
  input         auto_stream_in_valid,
  input  [31:0] auto_stream_in_bits_data,
  input         auto_stream_in_bits_last,
  input         auto_stream_out_ready,
  output        auto_stream_out_valid,
  output [31:0] auto_stream_out_bits_data,
  output        auto_stream_out_bits_last
);
  wire  fft_clock; // @[FFTBlock.scala 53:21]
  wire  fft_reset; // @[FFTBlock.scala 53:21]
  wire  fft_io_in_ready; // @[FFTBlock.scala 53:21]
  wire  fft_io_in_valid; // @[FFTBlock.scala 53:21]
  wire [15:0] fft_io_in_bits_real; // @[FFTBlock.scala 53:21]
  wire [15:0] fft_io_in_bits_imag; // @[FFTBlock.scala 53:21]
  wire  fft_io_out_ready; // @[FFTBlock.scala 53:21]
  wire  fft_io_out_valid; // @[FFTBlock.scala 53:21]
  wire [15:0] fft_io_out_bits_real; // @[FFTBlock.scala 53:21]
  wire [15:0] fft_io_out_bits_imag; // @[FFTBlock.scala 53:21]
  wire  fft_io_lastOut; // @[FFTBlock.scala 53:21]
  wire  fft_io_lastIn; // @[FFTBlock.scala 53:21]
  wire [6:0] fft_io_fftSize; // @[FFTBlock.scala 53:21]
  wire  fft_io_busy; // @[FFTBlock.scala 53:21]
  wire  Queue_clock; // @[Decoupled.scala 296:21]
  wire  Queue_reset; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_bits_read; // @[Decoupled.scala 296:21]
  wire [31:0] Queue_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_bits_extra; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_bits_read; // @[Decoupled.scala 296:21]
  wire [31:0] Queue_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_bits_extra; // @[Decoupled.scala 296:21]
  reg [2:0] fftSize; // @[FFTBlock.scala 59:34]
  reg [31:0] _RAND_0;
  reg  fftDir; // @[FFTBlock.scala 60:34]
  reg [31:0] _RAND_1;
  reg [6:0] keepMSBorLSBReg; // @[FFTBlock.scala 61:34]
  reg [31:0] _RAND_2;
  reg  busy; // @[FFTBlock.scala 64:34]
  reg [31:0] _RAND_3;
  wire  _T_2 = auto_mem_in_aw_valid & auto_mem_in_w_valid; // @[RegisterRouter.scala 40:39]
  wire  _T_3 = auto_mem_in_ar_valid | _T_2; // @[RegisterRouter.scala 40:26]
  wire  _T_4 = ~auto_mem_in_ar_valid; // @[RegisterRouter.scala 42:29]
  wire  _T_47_ready = Queue_io_enq_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 299:17]
  wire [29:0] _T_11 = auto_mem_in_ar_valid ? auto_mem_in_ar_bits_addr : auto_mem_in_aw_bits_addr; // @[RegisterRouter.scala 48:19]
  wire [2:0] _T_226 = {_T_11[4],_T_11[3],_T_11[2]}; // @[Cat.scala 29:58]
  wire [5:0] _T_51 = _T_11[7:2] & 6'h38; // @[RegisterRouter.scala 59:16]
  wire  _T_61 = _T_51 == 6'h0; // @[RegisterRouter.scala 59:16]
  wire  _T_5 = _T_47_ready & _T_4; // @[RegisterRouter.scala 42:26]
  wire [1:0] _T_14 = 2'h1 << auto_mem_in_ar_bits_size[0]; // @[OneHot.scala 65:12]
  wire [1:0] _T_16 = _T_14 | 2'h1; // @[Misc.scala 200:81]
  wire  _T_17 = auto_mem_in_ar_bits_size >= 3'h2; // @[Misc.scala 204:21]
  wire  _T_20 = ~auto_mem_in_ar_bits_addr[1]; // @[Misc.scala 209:20]
  wire  _T_22 = _T_16[1] & _T_20; // @[Misc.scala 213:38]
  wire  _T_23 = _T_17 | _T_22; // @[Misc.scala 213:29]
  wire  _T_25 = _T_16[1] & auto_mem_in_ar_bits_addr[1]; // @[Misc.scala 213:38]
  wire  _T_26 = _T_17 | _T_25; // @[Misc.scala 213:29]
  wire  _T_29 = ~auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 209:20]
  wire  _T_30 = _T_20 & _T_29; // @[Misc.scala 212:27]
  wire  _T_31 = _T_16[0] & _T_30; // @[Misc.scala 213:38]
  wire  _T_32 = _T_23 | _T_31; // @[Misc.scala 213:29]
  wire  _T_33 = _T_20 & auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  wire  _T_34 = _T_16[0] & _T_33; // @[Misc.scala 213:38]
  wire  _T_35 = _T_23 | _T_34; // @[Misc.scala 213:29]
  wire  _T_36 = auto_mem_in_ar_bits_addr[1] & _T_29; // @[Misc.scala 212:27]
  wire  _T_37 = _T_16[0] & _T_36; // @[Misc.scala 213:38]
  wire  _T_38 = _T_26 | _T_37; // @[Misc.scala 213:29]
  wire  _T_39 = auto_mem_in_ar_bits_addr[1] & auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  wire  _T_40 = _T_16[0] & _T_39; // @[Misc.scala 213:38]
  wire  _T_41 = _T_26 | _T_40; // @[Misc.scala 213:29]
  wire [3:0] _T_44 = {_T_41,_T_38,_T_35,_T_32}; // @[Cat.scala 29:58]
  wire [3:0] _T_46 = auto_mem_in_ar_valid ? _T_44 : auto_mem_in_w_bits_strb; // @[RegisterRouter.scala 54:25]
  wire [7:0] _T_71 = _T_46[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_73 = _T_46[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_75 = _T_46[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_77 = _T_46[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_80 = {_T_77,_T_75,_T_73,_T_71}; // @[Cat.scala 29:58]
  wire  _T_99 = _T_80[2:0] == 3'h7; // @[RegisterRouter.scala 59:16]
  wire  _T_245 = _T_3 & _T_47_ready; // @[RegisterRouter.scala 59:16]
  wire [7:0] _T_227 = 8'h1 << _T_226; // @[OneHot.scala 58:35]
  wire  _T_292 = _T_245 & _T_4; // @[RegisterRouter.scala 59:16]
  wire  _T_294 = _T_292 & _T_227[0]; // @[RegisterRouter.scala 59:16]
  wire  _T_295 = _T_294 & _T_61; // @[RegisterRouter.scala 59:16]
  wire  _T_106 = _T_295 & _T_99; // @[RegisterRouter.scala 59:16]
  wire  _T_299 = _T_292 & _T_227[1]; // @[RegisterRouter.scala 59:16]
  wire  _T_300 = _T_299 & _T_61; // @[RegisterRouter.scala 59:16]
  wire  _T_129 = _T_300 & _T_80[0]; // @[RegisterRouter.scala 59:16]
  wire  _GEN_1 = _T_129 ? auto_mem_in_w_bits_data[0] : fftDir; // @[RegField.scala 134:88]
  wire  _T_145 = _T_80[6:0] == 7'h7f; // @[RegisterRouter.scala 59:16]
  wire  _T_304 = _T_292 & _T_227[2]; // @[RegisterRouter.scala 59:16]
  wire  _T_305 = _T_304 & _T_61; // @[RegisterRouter.scala 59:16]
  wire  _T_152 = _T_305 & _T_145; // @[RegisterRouter.scala 59:16]
  wire  _GEN_36 = 3'h1 == _T_226 ? _T_61 : _T_61; // @[MuxLiteral.scala 48:10]
  wire  _GEN_37 = 3'h2 == _T_226 ? _T_61 : _GEN_36; // @[MuxLiteral.scala 48:10]
  wire  _GEN_38 = 3'h3 == _T_226 ? _T_61 : _GEN_37; // @[MuxLiteral.scala 48:10]
  wire  _GEN_39 = 3'h4 == _T_226 ? _T_61 : _GEN_38; // @[MuxLiteral.scala 48:10]
  wire  _GEN_51 = 3'h5 == _T_226; // @[MuxLiteral.scala 48:10]
  wire  _GEN_40 = _GEN_51 | _GEN_39; // @[MuxLiteral.scala 48:10]
  wire  _GEN_52 = 3'h6 == _T_226; // @[MuxLiteral.scala 48:10]
  wire  _GEN_41 = _GEN_52 | _GEN_40; // @[MuxLiteral.scala 48:10]
  wire  _GEN_53 = 3'h7 == _T_226; // @[MuxLiteral.scala 48:10]
  wire  _GEN_42 = _GEN_53 | _GEN_41; // @[MuxLiteral.scala 48:10]
  wire [6:0] _T_437_0 = {{4'd0}, fftSize}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [6:0] _T_437_1 = {{6'd0}, fftDir}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [6:0] _GEN_44 = 3'h1 == _T_226 ? _T_437_1 : _T_437_0; // @[MuxLiteral.scala 48:10]
  wire [6:0] _GEN_45 = 3'h2 == _T_226 ? keepMSBorLSBReg : _GEN_44; // @[MuxLiteral.scala 48:10]
  wire [6:0] _T_437_3 = {{6'd0}, busy}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [6:0] _GEN_46 = 3'h3 == _T_226 ? _T_437_3 : _GEN_45; // @[MuxLiteral.scala 48:10]
  wire [6:0] _GEN_47 = 3'h4 == _T_226 ? 7'h0 : _GEN_46; // @[MuxLiteral.scala 48:10]
  wire [6:0] _GEN_48 = 3'h5 == _T_226 ? 7'h0 : _GEN_47; // @[MuxLiteral.scala 48:10]
  wire [6:0] _GEN_49 = 3'h6 == _T_226 ? 7'h0 : _GEN_48; // @[MuxLiteral.scala 48:10]
  wire [6:0] _GEN_50 = 3'h7 == _T_226 ? 7'h0 : _GEN_49; // @[MuxLiteral.scala 48:10]
  wire [6:0] _T_439 = _GEN_42 ? _GEN_50 : 7'h0; // @[RegisterRouter.scala 59:16]
  wire  _T_440_bits_read = Queue_io_deq_bits_read; // @[Decoupled.scala 317:19 Decoupled.scala 318:14]
  wire  _T_440_valid = Queue_io_deq_valid; // @[Decoupled.scala 317:19 Decoupled.scala 319:15]
  wire  _T_443 = ~_T_440_bits_read; // @[RegisterRouter.scala 65:29]
  SDFFFT_128_16 fft ( // @[FFTBlock.scala 53:21]
    .clock(fft_clock),
    .reset(fft_reset),
    .io_in_ready(fft_io_in_ready),
    .io_in_valid(fft_io_in_valid),
    .io_in_bits_real(fft_io_in_bits_real),
    .io_in_bits_imag(fft_io_in_bits_imag),
    .io_out_ready(fft_io_out_ready),
    .io_out_valid(fft_io_out_valid),
    .io_out_bits_real(fft_io_out_bits_real),
    .io_out_bits_imag(fft_io_out_bits_imag),
    .io_lastOut(fft_io_lastOut),
    .io_lastIn(fft_io_lastIn),
    .io_fftSize(fft_io_fftSize),
    .io_busy(fft_io_busy)
  );
  Queue Queue ( // @[Decoupled.scala 296:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_read(Queue_io_enq_bits_read),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_extra(Queue_io_enq_bits_extra),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_read(Queue_io_deq_bits_read),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_extra(Queue_io_deq_bits_extra)
  );
  assign auto_mem_in_aw_ready = _T_5 & auto_mem_in_w_valid; // @[LazyModule.scala 173:31]
  assign auto_mem_in_w_ready = _T_5 & auto_mem_in_aw_valid; // @[LazyModule.scala 173:31]
  assign auto_mem_in_b_valid = _T_440_valid & _T_443; // @[LazyModule.scala 173:31]
  assign auto_mem_in_b_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_mem_in_ar_ready = Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_valid = _T_440_valid & _T_440_bits_read; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 173:31]
  assign auto_stream_in_ready = fft_io_in_ready; // @[LazyModule.scala 173:31]
  assign auto_stream_out_valid = fft_io_out_valid; // @[LazyModule.scala 173:49]
  assign auto_stream_out_bits_data = {fft_io_out_bits_real,fft_io_out_bits_imag}; // @[LazyModule.scala 173:49]
  assign auto_stream_out_bits_last = fft_io_lastOut; // @[LazyModule.scala 173:49]
  assign fft_clock = clock;
  assign fft_reset = reset;
  assign fft_io_in_valid = auto_stream_in_valid; // @[FFTBlock.scala 103:24]
  assign fft_io_in_bits_real = auto_stream_in_bits_data[31:16]; // @[FFTBlock.scala 104:24]
  assign fft_io_in_bits_imag = auto_stream_in_bits_data[15:0]; // @[FFTBlock.scala 104:24]
  assign fft_io_out_ready = auto_stream_out_ready; // @[FFTBlock.scala 111:22]
  assign fft_io_lastIn = auto_stream_in_bits_last; // @[FFTBlock.scala 106:24]
  assign fft_io_fftSize = {{4'd0}, fftSize}; // @[FFTBlock.scala 71:26]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_mem_in_ar_valid | _T_2; // @[Decoupled.scala 297:22]
  assign Queue_io_enq_bits_read = auto_mem_in_ar_valid; // @[Decoupled.scala 298:21]
  assign Queue_io_enq_bits_data = {{25'd0}, _T_439}; // @[Decoupled.scala 298:21]
  assign Queue_io_enq_bits_extra = auto_mem_in_ar_valid ? auto_mem_in_ar_bits_id : auto_mem_in_aw_bits_id; // @[Decoupled.scala 298:21]
  assign Queue_io_deq_ready = _T_440_bits_read ? auto_mem_in_r_ready : auto_mem_in_b_ready; // @[Decoupled.scala 320:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  fftSize = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  fftDir = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  keepMSBorLSBReg = _RAND_2[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  busy = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      fftSize <= 3'h7;
    end else if (_T_106) begin
      fftSize <= auto_mem_in_w_bits_data[2:0];
    end
    fftDir <= reset | _GEN_1;
    if (reset) begin
      keepMSBorLSBReg <= 7'h0;
    end else if (_T_152) begin
      keepMSBorLSBReg <= auto_mem_in_w_bits_data[6:0];
    end
    if (reset) begin
      busy <= 1'h0;
    end else begin
      busy <= fft_io_busy;
    end
  end
endmodule
module AXI4Splitter_3(
  input         clock,
  input         reset,
  output        auto_mem_in_aw_ready,
  input         auto_mem_in_aw_valid,
  input         auto_mem_in_aw_bits_id,
  input  [29:0] auto_mem_in_aw_bits_addr,
  output        auto_mem_in_w_ready,
  input         auto_mem_in_w_valid,
  input  [31:0] auto_mem_in_w_bits_data,
  input  [3:0]  auto_mem_in_w_bits_strb,
  input         auto_mem_in_b_ready,
  output        auto_mem_in_b_valid,
  output        auto_mem_in_b_bits_id,
  output        auto_mem_in_ar_ready,
  input         auto_mem_in_ar_valid,
  input         auto_mem_in_ar_bits_id,
  input  [29:0] auto_mem_in_ar_bits_addr,
  input  [2:0]  auto_mem_in_ar_bits_size,
  input         auto_mem_in_r_ready,
  output        auto_mem_in_r_valid,
  output        auto_mem_in_r_bits_id,
  output [31:0] auto_mem_in_r_bits_data,
  output        auto_stream_in_ready,
  input         auto_stream_in_valid,
  input  [31:0] auto_stream_in_bits_data,
  input         auto_stream_in_bits_last,
  input         auto_stream_out_1_ready,
  output        auto_stream_out_1_valid,
  output [31:0] auto_stream_out_1_bits_data,
  output        auto_stream_out_1_bits_last,
  input         auto_stream_out_0_ready,
  output        auto_stream_out_0_valid,
  output [31:0] auto_stream_out_0_bits_data,
  output        auto_stream_out_0_bits_last
);
  wire  Queue_clock; // @[Decoupled.scala 296:21]
  wire  Queue_reset; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_bits_read; // @[Decoupled.scala 296:21]
  wire [31:0] Queue_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_bits_extra; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_bits_read; // @[Decoupled.scala 296:21]
  wire [31:0] Queue_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_bits_extra; // @[Decoupled.scala 296:21]
  reg [31:0] ctrlReg; // @[Splitter.scala 27:26]
  reg [31:0] _RAND_0;
  reg [31:0] maskReg; // @[Splitter.scala 28:26]
  reg [31:0] _RAND_1;
  wire  _T_4 = auto_mem_in_aw_valid & auto_mem_in_w_valid; // @[RegisterRouter.scala 40:39]
  wire  _T_5 = auto_mem_in_ar_valid | _T_4; // @[RegisterRouter.scala 40:26]
  wire  _T_6 = ~auto_mem_in_ar_valid; // @[RegisterRouter.scala 42:29]
  wire  _T_49_ready = Queue_io_enq_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 299:17]
  wire [29:0] _T_13 = auto_mem_in_ar_valid ? auto_mem_in_ar_bits_addr : auto_mem_in_aw_bits_addr; // @[RegisterRouter.scala 48:19]
  wire [1:0] _T_53 = _T_13[3:2] & 2'h2; // @[RegisterRouter.scala 59:16]
  wire  _T_55 = _T_53 == 2'h0; // @[RegisterRouter.scala 59:16]
  wire  _T_7 = _T_49_ready & _T_6; // @[RegisterRouter.scala 42:26]
  wire [1:0] _T_16 = 2'h1 << auto_mem_in_ar_bits_size[0]; // @[OneHot.scala 65:12]
  wire [1:0] _T_18 = _T_16 | 2'h1; // @[Misc.scala 200:81]
  wire  _T_19 = auto_mem_in_ar_bits_size >= 3'h2; // @[Misc.scala 204:21]
  wire  _T_22 = ~auto_mem_in_ar_bits_addr[1]; // @[Misc.scala 209:20]
  wire  _T_24 = _T_18[1] & _T_22; // @[Misc.scala 213:38]
  wire  _T_25 = _T_19 | _T_24; // @[Misc.scala 213:29]
  wire  _T_27 = _T_18[1] & auto_mem_in_ar_bits_addr[1]; // @[Misc.scala 213:38]
  wire  _T_28 = _T_19 | _T_27; // @[Misc.scala 213:29]
  wire  _T_31 = ~auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 209:20]
  wire  _T_32 = _T_22 & _T_31; // @[Misc.scala 212:27]
  wire  _T_33 = _T_18[0] & _T_32; // @[Misc.scala 213:38]
  wire  _T_34 = _T_25 | _T_33; // @[Misc.scala 213:29]
  wire  _T_35 = _T_22 & auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  wire  _T_36 = _T_18[0] & _T_35; // @[Misc.scala 213:38]
  wire  _T_37 = _T_25 | _T_36; // @[Misc.scala 213:29]
  wire  _T_38 = auto_mem_in_ar_bits_addr[1] & _T_31; // @[Misc.scala 212:27]
  wire  _T_39 = _T_18[0] & _T_38; // @[Misc.scala 213:38]
  wire  _T_40 = _T_28 | _T_39; // @[Misc.scala 213:29]
  wire  _T_41 = auto_mem_in_ar_bits_addr[1] & auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  wire  _T_42 = _T_18[0] & _T_41; // @[Misc.scala 213:38]
  wire  _T_43 = _T_28 | _T_42; // @[Misc.scala 213:29]
  wire [3:0] _T_46 = {_T_43,_T_40,_T_37,_T_34}; // @[Cat.scala 29:58]
  wire [3:0] _T_48 = auto_mem_in_ar_valid ? _T_46 : auto_mem_in_w_bits_strb; // @[RegisterRouter.scala 54:25]
  wire [7:0] _T_67 = _T_48[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_69 = _T_48[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_71 = _T_48[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_73 = _T_48[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_76 = {_T_73,_T_71,_T_69,_T_67}; // @[Cat.scala 29:58]
  wire  _T_95 = _T_76 == 32'hffffffff; // @[RegisterRouter.scala 59:16]
  wire  _T_148 = _T_5 & _T_49_ready; // @[RegisterRouter.scala 59:16]
  wire [1:0] _T_142 = 2'h1 << _T_13[2]; // @[OneHot.scala 58:35]
  wire  _T_165 = _T_148 & _T_6; // @[RegisterRouter.scala 59:16]
  wire  _T_172 = _T_165 & _T_142[1]; // @[RegisterRouter.scala 59:16]
  wire  _T_173 = _T_172 & _T_55; // @[RegisterRouter.scala 59:16]
  wire  _T_102 = _T_173 & _T_95; // @[RegisterRouter.scala 59:16]
  wire  _T_167 = _T_165 & _T_142[0]; // @[RegisterRouter.scala 59:16]
  wire  _T_168 = _T_167 & _T_55; // @[RegisterRouter.scala 59:16]
  wire  _T_125 = _T_168 & _T_95; // @[RegisterRouter.scala 59:16]
  wire  _GEN_11 = _T_13[2] ? _T_55 : _T_55; // @[MuxLiteral.scala 48:10]
  wire [31:0] _GEN_13 = _T_13[2] ? maskReg : ctrlReg; // @[MuxLiteral.scala 48:10]
  wire  _T_223_bits_read = Queue_io_deq_bits_read; // @[Decoupled.scala 317:19 Decoupled.scala 318:14]
  wire  _T_223_valid = Queue_io_deq_valid; // @[Decoupled.scala 317:19 Decoupled.scala 319:15]
  wire  _T_226 = ~_T_223_bits_read; // @[RegisterRouter.scala 65:29]
  wire  readyOR = auto_stream_out_0_ready | auto_stream_out_1_ready; // @[Splitter.scala 45:34]
  wire  readyAND = auto_stream_out_0_ready & auto_stream_out_1_ready; // @[Splitter.scala 46:34]
  wire  _T_229 = ctrlReg == 32'h0; // @[Splitter.scala 49:19]
  wire  _T_230 = ctrlReg == 32'h1; // @[Splitter.scala 52:24]
  wire  _GEN_14 = _T_230 & readyOR; // @[Splitter.scala 52:33]
  wire  _T_233 = ~maskReg[0]; // @[Splitter.scala 62:34]
  wire  _T_237 = ~maskReg[1]; // @[Splitter.scala 62:34]
  Queue Queue ( // @[Decoupled.scala 296:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_read(Queue_io_enq_bits_read),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_extra(Queue_io_enq_bits_extra),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_read(Queue_io_deq_bits_read),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_extra(Queue_io_deq_bits_extra)
  );
  assign auto_mem_in_aw_ready = _T_7 & auto_mem_in_w_valid; // @[LazyModule.scala 173:31]
  assign auto_mem_in_w_ready = _T_7 & auto_mem_in_aw_valid; // @[LazyModule.scala 173:31]
  assign auto_mem_in_b_valid = _T_223_valid & _T_226; // @[LazyModule.scala 173:31]
  assign auto_mem_in_b_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_mem_in_ar_ready = Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_valid = _T_223_valid & _T_223_bits_read; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 173:31]
  assign auto_stream_in_ready = _T_229 ? readyAND : _GEN_14; // @[LazyModule.scala 173:31]
  assign auto_stream_out_1_valid = auto_stream_in_valid & _T_237; // @[LazyModule.scala 173:49]
  assign auto_stream_out_1_bits_data = auto_stream_in_bits_data; // @[LazyModule.scala 173:49]
  assign auto_stream_out_1_bits_last = auto_stream_in_bits_last; // @[LazyModule.scala 173:49]
  assign auto_stream_out_0_valid = auto_stream_in_valid & _T_233; // @[LazyModule.scala 173:49]
  assign auto_stream_out_0_bits_data = auto_stream_in_bits_data; // @[LazyModule.scala 173:49]
  assign auto_stream_out_0_bits_last = auto_stream_in_bits_last; // @[LazyModule.scala 173:49]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_mem_in_ar_valid | _T_4; // @[Decoupled.scala 297:22]
  assign Queue_io_enq_bits_read = auto_mem_in_ar_valid; // @[Decoupled.scala 298:21]
  assign Queue_io_enq_bits_data = _GEN_11 ? _GEN_13 : 32'h0; // @[Decoupled.scala 298:21]
  assign Queue_io_enq_bits_extra = auto_mem_in_ar_valid ? auto_mem_in_ar_bits_id : auto_mem_in_aw_bits_id; // @[Decoupled.scala 298:21]
  assign Queue_io_deq_ready = _T_223_bits_read ? auto_mem_in_r_ready : auto_mem_in_b_ready; // @[Decoupled.scala 320:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ctrlReg = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  maskReg = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      ctrlReg <= 32'h0;
    end else if (_T_125) begin
      ctrlReg <= auto_mem_in_w_bits_data;
    end
    if (reset) begin
      maskReg <= 32'h0;
    end else if (_T_102) begin
      maskReg <= auto_mem_in_w_bits_data;
    end
  end
endmodule
module AXI4StreamMux_4(
  input         clock,
  input         reset,
  output        auto_register_in_aw_ready,
  input         auto_register_in_aw_valid,
  input         auto_register_in_aw_bits_id,
  input  [29:0] auto_register_in_aw_bits_addr,
  output        auto_register_in_w_ready,
  input         auto_register_in_w_valid,
  input  [31:0] auto_register_in_w_bits_data,
  input  [3:0]  auto_register_in_w_bits_strb,
  input         auto_register_in_b_ready,
  output        auto_register_in_b_valid,
  output        auto_register_in_b_bits_id,
  output        auto_register_in_ar_ready,
  input         auto_register_in_ar_valid,
  input         auto_register_in_ar_bits_id,
  input  [29:0] auto_register_in_ar_bits_addr,
  input  [2:0]  auto_register_in_ar_bits_size,
  input         auto_register_in_r_ready,
  output        auto_register_in_r_valid,
  output        auto_register_in_r_bits_id,
  output [31:0] auto_register_in_r_bits_data,
  output        auto_stream_in_2_ready,
  input         auto_stream_in_2_valid,
  input  [31:0] auto_stream_in_2_bits_data,
  input         auto_stream_in_2_bits_last,
  output        auto_stream_in_1_ready,
  input         auto_stream_in_1_valid,
  input  [31:0] auto_stream_in_1_bits_data,
  input         auto_stream_in_1_bits_last,
  output        auto_stream_in_0_ready,
  input         auto_stream_in_0_valid,
  input  [31:0] auto_stream_in_0_bits_data,
  input         auto_stream_in_0_bits_last,
  input         auto_stream_out_0_ready,
  output        auto_stream_out_0_valid,
  output [31:0] auto_stream_out_0_bits_data,
  output        auto_stream_out_0_bits_last
);
  wire  Queue_clock; // @[Decoupled.scala 296:21]
  wire  Queue_reset; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_bits_read; // @[Decoupled.scala 296:21]
  wire [31:0] Queue_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_bits_extra; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_bits_read; // @[Decoupled.scala 296:21]
  wire [31:0] Queue_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_bits_extra; // @[Decoupled.scala 296:21]
  reg [2:0] sels_0; // @[Mux.scala 32:23]
  reg [31:0] _RAND_0;
  reg [2:0] sels_1; // @[Mux.scala 32:23]
  reg [31:0] _RAND_1;
  wire  _T_3 = sels_0 == 3'h0; // @[Mux.scala 45:28]
  wire  _GEN_7 = _T_3 & auto_stream_in_0_valid; // @[Mux.scala 45:41]
  wire  _GEN_8 = _T_3 & auto_stream_out_0_ready; // @[Mux.scala 45:41]
  wire  _T_4 = sels_0 == 3'h1; // @[Mux.scala 45:28]
  wire  _GEN_12 = _T_4 ? auto_stream_in_1_bits_last : auto_stream_in_0_bits_last; // @[Mux.scala 45:41]
  wire [31:0] _GEN_15 = _T_4 ? auto_stream_in_1_bits_data : auto_stream_in_0_bits_data; // @[Mux.scala 45:41]
  wire  _GEN_16 = _T_4 ? auto_stream_in_1_valid : _GEN_7; // @[Mux.scala 45:41]
  wire  _GEN_17 = _T_4 & auto_stream_out_0_ready; // @[Mux.scala 45:41]
  wire  _T_5 = sels_0 == 3'h2; // @[Mux.scala 45:28]
  wire  _GEN_21 = _T_5 ? auto_stream_in_2_bits_last : _GEN_12; // @[Mux.scala 45:41]
  wire [31:0] _GEN_24 = _T_5 ? auto_stream_in_2_bits_data : _GEN_15; // @[Mux.scala 45:41]
  wire  _GEN_25 = _T_5 ? auto_stream_in_2_valid : _GEN_16; // @[Mux.scala 45:41]
  wire  _GEN_26 = _T_5 & auto_stream_out_0_ready; // @[Mux.scala 45:41]
  wire  _T_6 = sels_0 == 3'h3; // @[Mux.scala 45:28]
  wire  _GEN_30 = _T_6 ? 1'h0 : _GEN_21; // @[Mux.scala 45:41]
  wire [31:0] _GEN_33 = _T_6 ? 32'hffffffff : _GEN_24; // @[Mux.scala 45:41]
  wire  _GEN_34 = _T_6 | _GEN_25; // @[Mux.scala 45:41]
  wire  _T_7 = sels_0 == 3'h4; // @[Mux.scala 45:28]
  wire  _T_8 = sels_0 == sels_1; // @[Mux.scala 40:46]
  wire [2:0] _T_10 = _T_8 ? 3'h5 : sels_1; // @[Mux.scala 41:29]
  wire  _T_11 = _T_10 == 3'h0; // @[Mux.scala 45:28]
  wire  _T_12 = _T_10 == 3'h1; // @[Mux.scala 45:28]
  wire  _T_13 = _T_10 == 3'h2; // @[Mux.scala 45:28]
  wire  _T_17 = auto_register_in_aw_valid & auto_register_in_w_valid; // @[RegisterRouter.scala 40:39]
  wire  _T_18 = auto_register_in_ar_valid | _T_17; // @[RegisterRouter.scala 40:26]
  wire  _T_19 = ~auto_register_in_ar_valid; // @[RegisterRouter.scala 42:29]
  wire  _T_62_ready = Queue_io_enq_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 299:17]
  wire [29:0] _T_26 = auto_register_in_ar_valid ? auto_register_in_ar_bits_addr : auto_register_in_aw_bits_addr; // @[RegisterRouter.scala 48:19]
  wire [1:0] _T_66 = _T_26[3:2] & 2'h2; // @[RegisterRouter.scala 59:16]
  wire  _T_68 = _T_66 == 2'h0; // @[RegisterRouter.scala 59:16]
  wire  _T_20 = _T_62_ready & _T_19; // @[RegisterRouter.scala 42:26]
  wire [1:0] _T_29 = 2'h1 << auto_register_in_ar_bits_size[0]; // @[OneHot.scala 65:12]
  wire [1:0] _T_31 = _T_29 | 2'h1; // @[Misc.scala 200:81]
  wire  _T_32 = auto_register_in_ar_bits_size >= 3'h2; // @[Misc.scala 204:21]
  wire  _T_35 = ~auto_register_in_ar_bits_addr[1]; // @[Misc.scala 209:20]
  wire  _T_37 = _T_31[1] & _T_35; // @[Misc.scala 213:38]
  wire  _T_38 = _T_32 | _T_37; // @[Misc.scala 213:29]
  wire  _T_40 = _T_31[1] & auto_register_in_ar_bits_addr[1]; // @[Misc.scala 213:38]
  wire  _T_41 = _T_32 | _T_40; // @[Misc.scala 213:29]
  wire  _T_44 = ~auto_register_in_ar_bits_addr[0]; // @[Misc.scala 209:20]
  wire  _T_45 = _T_35 & _T_44; // @[Misc.scala 212:27]
  wire  _T_46 = _T_31[0] & _T_45; // @[Misc.scala 213:38]
  wire  _T_47 = _T_38 | _T_46; // @[Misc.scala 213:29]
  wire  _T_48 = _T_35 & auto_register_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  wire  _T_49 = _T_31[0] & _T_48; // @[Misc.scala 213:38]
  wire  _T_50 = _T_38 | _T_49; // @[Misc.scala 213:29]
  wire  _T_51 = auto_register_in_ar_bits_addr[1] & _T_44; // @[Misc.scala 212:27]
  wire  _T_52 = _T_31[0] & _T_51; // @[Misc.scala 213:38]
  wire  _T_53 = _T_41 | _T_52; // @[Misc.scala 213:29]
  wire  _T_54 = auto_register_in_ar_bits_addr[1] & auto_register_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  wire  _T_55 = _T_31[0] & _T_54; // @[Misc.scala 213:38]
  wire  _T_56 = _T_41 | _T_55; // @[Misc.scala 213:29]
  wire [3:0] _T_59 = {_T_56,_T_53,_T_50,_T_47}; // @[Cat.scala 29:58]
  wire [3:0] _T_61 = auto_register_in_ar_valid ? _T_59 : auto_register_in_w_bits_strb; // @[RegisterRouter.scala 54:25]
  wire [7:0] _T_80 = _T_61[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_82 = _T_61[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_84 = _T_61[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_86 = _T_61[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_89 = {_T_86,_T_84,_T_82,_T_80}; // @[Cat.scala 29:58]
  wire  _T_108 = _T_89[2:0] == 3'h7; // @[RegisterRouter.scala 59:16]
  wire  _T_161 = _T_18 & _T_62_ready; // @[RegisterRouter.scala 59:16]
  wire [1:0] _T_155 = 2'h1 << _T_26[2]; // @[OneHot.scala 58:35]
  wire  _T_178 = _T_161 & _T_19; // @[RegisterRouter.scala 59:16]
  wire  _T_185 = _T_178 & _T_155[1]; // @[RegisterRouter.scala 59:16]
  wire  _T_186 = _T_185 & _T_68; // @[RegisterRouter.scala 59:16]
  wire  _T_115 = _T_186 & _T_108; // @[RegisterRouter.scala 59:16]
  wire  _T_180 = _T_178 & _T_155[0]; // @[RegisterRouter.scala 59:16]
  wire  _T_181 = _T_180 & _T_68; // @[RegisterRouter.scala 59:16]
  wire  _T_138 = _T_181 & _T_108; // @[RegisterRouter.scala 59:16]
  wire  _GEN_101 = _T_26[2] ? _T_68 : _T_68; // @[MuxLiteral.scala 48:10]
  wire [2:0] _GEN_103 = _T_26[2] ? sels_1 : sels_0; // @[MuxLiteral.scala 48:10]
  wire [2:0] _T_235 = _GEN_101 ? _GEN_103 : 3'h0; // @[RegisterRouter.scala 59:16]
  wire  _T_236_bits_read = Queue_io_deq_bits_read; // @[Decoupled.scala 317:19 Decoupled.scala 318:14]
  wire  _T_236_valid = Queue_io_deq_valid; // @[Decoupled.scala 317:19 Decoupled.scala 319:15]
  wire  _T_239 = ~_T_236_bits_read; // @[RegisterRouter.scala 65:29]
  Queue Queue ( // @[Decoupled.scala 296:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_read(Queue_io_enq_bits_read),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_extra(Queue_io_enq_bits_extra),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_read(Queue_io_deq_bits_read),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_extra(Queue_io_deq_bits_extra)
  );
  assign auto_register_in_aw_ready = _T_20 & auto_register_in_w_valid; // @[LazyModule.scala 173:31]
  assign auto_register_in_w_ready = _T_20 & auto_register_in_aw_valid; // @[LazyModule.scala 173:31]
  assign auto_register_in_b_valid = _T_236_valid & _T_239; // @[LazyModule.scala 173:31]
  assign auto_register_in_b_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_register_in_ar_ready = Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_register_in_r_valid = _T_236_valid & _T_236_bits_read; // @[LazyModule.scala 173:31]
  assign auto_register_in_r_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_register_in_r_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 173:31]
  assign auto_stream_in_2_ready = _T_13 | _GEN_26; // @[LazyModule.scala 173:31]
  assign auto_stream_in_1_ready = _T_12 | _GEN_17; // @[LazyModule.scala 173:31]
  assign auto_stream_in_0_ready = _T_11 | _GEN_8; // @[LazyModule.scala 173:31]
  assign auto_stream_out_0_valid = _T_7 | _GEN_34; // @[LazyModule.scala 173:49]
  assign auto_stream_out_0_bits_data = _T_7 ? 32'h0 : _GEN_33; // @[LazyModule.scala 173:49]
  assign auto_stream_out_0_bits_last = _T_7 ? 1'h0 : _GEN_30; // @[LazyModule.scala 173:49]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_register_in_ar_valid | _T_17; // @[Decoupled.scala 297:22]
  assign Queue_io_enq_bits_read = auto_register_in_ar_valid; // @[Decoupled.scala 298:21]
  assign Queue_io_enq_bits_data = {{29'd0}, _T_235}; // @[Decoupled.scala 298:21]
  assign Queue_io_enq_bits_extra = auto_register_in_ar_valid ? auto_register_in_ar_bits_id : auto_register_in_aw_bits_id; // @[Decoupled.scala 298:21]
  assign Queue_io_deq_ready = _T_236_bits_read ? auto_register_in_r_ready : auto_register_in_b_ready; // @[Decoupled.scala 320:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  sels_0 = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  sels_1 = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      sels_0 <= 3'h5;
    end else if (_T_138) begin
      sels_0 <= auto_register_in_w_bits_data[2:0];
    end
    if (reset) begin
      sels_1 <= 3'h5;
    end else if (_T_115) begin
      sels_1 <= auto_register_in_w_bits_data[2:0];
    end
  end
endmodule
module AXI4StreamMux_5(
  input         clock,
  input         reset,
  output        auto_register_in_aw_ready,
  input         auto_register_in_aw_valid,
  input         auto_register_in_aw_bits_id,
  input  [29:0] auto_register_in_aw_bits_addr,
  output        auto_register_in_w_ready,
  input         auto_register_in_w_valid,
  input  [31:0] auto_register_in_w_bits_data,
  input  [3:0]  auto_register_in_w_bits_strb,
  input         auto_register_in_b_ready,
  output        auto_register_in_b_valid,
  output        auto_register_in_b_bits_id,
  output        auto_register_in_ar_ready,
  input         auto_register_in_ar_valid,
  input         auto_register_in_ar_bits_id,
  input  [29:0] auto_register_in_ar_bits_addr,
  input  [2:0]  auto_register_in_ar_bits_size,
  input         auto_register_in_r_ready,
  output        auto_register_in_r_valid,
  output        auto_register_in_r_bits_id,
  output [31:0] auto_register_in_r_bits_data,
  output        auto_stream_in_ready,
  input         auto_stream_in_valid,
  input  [31:0] auto_stream_in_bits_data,
  input         auto_stream_in_bits_last,
  input         auto_stream_out_1_ready,
  output        auto_stream_out_1_valid,
  output [31:0] auto_stream_out_1_bits_data,
  output        auto_stream_out_1_bits_last
);
  wire  Queue_clock; // @[Decoupled.scala 296:21]
  wire  Queue_reset; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_bits_read; // @[Decoupled.scala 296:21]
  wire [31:0] Queue_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_bits_extra; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_bits_read; // @[Decoupled.scala 296:21]
  wire [31:0] Queue_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_bits_extra; // @[Decoupled.scala 296:21]
  reg  sels_0; // @[Mux.scala 32:23]
  reg [31:0] _RAND_0;
  reg  sels_1; // @[Mux.scala 32:23]
  reg [31:0] _RAND_1;
  wire  _T_3 = ~sels_0; // @[Mux.scala 45:28]
  wire  _T_4 = sels_0 == sels_1; // @[Mux.scala 40:46]
  wire  _T_6 = _T_4 | sels_1; // @[Mux.scala 41:29]
  wire  _T_7 = ~_T_6; // @[Mux.scala 45:28]
  wire  _T_9 = auto_register_in_aw_valid & auto_register_in_w_valid; // @[RegisterRouter.scala 40:39]
  wire  _T_10 = auto_register_in_ar_valid | _T_9; // @[RegisterRouter.scala 40:26]
  wire  _T_11 = ~auto_register_in_ar_valid; // @[RegisterRouter.scala 42:29]
  wire  _T_54_ready = Queue_io_enq_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 299:17]
  wire [29:0] _T_18 = auto_register_in_ar_valid ? auto_register_in_ar_bits_addr : auto_register_in_aw_bits_addr; // @[RegisterRouter.scala 48:19]
  wire [1:0] _T_58 = _T_18[3:2] & 2'h2; // @[RegisterRouter.scala 59:16]
  wire  _T_60 = _T_58 == 2'h0; // @[RegisterRouter.scala 59:16]
  wire  _T_12 = _T_54_ready & _T_11; // @[RegisterRouter.scala 42:26]
  wire [1:0] _T_21 = 2'h1 << auto_register_in_ar_bits_size[0]; // @[OneHot.scala 65:12]
  wire [1:0] _T_23 = _T_21 | 2'h1; // @[Misc.scala 200:81]
  wire  _T_24 = auto_register_in_ar_bits_size >= 3'h2; // @[Misc.scala 204:21]
  wire  _T_27 = ~auto_register_in_ar_bits_addr[1]; // @[Misc.scala 209:20]
  wire  _T_29 = _T_23[1] & _T_27; // @[Misc.scala 213:38]
  wire  _T_30 = _T_24 | _T_29; // @[Misc.scala 213:29]
  wire  _T_32 = _T_23[1] & auto_register_in_ar_bits_addr[1]; // @[Misc.scala 213:38]
  wire  _T_33 = _T_24 | _T_32; // @[Misc.scala 213:29]
  wire  _T_36 = ~auto_register_in_ar_bits_addr[0]; // @[Misc.scala 209:20]
  wire  _T_37 = _T_27 & _T_36; // @[Misc.scala 212:27]
  wire  _T_38 = _T_23[0] & _T_37; // @[Misc.scala 213:38]
  wire  _T_39 = _T_30 | _T_38; // @[Misc.scala 213:29]
  wire  _T_40 = _T_27 & auto_register_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  wire  _T_41 = _T_23[0] & _T_40; // @[Misc.scala 213:38]
  wire  _T_42 = _T_30 | _T_41; // @[Misc.scala 213:29]
  wire  _T_43 = auto_register_in_ar_bits_addr[1] & _T_36; // @[Misc.scala 212:27]
  wire  _T_44 = _T_23[0] & _T_43; // @[Misc.scala 213:38]
  wire  _T_45 = _T_33 | _T_44; // @[Misc.scala 213:29]
  wire  _T_46 = auto_register_in_ar_bits_addr[1] & auto_register_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  wire  _T_47 = _T_23[0] & _T_46; // @[Misc.scala 213:38]
  wire  _T_48 = _T_33 | _T_47; // @[Misc.scala 213:29]
  wire [3:0] _T_51 = {_T_48,_T_45,_T_42,_T_39}; // @[Cat.scala 29:58]
  wire [3:0] _T_53 = auto_register_in_ar_valid ? _T_51 : auto_register_in_w_bits_strb; // @[RegisterRouter.scala 54:25]
  wire [7:0] _T_72 = _T_53[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_74 = _T_53[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_76 = _T_53[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_78 = _T_53[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_81 = {_T_78,_T_76,_T_74,_T_72}; // @[Cat.scala 29:58]
  wire  _T_153 = _T_10 & _T_54_ready; // @[RegisterRouter.scala 59:16]
  wire [1:0] _T_147 = 2'h1 << _T_18[2]; // @[OneHot.scala 58:35]
  wire  _T_170 = _T_153 & _T_11; // @[RegisterRouter.scala 59:16]
  wire  _T_177 = _T_170 & _T_147[1]; // @[RegisterRouter.scala 59:16]
  wire  _T_178 = _T_177 & _T_60; // @[RegisterRouter.scala 59:16]
  wire  _T_107 = _T_178 & _T_81[0]; // @[RegisterRouter.scala 59:16]
  wire  _GEN_18 = _T_107 ? auto_register_in_w_bits_data[0] : sels_1; // @[RegField.scala 134:88]
  wire  _T_172 = _T_170 & _T_147[0]; // @[RegisterRouter.scala 59:16]
  wire  _T_173 = _T_172 & _T_60; // @[RegisterRouter.scala 59:16]
  wire  _T_130 = _T_173 & _T_81[0]; // @[RegisterRouter.scala 59:16]
  wire  _GEN_19 = _T_130 ? auto_register_in_w_bits_data[0] : sels_0; // @[RegField.scala 134:88]
  wire  _GEN_29 = _T_18[2] ? _T_60 : _T_60; // @[MuxLiteral.scala 48:10]
  wire  _GEN_31 = _T_18[2] ? sels_1 : sels_0; // @[MuxLiteral.scala 48:10]
  wire  _T_227 = _GEN_29 & _GEN_31; // @[RegisterRouter.scala 59:16]
  wire  _T_228_bits_read = Queue_io_deq_bits_read; // @[Decoupled.scala 317:19 Decoupled.scala 318:14]
  wire  _T_228_valid = Queue_io_deq_valid; // @[Decoupled.scala 317:19 Decoupled.scala 319:15]
  wire  _T_231 = ~_T_228_bits_read; // @[RegisterRouter.scala 65:29]
  Queue Queue ( // @[Decoupled.scala 296:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_read(Queue_io_enq_bits_read),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_extra(Queue_io_enq_bits_extra),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_read(Queue_io_deq_bits_read),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_extra(Queue_io_deq_bits_extra)
  );
  assign auto_register_in_aw_ready = _T_12 & auto_register_in_w_valid; // @[LazyModule.scala 173:31]
  assign auto_register_in_w_ready = _T_12 & auto_register_in_aw_valid; // @[LazyModule.scala 173:31]
  assign auto_register_in_b_valid = _T_228_valid & _T_231; // @[LazyModule.scala 173:31]
  assign auto_register_in_b_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_register_in_ar_ready = Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_register_in_r_valid = _T_228_valid & _T_228_bits_read; // @[LazyModule.scala 173:31]
  assign auto_register_in_r_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_register_in_r_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 173:31]
  assign auto_stream_in_ready = _T_7 ? auto_stream_out_1_ready : _T_3; // @[LazyModule.scala 173:31]
  assign auto_stream_out_1_valid = _T_7 & auto_stream_in_valid; // @[LazyModule.scala 173:49]
  assign auto_stream_out_1_bits_data = auto_stream_in_bits_data; // @[LazyModule.scala 173:49]
  assign auto_stream_out_1_bits_last = auto_stream_in_bits_last; // @[LazyModule.scala 173:49]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_register_in_ar_valid | _T_9; // @[Decoupled.scala 297:22]
  assign Queue_io_enq_bits_read = auto_register_in_ar_valid; // @[Decoupled.scala 298:21]
  assign Queue_io_enq_bits_data = {{31'd0}, _T_227}; // @[Decoupled.scala 298:21]
  assign Queue_io_enq_bits_extra = auto_register_in_ar_valid ? auto_register_in_ar_bits_id : auto_register_in_aw_bits_id; // @[Decoupled.scala 298:21]
  assign Queue_io_deq_ready = _T_228_bits_read ? auto_register_in_r_ready : auto_register_in_b_ready; // @[Decoupled.scala 320:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  sels_0 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  sels_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    sels_0 <= reset | _GEN_19;
    sels_1 <= reset | _GEN_18;
  end
endmodule
module Queue_15(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [15:0] io_enq_bits_real,
  input  [15:0] io_enq_bits_imag,
  input         io_deq_ready,
  output        io_deq_valid,
  output [15:0] io_deq_bits_real,
  output [15:0] io_deq_bits_imag
);
  reg [15:0] _T_4_real [0:4]; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_0;
  wire [15:0] _T_4_real__T_26_data; // @[Decoupled.scala 218:24]
  wire [2:0] _T_4_real__T_26_addr; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_1;
  wire [15:0] _T_4_real__T_16_data; // @[Decoupled.scala 218:24]
  wire [2:0] _T_4_real__T_16_addr; // @[Decoupled.scala 218:24]
  wire  _T_4_real__T_16_mask; // @[Decoupled.scala 218:24]
  wire  _T_4_real__T_16_en; // @[Decoupled.scala 218:24]
  reg [15:0] _T_4_imag [0:4]; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_2;
  wire [15:0] _T_4_imag__T_26_data; // @[Decoupled.scala 218:24]
  wire [2:0] _T_4_imag__T_26_addr; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_3;
  wire [15:0] _T_4_imag__T_16_data; // @[Decoupled.scala 218:24]
  wire [2:0] _T_4_imag__T_16_addr; // @[Decoupled.scala 218:24]
  wire  _T_4_imag__T_16_mask; // @[Decoupled.scala 218:24]
  wire  _T_4_imag__T_16_en; // @[Decoupled.scala 218:24]
  reg [2:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_4;
  reg [2:0] value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  reg  _T_5; // @[Decoupled.scala 221:35]
  reg [31:0] _RAND_6;
  wire  _T_6 = value == value_1; // @[Decoupled.scala 223:41]
  wire  _T_7 = ~_T_5; // @[Decoupled.scala 224:36]
  wire  _T_8 = _T_6 & _T_7; // @[Decoupled.scala 224:33]
  wire  _T_9 = _T_6 & _T_5; // @[Decoupled.scala 225:32]
  wire  _T_10 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  _T_12 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire  wrap = value == 3'h4; // @[Counter.scala 38:24]
  wire [2:0] _T_18 = value + 3'h1; // @[Counter.scala 39:22]
  wire  wrap_1 = value_1 == 3'h4; // @[Counter.scala 38:24]
  wire [2:0] _T_20 = value_1 + 3'h1; // @[Counter.scala 39:22]
  wire  _T_21 = _T_10 != _T_12; // @[Decoupled.scala 236:16]
  assign _T_4_real__T_26_addr = value_1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_4_real__T_26_data = _T_4_real[_T_4_real__T_26_addr]; // @[Decoupled.scala 218:24]
  `else
  assign _T_4_real__T_26_data = _T_4_real__T_26_addr >= 3'h5 ? _RAND_1[15:0] : _T_4_real[_T_4_real__T_26_addr]; // @[Decoupled.scala 218:24]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_4_real__T_16_data = io_enq_bits_real;
  assign _T_4_real__T_16_addr = value;
  assign _T_4_real__T_16_mask = 1'h1;
  assign _T_4_real__T_16_en = io_enq_ready & io_enq_valid;
  assign _T_4_imag__T_26_addr = value_1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_4_imag__T_26_data = _T_4_imag[_T_4_imag__T_26_addr]; // @[Decoupled.scala 218:24]
  `else
  assign _T_4_imag__T_26_data = _T_4_imag__T_26_addr >= 3'h5 ? _RAND_3[15:0] : _T_4_imag[_T_4_imag__T_26_addr]; // @[Decoupled.scala 218:24]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_4_imag__T_16_data = io_enq_bits_imag;
  assign _T_4_imag__T_16_addr = value;
  assign _T_4_imag__T_16_mask = 1'h1;
  assign _T_4_imag__T_16_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~_T_9; // @[Decoupled.scala 241:16]
  assign io_deq_valid = ~_T_8; // @[Decoupled.scala 240:16]
  assign io_deq_bits_real = _T_4_real__T_26_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_imag = _T_4_imag__T_26_data; // @[Decoupled.scala 242:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 5; initvar = initvar+1)
    _T_4_real[initvar] = _RAND_0[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  _RAND_2 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 5; initvar = initvar+1)
    _T_4_imag[initvar] = _RAND_2[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  value = _RAND_4[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value_1 = _RAND_5[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_5 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T_4_real__T_16_en & _T_4_real__T_16_mask) begin
      _T_4_real[_T_4_real__T_16_addr] <= _T_4_real__T_16_data; // @[Decoupled.scala 218:24]
    end
    if(_T_4_imag__T_16_en & _T_4_imag__T_16_mask) begin
      _T_4_imag[_T_4_imag__T_16_addr] <= _T_4_imag__T_16_data; // @[Decoupled.scala 218:24]
    end
    if (reset) begin
      value <= 3'h0;
    end else if (_T_10) begin
      if (wrap) begin
        value <= 3'h0;
      end else begin
        value <= _T_18;
      end
    end
    if (reset) begin
      value_1 <= 3'h0;
    end else if (_T_12) begin
      if (wrap_1) begin
        value_1 <= 3'h0;
      end else begin
        value_1 <= _T_20;
      end
    end
    if (reset) begin
      _T_5 <= 1'h0;
    end else if (_T_21) begin
      _T_5 <= _T_10;
    end
  end
endmodule
module Queue_16(
  input   clock,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input   io_enq_bits,
  input   io_deq_ready,
  output  io_deq_valid,
  output  io_deq_bits
);
  reg  _T [0:4]; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_0;
  wire  _T__T_18_data; // @[Decoupled.scala 218:24]
  wire [2:0] _T__T_18_addr; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_1;
  wire  _T__T_10_data; // @[Decoupled.scala 218:24]
  wire [2:0] _T__T_10_addr; // @[Decoupled.scala 218:24]
  wire  _T__T_10_mask; // @[Decoupled.scala 218:24]
  wire  _T__T_10_en; // @[Decoupled.scala 218:24]
  reg [2:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_2;
  reg [2:0] value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_3;
  reg  _T_1; // @[Decoupled.scala 221:35]
  reg [31:0] _RAND_4;
  wire  _T_2 = value == value_1; // @[Decoupled.scala 223:41]
  wire  _T_3 = ~_T_1; // @[Decoupled.scala 224:36]
  wire  _T_4 = _T_2 & _T_3; // @[Decoupled.scala 224:33]
  wire  _T_5 = _T_2 & _T_1; // @[Decoupled.scala 225:32]
  wire  _T_6 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  _T_8 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire  wrap = value == 3'h4; // @[Counter.scala 38:24]
  wire [2:0] _T_12 = value + 3'h1; // @[Counter.scala 39:22]
  wire  wrap_1 = value_1 == 3'h4; // @[Counter.scala 38:24]
  wire [2:0] _T_14 = value_1 + 3'h1; // @[Counter.scala 39:22]
  wire  _T_15 = _T_6 != _T_8; // @[Decoupled.scala 236:16]
  assign _T__T_18_addr = value_1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__T_18_data = _T[_T__T_18_addr]; // @[Decoupled.scala 218:24]
  `else
  assign _T__T_18_data = _T__T_18_addr >= 3'h5 ? _RAND_1[0:0] : _T[_T__T_18_addr]; // @[Decoupled.scala 218:24]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__T_10_data = io_enq_bits;
  assign _T__T_10_addr = value;
  assign _T__T_10_mask = 1'h1;
  assign _T__T_10_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~_T_5; // @[Decoupled.scala 241:16]
  assign io_deq_valid = ~_T_4; // @[Decoupled.scala 240:16]
  assign io_deq_bits = _T__T_18_data; // @[Decoupled.scala 242:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 5; initvar = initvar+1)
    _T[initvar] = _RAND_0[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  value = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  value_1 = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T__T_10_en & _T__T_10_mask) begin
      _T[_T__T_10_addr] <= _T__T_10_data; // @[Decoupled.scala 218:24]
    end
    if (reset) begin
      value <= 3'h0;
    end else if (_T_6) begin
      if (wrap) begin
        value <= 3'h0;
      end else begin
        value <= _T_12;
      end
    end
    if (reset) begin
      value_1 <= 3'h0;
    end else if (_T_8) begin
      if (wrap_1) begin
        value_1 <= 3'h0;
      end else begin
        value_1 <= _T_14;
      end
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else if (_T_15) begin
      _T_1 <= _T_6;
    end
  end
endmodule
module LogMagMux(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [15:0] io_in_bits_real,
  input  [15:0] io_in_bits_imag,
  input         io_lastIn,
  input         io_out_ready,
  output        io_out_valid,
  output [15:0] io_out_bits_real,
  output [15:0] io_out_bits_imag,
  input  [1:0]  io_sel,
  output        io_lastOut
);
  wire  Queue_clock; // @[Skid.scala 21:23]
  wire  Queue_reset; // @[Skid.scala 21:23]
  wire  Queue_io_enq_ready; // @[Skid.scala 21:23]
  wire  Queue_io_enq_valid; // @[Skid.scala 21:23]
  wire [15:0] Queue_io_enq_bits_real; // @[Skid.scala 21:23]
  wire [15:0] Queue_io_enq_bits_imag; // @[Skid.scala 21:23]
  wire  Queue_io_deq_ready; // @[Skid.scala 21:23]
  wire  Queue_io_deq_valid; // @[Skid.scala 21:23]
  wire [15:0] Queue_io_deq_bits_real; // @[Skid.scala 21:23]
  wire [15:0] Queue_io_deq_bits_imag; // @[Skid.scala 21:23]
  wire  Queue_1_clock; // @[Skid.scala 21:23]
  wire  Queue_1_reset; // @[Skid.scala 21:23]
  wire  Queue_1_io_enq_ready; // @[Skid.scala 21:23]
  wire  Queue_1_io_enq_valid; // @[Skid.scala 21:23]
  wire  Queue_1_io_enq_bits; // @[Skid.scala 21:23]
  wire  Queue_1_io_deq_ready; // @[Skid.scala 21:23]
  wire  Queue_1_io_deq_valid; // @[Skid.scala 21:23]
  wire  Queue_1_io_deq_bits; // @[Skid.scala 21:23]
  wire [15:0] _T_7 = 16'sh0 - $signed(io_in_bits_real); // @[FixedPointTypeClass.scala 30:68]
  wire [15:0] absInReal = io_in_bits_real[15] ? $signed(_T_7) : $signed(io_in_bits_real); // @[FixedPointTypeClass.scala 247:8]
  wire [15:0] _T_11 = 16'sh0 - $signed(io_in_bits_imag); // @[FixedPointTypeClass.scala 30:68]
  wire [15:0] absInImag = io_in_bits_imag[15] ? $signed(_T_11) : $signed(io_in_bits_imag); // @[FixedPointTypeClass.scala 247:8]
  wire  _T_12 = $signed(absInReal) > $signed(absInImag); // @[FixedPointTypeClass.scala 55:59]
  wire [15:0] u = _T_12 ? $signed(absInReal) : $signed(absInImag); // @[Order.scala 56:31]
  wire  _T_13 = $signed(absInReal) < $signed(absInImag); // @[FixedPointTypeClass.scala 53:59]
  wire [15:0] v = _T_13 ? $signed(absInReal) : $signed(absInImag); // @[Order.scala 55:31]
  wire [12:0] _T_14 = v[15:3]; // @[FixedPointTypeClass.scala 117:50]
  wire [15:0] _GEN_559 = {{3{_T_14[12]}},_T_14}; // @[FixedPointTypeClass.scala 24:22]
  reg [16:0] _T_16; // @[Reg.scala 15:16]
  reg [31:0] _RAND_0;
  reg [16:0] jplMagOp1; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1;
  wire [12:0] _T_17 = u[15:3]; // @[FixedPointTypeClass.scala 117:50]
  wire [15:0] _GEN_560 = {{3{_T_17[12]}},_T_17}; // @[FixedPointTypeClass.scala 33:22]
  reg [16:0] tmpOp2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2;
  reg [14:0] _T_20; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3;
  wire [16:0] _GEN_561 = {{2{_T_20[14]}},_T_20}; // @[FixedPointTypeClass.scala 24:22]
  reg [17:0] jplMagOp2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4;
  reg [31:0] _T_23; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5;
  wire [32:0] _T_24 = {$signed(_T_23), 1'h0}; // @[FixedPointTypeClass.scala 153:43]
  reg [31:0] _T_26; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6;
  wire [32:0] _T_27 = {$signed(_T_26), 1'h0}; // @[FixedPointTypeClass.scala 153:43]
  reg [33:0] _T_29; // @[Reg.scala 15:16]
  reg [63:0] _RAND_7;
  reg [33:0] _T_30; // @[Reg.scala 15:16]
  reg [63:0] _RAND_8;
  reg [33:0] _T_31; // @[Reg.scala 15:16]
  reg [63:0] _RAND_9;
  wire [17:0] _GEN_562 = {{1{jplMagOp1[16]}},jplMagOp1}; // @[FixedPointTypeClass.scala 55:59]
  wire  _T_32 = $signed(_GEN_562) > $signed(jplMagOp2); // @[FixedPointTypeClass.scala 55:59]
  reg [17:0] _T_33; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10;
  reg [17:0] jplMag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11;
  wire [17:0] _T_34 = jplMag; // @[LogMagMux.scala 113:35]
  wire  _T_37 = _T_34[17:16] != 2'h0; // @[CircuitMath.scala 37:22]
  wire  _T_41 = _T_34[15:8] != 8'h0; // @[CircuitMath.scala 37:22]
  wire  _T_44 = _T_34[15:12] != 4'h0; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_48 = _T_34[14] ? 2'h2 : {{1'd0}, _T_34[13]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_49 = _T_34[15] ? 2'h3 : _T_48; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_53 = _T_34[10] ? 2'h2 : {{1'd0}, _T_34[9]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_54 = _T_34[11] ? 2'h3 : _T_53; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_55 = _T_44 ? _T_49 : _T_54; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_56 = {_T_44,_T_55}; // @[Cat.scala 29:58]
  wire  _T_59 = _T_34[7:4] != 4'h0; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_63 = _T_34[6] ? 2'h2 : {{1'd0}, _T_34[5]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_64 = _T_34[7] ? 2'h3 : _T_63; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_68 = _T_34[2] ? 2'h2 : {{1'd0}, _T_34[1]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_69 = _T_34[3] ? 2'h3 : _T_68; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_70 = _T_59 ? _T_64 : _T_69; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_71 = {_T_59,_T_70}; // @[Cat.scala 29:58]
  wire [2:0] _T_72 = _T_41 ? _T_56 : _T_71; // @[CircuitMath.scala 38:21]
  wire [3:0] _T_73 = {_T_41,_T_72}; // @[Cat.scala 29:58]
  wire [3:0] _T_74 = _T_37 ? {{3'd0}, _T_34[17]} : _T_73; // @[CircuitMath.scala 38:21]
  wire [4:0] logUInt = {_T_37,_T_74}; // @[Cat.scala 29:58]
  wire [17:0] _T_589 = _T_32 ? $signed({{1{jplMagOp1[16]}},jplMagOp1}) : $signed(jplMagOp2); // @[LogMagMux.scala 131:50]
  wire [31:0] _T_590 = 32'h1 << logUInt; // @[UIntTypeClass.scala 124:39]
  reg [17:0] noLeadOne; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12;
  wire [4:0] _T_596 = 5'h10 - logUInt; // @[LogMagMux.scala 132:44]
  reg [4:0] shiftNum; // @[Reg.scala 15:16]
  reg [31:0] _RAND_13;
  wire [48:0] _GEN_563 = {{31'd0}, noLeadOne}; // @[UIntTypeClass.scala 124:39]
  wire [48:0] _T_599 = _GEN_563 << shiftNum; // @[UIntTypeClass.scala 124:39]
  wire [8:0] logLookUpAddr = _T_599[14:6]; // @[LogMagMux.scala 134:74]
  wire [9:0] _GEN_15 = 9'h1 == logLookUpAddr ? $signed(10'sh1) : $signed(10'sh0); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_16 = 9'h2 == logLookUpAddr ? $signed(10'sh3) : $signed(_GEN_15); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_17 = 9'h3 == logLookUpAddr ? $signed(10'sh4) : $signed(_GEN_16); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_18 = 9'h4 == logLookUpAddr ? $signed(10'sh6) : $signed(_GEN_17); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_19 = 9'h5 == logLookUpAddr ? $signed(10'sh7) : $signed(_GEN_18); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_20 = 9'h6 == logLookUpAddr ? $signed(10'sh9) : $signed(_GEN_19); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_21 = 9'h7 == logLookUpAddr ? $signed(10'sha) : $signed(_GEN_20); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_22 = 9'h8 == logLookUpAddr ? $signed(10'shb) : $signed(_GEN_21); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_23 = 9'h9 == logLookUpAddr ? $signed(10'shd) : $signed(_GEN_22); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_24 = 9'ha == logLookUpAddr ? $signed(10'she) : $signed(_GEN_23); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_25 = 9'hb == logLookUpAddr ? $signed(10'sh10) : $signed(_GEN_24); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_26 = 9'hc == logLookUpAddr ? $signed(10'sh11) : $signed(_GEN_25); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_27 = 9'hd == logLookUpAddr ? $signed(10'sh13) : $signed(_GEN_26); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_28 = 9'he == logLookUpAddr ? $signed(10'sh14) : $signed(_GEN_27); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_29 = 9'hf == logLookUpAddr ? $signed(10'sh15) : $signed(_GEN_28); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_30 = 9'h10 == logLookUpAddr ? $signed(10'sh17) : $signed(_GEN_29); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_31 = 9'h11 == logLookUpAddr ? $signed(10'sh18) : $signed(_GEN_30); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_32 = 9'h12 == logLookUpAddr ? $signed(10'sh1a) : $signed(_GEN_31); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_33 = 9'h13 == logLookUpAddr ? $signed(10'sh1b) : $signed(_GEN_32); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_34 = 9'h14 == logLookUpAddr ? $signed(10'sh1c) : $signed(_GEN_33); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_35 = 9'h15 == logLookUpAddr ? $signed(10'sh1e) : $signed(_GEN_34); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_36 = 9'h16 == logLookUpAddr ? $signed(10'sh1f) : $signed(_GEN_35); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_37 = 9'h17 == logLookUpAddr ? $signed(10'sh20) : $signed(_GEN_36); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_38 = 9'h18 == logLookUpAddr ? $signed(10'sh22) : $signed(_GEN_37); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_39 = 9'h19 == logLookUpAddr ? $signed(10'sh23) : $signed(_GEN_38); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_40 = 9'h1a == logLookUpAddr ? $signed(10'sh25) : $signed(_GEN_39); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_41 = 9'h1b == logLookUpAddr ? $signed(10'sh26) : $signed(_GEN_40); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_42 = 9'h1c == logLookUpAddr ? $signed(10'sh27) : $signed(_GEN_41); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_43 = 9'h1d == logLookUpAddr ? $signed(10'sh29) : $signed(_GEN_42); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_44 = 9'h1e == logLookUpAddr ? $signed(10'sh2a) : $signed(_GEN_43); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_45 = 9'h1f == logLookUpAddr ? $signed(10'sh2b) : $signed(_GEN_44); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_46 = 9'h20 == logLookUpAddr ? $signed(10'sh2d) : $signed(_GEN_45); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_47 = 9'h21 == logLookUpAddr ? $signed(10'sh2e) : $signed(_GEN_46); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_48 = 9'h22 == logLookUpAddr ? $signed(10'sh2f) : $signed(_GEN_47); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_49 = 9'h23 == logLookUpAddr ? $signed(10'sh31) : $signed(_GEN_48); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_50 = 9'h24 == logLookUpAddr ? $signed(10'sh32) : $signed(_GEN_49); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_51 = 9'h25 == logLookUpAddr ? $signed(10'sh34) : $signed(_GEN_50); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_52 = 9'h26 == logLookUpAddr ? $signed(10'sh35) : $signed(_GEN_51); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_53 = 9'h27 == logLookUpAddr ? $signed(10'sh36) : $signed(_GEN_52); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_54 = 9'h28 == logLookUpAddr ? $signed(10'sh38) : $signed(_GEN_53); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_55 = 9'h29 == logLookUpAddr ? $signed(10'sh39) : $signed(_GEN_54); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_56 = 9'h2a == logLookUpAddr ? $signed(10'sh3a) : $signed(_GEN_55); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_57 = 9'h2b == logLookUpAddr ? $signed(10'sh3c) : $signed(_GEN_56); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_58 = 9'h2c == logLookUpAddr ? $signed(10'sh3d) : $signed(_GEN_57); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_59 = 9'h2d == logLookUpAddr ? $signed(10'sh3e) : $signed(_GEN_58); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_60 = 9'h2e == logLookUpAddr ? $signed(10'sh40) : $signed(_GEN_59); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_61 = 9'h2f == logLookUpAddr ? $signed(10'sh41) : $signed(_GEN_60); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_62 = 9'h30 == logLookUpAddr ? $signed(10'sh42) : $signed(_GEN_61); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_63 = 9'h31 == logLookUpAddr ? $signed(10'sh44) : $signed(_GEN_62); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_64 = 9'h32 == logLookUpAddr ? $signed(10'sh45) : $signed(_GEN_63); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_65 = 9'h33 == logLookUpAddr ? $signed(10'sh46) : $signed(_GEN_64); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_66 = 9'h34 == logLookUpAddr ? $signed(10'sh47) : $signed(_GEN_65); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_67 = 9'h35 == logLookUpAddr ? $signed(10'sh49) : $signed(_GEN_66); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_68 = 9'h36 == logLookUpAddr ? $signed(10'sh4a) : $signed(_GEN_67); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_69 = 9'h37 == logLookUpAddr ? $signed(10'sh4b) : $signed(_GEN_68); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_70 = 9'h38 == logLookUpAddr ? $signed(10'sh4d) : $signed(_GEN_69); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_71 = 9'h39 == logLookUpAddr ? $signed(10'sh4e) : $signed(_GEN_70); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_72 = 9'h3a == logLookUpAddr ? $signed(10'sh4f) : $signed(_GEN_71); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_73 = 9'h3b == logLookUpAddr ? $signed(10'sh51) : $signed(_GEN_72); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_74 = 9'h3c == logLookUpAddr ? $signed(10'sh52) : $signed(_GEN_73); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_75 = 9'h3d == logLookUpAddr ? $signed(10'sh53) : $signed(_GEN_74); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_76 = 9'h3e == logLookUpAddr ? $signed(10'sh54) : $signed(_GEN_75); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_77 = 9'h3f == logLookUpAddr ? $signed(10'sh56) : $signed(_GEN_76); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_78 = 9'h40 == logLookUpAddr ? $signed(10'sh57) : $signed(_GEN_77); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_79 = 9'h41 == logLookUpAddr ? $signed(10'sh58) : $signed(_GEN_78); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_80 = 9'h42 == logLookUpAddr ? $signed(10'sh5a) : $signed(_GEN_79); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_81 = 9'h43 == logLookUpAddr ? $signed(10'sh5b) : $signed(_GEN_80); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_82 = 9'h44 == logLookUpAddr ? $signed(10'sh5c) : $signed(_GEN_81); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_83 = 9'h45 == logLookUpAddr ? $signed(10'sh5d) : $signed(_GEN_82); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_84 = 9'h46 == logLookUpAddr ? $signed(10'sh5f) : $signed(_GEN_83); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_85 = 9'h47 == logLookUpAddr ? $signed(10'sh60) : $signed(_GEN_84); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_86 = 9'h48 == logLookUpAddr ? $signed(10'sh61) : $signed(_GEN_85); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_87 = 9'h49 == logLookUpAddr ? $signed(10'sh62) : $signed(_GEN_86); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_88 = 9'h4a == logLookUpAddr ? $signed(10'sh64) : $signed(_GEN_87); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_89 = 9'h4b == logLookUpAddr ? $signed(10'sh65) : $signed(_GEN_88); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_90 = 9'h4c == logLookUpAddr ? $signed(10'sh66) : $signed(_GEN_89); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_91 = 9'h4d == logLookUpAddr ? $signed(10'sh67) : $signed(_GEN_90); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_92 = 9'h4e == logLookUpAddr ? $signed(10'sh69) : $signed(_GEN_91); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_93 = 9'h4f == logLookUpAddr ? $signed(10'sh6a) : $signed(_GEN_92); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_94 = 9'h50 == logLookUpAddr ? $signed(10'sh6b) : $signed(_GEN_93); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_95 = 9'h51 == logLookUpAddr ? $signed(10'sh6c) : $signed(_GEN_94); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_96 = 9'h52 == logLookUpAddr ? $signed(10'sh6e) : $signed(_GEN_95); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_97 = 9'h53 == logLookUpAddr ? $signed(10'sh6f) : $signed(_GEN_96); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_98 = 9'h54 == logLookUpAddr ? $signed(10'sh70) : $signed(_GEN_97); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_99 = 9'h55 == logLookUpAddr ? $signed(10'sh71) : $signed(_GEN_98); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_100 = 9'h56 == logLookUpAddr ? $signed(10'sh73) : $signed(_GEN_99); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_101 = 9'h57 == logLookUpAddr ? $signed(10'sh74) : $signed(_GEN_100); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_102 = 9'h58 == logLookUpAddr ? $signed(10'sh75) : $signed(_GEN_101); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_103 = 9'h59 == logLookUpAddr ? $signed(10'sh76) : $signed(_GEN_102); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_104 = 9'h5a == logLookUpAddr ? $signed(10'sh78) : $signed(_GEN_103); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_105 = 9'h5b == logLookUpAddr ? $signed(10'sh79) : $signed(_GEN_104); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_106 = 9'h5c == logLookUpAddr ? $signed(10'sh7a) : $signed(_GEN_105); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_107 = 9'h5d == logLookUpAddr ? $signed(10'sh7b) : $signed(_GEN_106); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_108 = 9'h5e == logLookUpAddr ? $signed(10'sh7d) : $signed(_GEN_107); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_109 = 9'h5f == logLookUpAddr ? $signed(10'sh7e) : $signed(_GEN_108); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_110 = 9'h60 == logLookUpAddr ? $signed(10'sh7f) : $signed(_GEN_109); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_111 = 9'h61 == logLookUpAddr ? $signed(10'sh80) : $signed(_GEN_110); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_112 = 9'h62 == logLookUpAddr ? $signed(10'sh81) : $signed(_GEN_111); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_113 = 9'h63 == logLookUpAddr ? $signed(10'sh83) : $signed(_GEN_112); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_114 = 9'h64 == logLookUpAddr ? $signed(10'sh84) : $signed(_GEN_113); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_115 = 9'h65 == logLookUpAddr ? $signed(10'sh85) : $signed(_GEN_114); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_116 = 9'h66 == logLookUpAddr ? $signed(10'sh86) : $signed(_GEN_115); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_117 = 9'h67 == logLookUpAddr ? $signed(10'sh87) : $signed(_GEN_116); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_118 = 9'h68 == logLookUpAddr ? $signed(10'sh89) : $signed(_GEN_117); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_119 = 9'h69 == logLookUpAddr ? $signed(10'sh8a) : $signed(_GEN_118); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_120 = 9'h6a == logLookUpAddr ? $signed(10'sh8b) : $signed(_GEN_119); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_121 = 9'h6b == logLookUpAddr ? $signed(10'sh8c) : $signed(_GEN_120); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_122 = 9'h6c == logLookUpAddr ? $signed(10'sh8d) : $signed(_GEN_121); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_123 = 9'h6d == logLookUpAddr ? $signed(10'sh8f) : $signed(_GEN_122); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_124 = 9'h6e == logLookUpAddr ? $signed(10'sh90) : $signed(_GEN_123); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_125 = 9'h6f == logLookUpAddr ? $signed(10'sh91) : $signed(_GEN_124); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_126 = 9'h70 == logLookUpAddr ? $signed(10'sh92) : $signed(_GEN_125); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_127 = 9'h71 == logLookUpAddr ? $signed(10'sh93) : $signed(_GEN_126); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_128 = 9'h72 == logLookUpAddr ? $signed(10'sh94) : $signed(_GEN_127); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_129 = 9'h73 == logLookUpAddr ? $signed(10'sh96) : $signed(_GEN_128); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_130 = 9'h74 == logLookUpAddr ? $signed(10'sh97) : $signed(_GEN_129); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_131 = 9'h75 == logLookUpAddr ? $signed(10'sh98) : $signed(_GEN_130); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_132 = 9'h76 == logLookUpAddr ? $signed(10'sh99) : $signed(_GEN_131); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_133 = 9'h77 == logLookUpAddr ? $signed(10'sh9a) : $signed(_GEN_132); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_134 = 9'h78 == logLookUpAddr ? $signed(10'sh9c) : $signed(_GEN_133); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_135 = 9'h79 == logLookUpAddr ? $signed(10'sh9d) : $signed(_GEN_134); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_136 = 9'h7a == logLookUpAddr ? $signed(10'sh9e) : $signed(_GEN_135); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_137 = 9'h7b == logLookUpAddr ? $signed(10'sh9f) : $signed(_GEN_136); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_138 = 9'h7c == logLookUpAddr ? $signed(10'sha0) : $signed(_GEN_137); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_139 = 9'h7d == logLookUpAddr ? $signed(10'sha1) : $signed(_GEN_138); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_140 = 9'h7e == logLookUpAddr ? $signed(10'sha3) : $signed(_GEN_139); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_141 = 9'h7f == logLookUpAddr ? $signed(10'sha4) : $signed(_GEN_140); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_142 = 9'h80 == logLookUpAddr ? $signed(10'sha5) : $signed(_GEN_141); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_143 = 9'h81 == logLookUpAddr ? $signed(10'sha6) : $signed(_GEN_142); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_144 = 9'h82 == logLookUpAddr ? $signed(10'sha7) : $signed(_GEN_143); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_145 = 9'h83 == logLookUpAddr ? $signed(10'sha8) : $signed(_GEN_144); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_146 = 9'h84 == logLookUpAddr ? $signed(10'sha9) : $signed(_GEN_145); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_147 = 9'h85 == logLookUpAddr ? $signed(10'shab) : $signed(_GEN_146); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_148 = 9'h86 == logLookUpAddr ? $signed(10'shac) : $signed(_GEN_147); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_149 = 9'h87 == logLookUpAddr ? $signed(10'shad) : $signed(_GEN_148); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_150 = 9'h88 == logLookUpAddr ? $signed(10'shae) : $signed(_GEN_149); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_151 = 9'h89 == logLookUpAddr ? $signed(10'shaf) : $signed(_GEN_150); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_152 = 9'h8a == logLookUpAddr ? $signed(10'shb0) : $signed(_GEN_151); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_153 = 9'h8b == logLookUpAddr ? $signed(10'shb1) : $signed(_GEN_152); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_154 = 9'h8c == logLookUpAddr ? $signed(10'shb3) : $signed(_GEN_153); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_155 = 9'h8d == logLookUpAddr ? $signed(10'shb4) : $signed(_GEN_154); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_156 = 9'h8e == logLookUpAddr ? $signed(10'shb5) : $signed(_GEN_155); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_157 = 9'h8f == logLookUpAddr ? $signed(10'shb6) : $signed(_GEN_156); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_158 = 9'h90 == logLookUpAddr ? $signed(10'shb7) : $signed(_GEN_157); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_159 = 9'h91 == logLookUpAddr ? $signed(10'shb8) : $signed(_GEN_158); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_160 = 9'h92 == logLookUpAddr ? $signed(10'shb9) : $signed(_GEN_159); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_161 = 9'h93 == logLookUpAddr ? $signed(10'shba) : $signed(_GEN_160); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_162 = 9'h94 == logLookUpAddr ? $signed(10'shbc) : $signed(_GEN_161); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_163 = 9'h95 == logLookUpAddr ? $signed(10'shbd) : $signed(_GEN_162); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_164 = 9'h96 == logLookUpAddr ? $signed(10'shbe) : $signed(_GEN_163); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_165 = 9'h97 == logLookUpAddr ? $signed(10'shbf) : $signed(_GEN_164); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_166 = 9'h98 == logLookUpAddr ? $signed(10'shc0) : $signed(_GEN_165); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_167 = 9'h99 == logLookUpAddr ? $signed(10'shc1) : $signed(_GEN_166); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_168 = 9'h9a == logLookUpAddr ? $signed(10'shc2) : $signed(_GEN_167); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_169 = 9'h9b == logLookUpAddr ? $signed(10'shc3) : $signed(_GEN_168); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_170 = 9'h9c == logLookUpAddr ? $signed(10'shc4) : $signed(_GEN_169); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_171 = 9'h9d == logLookUpAddr ? $signed(10'shc6) : $signed(_GEN_170); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_172 = 9'h9e == logLookUpAddr ? $signed(10'shc7) : $signed(_GEN_171); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_173 = 9'h9f == logLookUpAddr ? $signed(10'shc8) : $signed(_GEN_172); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_174 = 9'ha0 == logLookUpAddr ? $signed(10'shc9) : $signed(_GEN_173); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_175 = 9'ha1 == logLookUpAddr ? $signed(10'shca) : $signed(_GEN_174); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_176 = 9'ha2 == logLookUpAddr ? $signed(10'shcb) : $signed(_GEN_175); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_177 = 9'ha3 == logLookUpAddr ? $signed(10'shcc) : $signed(_GEN_176); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_178 = 9'ha4 == logLookUpAddr ? $signed(10'shcd) : $signed(_GEN_177); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_179 = 9'ha5 == logLookUpAddr ? $signed(10'shce) : $signed(_GEN_178); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_180 = 9'ha6 == logLookUpAddr ? $signed(10'shcf) : $signed(_GEN_179); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_181 = 9'ha7 == logLookUpAddr ? $signed(10'shd1) : $signed(_GEN_180); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_182 = 9'ha8 == logLookUpAddr ? $signed(10'shd2) : $signed(_GEN_181); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_183 = 9'ha9 == logLookUpAddr ? $signed(10'shd3) : $signed(_GEN_182); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_184 = 9'haa == logLookUpAddr ? $signed(10'shd4) : $signed(_GEN_183); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_185 = 9'hab == logLookUpAddr ? $signed(10'shd5) : $signed(_GEN_184); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_186 = 9'hac == logLookUpAddr ? $signed(10'shd6) : $signed(_GEN_185); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_187 = 9'had == logLookUpAddr ? $signed(10'shd7) : $signed(_GEN_186); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_188 = 9'hae == logLookUpAddr ? $signed(10'shd8) : $signed(_GEN_187); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_189 = 9'haf == logLookUpAddr ? $signed(10'shd9) : $signed(_GEN_188); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_190 = 9'hb0 == logLookUpAddr ? $signed(10'shda) : $signed(_GEN_189); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_191 = 9'hb1 == logLookUpAddr ? $signed(10'shdb) : $signed(_GEN_190); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_192 = 9'hb2 == logLookUpAddr ? $signed(10'shdc) : $signed(_GEN_191); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_193 = 9'hb3 == logLookUpAddr ? $signed(10'shdd) : $signed(_GEN_192); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_194 = 9'hb4 == logLookUpAddr ? $signed(10'shdf) : $signed(_GEN_193); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_195 = 9'hb5 == logLookUpAddr ? $signed(10'she0) : $signed(_GEN_194); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_196 = 9'hb6 == logLookUpAddr ? $signed(10'she1) : $signed(_GEN_195); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_197 = 9'hb7 == logLookUpAddr ? $signed(10'she2) : $signed(_GEN_196); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_198 = 9'hb8 == logLookUpAddr ? $signed(10'she3) : $signed(_GEN_197); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_199 = 9'hb9 == logLookUpAddr ? $signed(10'she4) : $signed(_GEN_198); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_200 = 9'hba == logLookUpAddr ? $signed(10'she5) : $signed(_GEN_199); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_201 = 9'hbb == logLookUpAddr ? $signed(10'she6) : $signed(_GEN_200); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_202 = 9'hbc == logLookUpAddr ? $signed(10'she7) : $signed(_GEN_201); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_203 = 9'hbd == logLookUpAddr ? $signed(10'she8) : $signed(_GEN_202); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_204 = 9'hbe == logLookUpAddr ? $signed(10'she9) : $signed(_GEN_203); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_205 = 9'hbf == logLookUpAddr ? $signed(10'shea) : $signed(_GEN_204); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_206 = 9'hc0 == logLookUpAddr ? $signed(10'sheb) : $signed(_GEN_205); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_207 = 9'hc1 == logLookUpAddr ? $signed(10'shec) : $signed(_GEN_206); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_208 = 9'hc2 == logLookUpAddr ? $signed(10'shed) : $signed(_GEN_207); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_209 = 9'hc3 == logLookUpAddr ? $signed(10'shee) : $signed(_GEN_208); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_210 = 9'hc4 == logLookUpAddr ? $signed(10'shef) : $signed(_GEN_209); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_211 = 9'hc5 == logLookUpAddr ? $signed(10'shf0) : $signed(_GEN_210); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_212 = 9'hc6 == logLookUpAddr ? $signed(10'shf1) : $signed(_GEN_211); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_213 = 9'hc7 == logLookUpAddr ? $signed(10'shf3) : $signed(_GEN_212); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_214 = 9'hc8 == logLookUpAddr ? $signed(10'shf4) : $signed(_GEN_213); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_215 = 9'hc9 == logLookUpAddr ? $signed(10'shf5) : $signed(_GEN_214); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_216 = 9'hca == logLookUpAddr ? $signed(10'shf6) : $signed(_GEN_215); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_217 = 9'hcb == logLookUpAddr ? $signed(10'shf7) : $signed(_GEN_216); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_218 = 9'hcc == logLookUpAddr ? $signed(10'shf8) : $signed(_GEN_217); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_219 = 9'hcd == logLookUpAddr ? $signed(10'shf9) : $signed(_GEN_218); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_220 = 9'hce == logLookUpAddr ? $signed(10'shfa) : $signed(_GEN_219); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_221 = 9'hcf == logLookUpAddr ? $signed(10'shfb) : $signed(_GEN_220); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_222 = 9'hd0 == logLookUpAddr ? $signed(10'shfc) : $signed(_GEN_221); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_223 = 9'hd1 == logLookUpAddr ? $signed(10'shfd) : $signed(_GEN_222); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_224 = 9'hd2 == logLookUpAddr ? $signed(10'shfe) : $signed(_GEN_223); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_225 = 9'hd3 == logLookUpAddr ? $signed(10'shff) : $signed(_GEN_224); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_226 = 9'hd4 == logLookUpAddr ? $signed(10'sh100) : $signed(_GEN_225); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_227 = 9'hd5 == logLookUpAddr ? $signed(10'sh101) : $signed(_GEN_226); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_228 = 9'hd6 == logLookUpAddr ? $signed(10'sh102) : $signed(_GEN_227); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_229 = 9'hd7 == logLookUpAddr ? $signed(10'sh103) : $signed(_GEN_228); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_230 = 9'hd8 == logLookUpAddr ? $signed(10'sh104) : $signed(_GEN_229); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_231 = 9'hd9 == logLookUpAddr ? $signed(10'sh105) : $signed(_GEN_230); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_232 = 9'hda == logLookUpAddr ? $signed(10'sh106) : $signed(_GEN_231); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_233 = 9'hdb == logLookUpAddr ? $signed(10'sh107) : $signed(_GEN_232); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_234 = 9'hdc == logLookUpAddr ? $signed(10'sh108) : $signed(_GEN_233); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_235 = 9'hdd == logLookUpAddr ? $signed(10'sh109) : $signed(_GEN_234); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_236 = 9'hde == logLookUpAddr ? $signed(10'sh10a) : $signed(_GEN_235); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_237 = 9'hdf == logLookUpAddr ? $signed(10'sh10b) : $signed(_GEN_236); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_238 = 9'he0 == logLookUpAddr ? $signed(10'sh10c) : $signed(_GEN_237); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_239 = 9'he1 == logLookUpAddr ? $signed(10'sh10d) : $signed(_GEN_238); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_240 = 9'he2 == logLookUpAddr ? $signed(10'sh10e) : $signed(_GEN_239); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_241 = 9'he3 == logLookUpAddr ? $signed(10'sh10f) : $signed(_GEN_240); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_242 = 9'he4 == logLookUpAddr ? $signed(10'sh110) : $signed(_GEN_241); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_243 = 9'he5 == logLookUpAddr ? $signed(10'sh111) : $signed(_GEN_242); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_244 = 9'he6 == logLookUpAddr ? $signed(10'sh112) : $signed(_GEN_243); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_245 = 9'he7 == logLookUpAddr ? $signed(10'sh113) : $signed(_GEN_244); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_246 = 9'he8 == logLookUpAddr ? $signed(10'sh114) : $signed(_GEN_245); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_247 = 9'he9 == logLookUpAddr ? $signed(10'sh115) : $signed(_GEN_246); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_248 = 9'hea == logLookUpAddr ? $signed(10'sh116) : $signed(_GEN_247); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_249 = 9'heb == logLookUpAddr ? $signed(10'sh117) : $signed(_GEN_248); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_250 = 9'hec == logLookUpAddr ? $signed(10'sh118) : $signed(_GEN_249); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_251 = 9'hed == logLookUpAddr ? $signed(10'sh119) : $signed(_GEN_250); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_252 = 9'hee == logLookUpAddr ? $signed(10'sh11a) : $signed(_GEN_251); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_253 = 9'hef == logLookUpAddr ? $signed(10'sh11b) : $signed(_GEN_252); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_254 = 9'hf0 == logLookUpAddr ? $signed(10'sh11c) : $signed(_GEN_253); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_255 = 9'hf1 == logLookUpAddr ? $signed(10'sh11d) : $signed(_GEN_254); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_256 = 9'hf2 == logLookUpAddr ? $signed(10'sh11e) : $signed(_GEN_255); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_257 = 9'hf3 == logLookUpAddr ? $signed(10'sh11f) : $signed(_GEN_256); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_258 = 9'hf4 == logLookUpAddr ? $signed(10'sh120) : $signed(_GEN_257); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_259 = 9'hf5 == logLookUpAddr ? $signed(10'sh121) : $signed(_GEN_258); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_260 = 9'hf6 == logLookUpAddr ? $signed(10'sh122) : $signed(_GEN_259); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_261 = 9'hf7 == logLookUpAddr ? $signed(10'sh123) : $signed(_GEN_260); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_262 = 9'hf8 == logLookUpAddr ? $signed(10'sh124) : $signed(_GEN_261); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_263 = 9'hf9 == logLookUpAddr ? $signed(10'sh125) : $signed(_GEN_262); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_264 = 9'hfa == logLookUpAddr ? $signed(10'sh126) : $signed(_GEN_263); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_265 = 9'hfb == logLookUpAddr ? $signed(10'sh127) : $signed(_GEN_264); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_266 = 9'hfc == logLookUpAddr ? $signed(10'sh128) : $signed(_GEN_265); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_267 = 9'hfd == logLookUpAddr ? $signed(10'sh129) : $signed(_GEN_266); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_268 = 9'hfe == logLookUpAddr ? $signed(10'sh12a) : $signed(_GEN_267); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_269 = 9'hff == logLookUpAddr ? $signed(10'sh12b) : $signed(_GEN_268); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_270 = 9'h100 == logLookUpAddr ? $signed(10'sh12c) : $signed(_GEN_269); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_271 = 9'h101 == logLookUpAddr ? $signed(10'sh12c) : $signed(_GEN_270); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_272 = 9'h102 == logLookUpAddr ? $signed(10'sh12d) : $signed(_GEN_271); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_273 = 9'h103 == logLookUpAddr ? $signed(10'sh12e) : $signed(_GEN_272); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_274 = 9'h104 == logLookUpAddr ? $signed(10'sh12f) : $signed(_GEN_273); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_275 = 9'h105 == logLookUpAddr ? $signed(10'sh130) : $signed(_GEN_274); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_276 = 9'h106 == logLookUpAddr ? $signed(10'sh131) : $signed(_GEN_275); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_277 = 9'h107 == logLookUpAddr ? $signed(10'sh132) : $signed(_GEN_276); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_278 = 9'h108 == logLookUpAddr ? $signed(10'sh133) : $signed(_GEN_277); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_279 = 9'h109 == logLookUpAddr ? $signed(10'sh134) : $signed(_GEN_278); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_280 = 9'h10a == logLookUpAddr ? $signed(10'sh135) : $signed(_GEN_279); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_281 = 9'h10b == logLookUpAddr ? $signed(10'sh136) : $signed(_GEN_280); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_282 = 9'h10c == logLookUpAddr ? $signed(10'sh137) : $signed(_GEN_281); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_283 = 9'h10d == logLookUpAddr ? $signed(10'sh138) : $signed(_GEN_282); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_284 = 9'h10e == logLookUpAddr ? $signed(10'sh139) : $signed(_GEN_283); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_285 = 9'h10f == logLookUpAddr ? $signed(10'sh13a) : $signed(_GEN_284); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_286 = 9'h110 == logLookUpAddr ? $signed(10'sh13b) : $signed(_GEN_285); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_287 = 9'h111 == logLookUpAddr ? $signed(10'sh13c) : $signed(_GEN_286); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_288 = 9'h112 == logLookUpAddr ? $signed(10'sh13d) : $signed(_GEN_287); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_289 = 9'h113 == logLookUpAddr ? $signed(10'sh13e) : $signed(_GEN_288); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_290 = 9'h114 == logLookUpAddr ? $signed(10'sh13e) : $signed(_GEN_289); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_291 = 9'h115 == logLookUpAddr ? $signed(10'sh13f) : $signed(_GEN_290); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_292 = 9'h116 == logLookUpAddr ? $signed(10'sh140) : $signed(_GEN_291); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_293 = 9'h117 == logLookUpAddr ? $signed(10'sh141) : $signed(_GEN_292); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_294 = 9'h118 == logLookUpAddr ? $signed(10'sh142) : $signed(_GEN_293); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_295 = 9'h119 == logLookUpAddr ? $signed(10'sh143) : $signed(_GEN_294); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_296 = 9'h11a == logLookUpAddr ? $signed(10'sh144) : $signed(_GEN_295); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_297 = 9'h11b == logLookUpAddr ? $signed(10'sh145) : $signed(_GEN_296); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_298 = 9'h11c == logLookUpAddr ? $signed(10'sh146) : $signed(_GEN_297); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_299 = 9'h11d == logLookUpAddr ? $signed(10'sh147) : $signed(_GEN_298); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_300 = 9'h11e == logLookUpAddr ? $signed(10'sh148) : $signed(_GEN_299); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_301 = 9'h11f == logLookUpAddr ? $signed(10'sh149) : $signed(_GEN_300); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_302 = 9'h120 == logLookUpAddr ? $signed(10'sh14a) : $signed(_GEN_301); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_303 = 9'h121 == logLookUpAddr ? $signed(10'sh14b) : $signed(_GEN_302); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_304 = 9'h122 == logLookUpAddr ? $signed(10'sh14b) : $signed(_GEN_303); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_305 = 9'h123 == logLookUpAddr ? $signed(10'sh14c) : $signed(_GEN_304); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_306 = 9'h124 == logLookUpAddr ? $signed(10'sh14d) : $signed(_GEN_305); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_307 = 9'h125 == logLookUpAddr ? $signed(10'sh14e) : $signed(_GEN_306); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_308 = 9'h126 == logLookUpAddr ? $signed(10'sh14f) : $signed(_GEN_307); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_309 = 9'h127 == logLookUpAddr ? $signed(10'sh150) : $signed(_GEN_308); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_310 = 9'h128 == logLookUpAddr ? $signed(10'sh151) : $signed(_GEN_309); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_311 = 9'h129 == logLookUpAddr ? $signed(10'sh152) : $signed(_GEN_310); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_312 = 9'h12a == logLookUpAddr ? $signed(10'sh153) : $signed(_GEN_311); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_313 = 9'h12b == logLookUpAddr ? $signed(10'sh154) : $signed(_GEN_312); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_314 = 9'h12c == logLookUpAddr ? $signed(10'sh155) : $signed(_GEN_313); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_315 = 9'h12d == logLookUpAddr ? $signed(10'sh156) : $signed(_GEN_314); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_316 = 9'h12e == logLookUpAddr ? $signed(10'sh156) : $signed(_GEN_315); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_317 = 9'h12f == logLookUpAddr ? $signed(10'sh157) : $signed(_GEN_316); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_318 = 9'h130 == logLookUpAddr ? $signed(10'sh158) : $signed(_GEN_317); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_319 = 9'h131 == logLookUpAddr ? $signed(10'sh159) : $signed(_GEN_318); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_320 = 9'h132 == logLookUpAddr ? $signed(10'sh15a) : $signed(_GEN_319); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_321 = 9'h133 == logLookUpAddr ? $signed(10'sh15b) : $signed(_GEN_320); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_322 = 9'h134 == logLookUpAddr ? $signed(10'sh15c) : $signed(_GEN_321); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_323 = 9'h135 == logLookUpAddr ? $signed(10'sh15d) : $signed(_GEN_322); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_324 = 9'h136 == logLookUpAddr ? $signed(10'sh15e) : $signed(_GEN_323); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_325 = 9'h137 == logLookUpAddr ? $signed(10'sh15f) : $signed(_GEN_324); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_326 = 9'h138 == logLookUpAddr ? $signed(10'sh15f) : $signed(_GEN_325); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_327 = 9'h139 == logLookUpAddr ? $signed(10'sh160) : $signed(_GEN_326); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_328 = 9'h13a == logLookUpAddr ? $signed(10'sh161) : $signed(_GEN_327); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_329 = 9'h13b == logLookUpAddr ? $signed(10'sh162) : $signed(_GEN_328); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_330 = 9'h13c == logLookUpAddr ? $signed(10'sh163) : $signed(_GEN_329); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_331 = 9'h13d == logLookUpAddr ? $signed(10'sh164) : $signed(_GEN_330); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_332 = 9'h13e == logLookUpAddr ? $signed(10'sh165) : $signed(_GEN_331); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_333 = 9'h13f == logLookUpAddr ? $signed(10'sh166) : $signed(_GEN_332); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_334 = 9'h140 == logLookUpAddr ? $signed(10'sh167) : $signed(_GEN_333); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_335 = 9'h141 == logLookUpAddr ? $signed(10'sh168) : $signed(_GEN_334); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_336 = 9'h142 == logLookUpAddr ? $signed(10'sh168) : $signed(_GEN_335); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_337 = 9'h143 == logLookUpAddr ? $signed(10'sh169) : $signed(_GEN_336); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_338 = 9'h144 == logLookUpAddr ? $signed(10'sh16a) : $signed(_GEN_337); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_339 = 9'h145 == logLookUpAddr ? $signed(10'sh16b) : $signed(_GEN_338); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_340 = 9'h146 == logLookUpAddr ? $signed(10'sh16c) : $signed(_GEN_339); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_341 = 9'h147 == logLookUpAddr ? $signed(10'sh16d) : $signed(_GEN_340); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_342 = 9'h148 == logLookUpAddr ? $signed(10'sh16e) : $signed(_GEN_341); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_343 = 9'h149 == logLookUpAddr ? $signed(10'sh16f) : $signed(_GEN_342); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_344 = 9'h14a == logLookUpAddr ? $signed(10'sh16f) : $signed(_GEN_343); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_345 = 9'h14b == logLookUpAddr ? $signed(10'sh170) : $signed(_GEN_344); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_346 = 9'h14c == logLookUpAddr ? $signed(10'sh171) : $signed(_GEN_345); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_347 = 9'h14d == logLookUpAddr ? $signed(10'sh172) : $signed(_GEN_346); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_348 = 9'h14e == logLookUpAddr ? $signed(10'sh173) : $signed(_GEN_347); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_349 = 9'h14f == logLookUpAddr ? $signed(10'sh174) : $signed(_GEN_348); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_350 = 9'h150 == logLookUpAddr ? $signed(10'sh175) : $signed(_GEN_349); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_351 = 9'h151 == logLookUpAddr ? $signed(10'sh176) : $signed(_GEN_350); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_352 = 9'h152 == logLookUpAddr ? $signed(10'sh176) : $signed(_GEN_351); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_353 = 9'h153 == logLookUpAddr ? $signed(10'sh177) : $signed(_GEN_352); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_354 = 9'h154 == logLookUpAddr ? $signed(10'sh178) : $signed(_GEN_353); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_355 = 9'h155 == logLookUpAddr ? $signed(10'sh179) : $signed(_GEN_354); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_356 = 9'h156 == logLookUpAddr ? $signed(10'sh17a) : $signed(_GEN_355); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_357 = 9'h157 == logLookUpAddr ? $signed(10'sh17b) : $signed(_GEN_356); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_358 = 9'h158 == logLookUpAddr ? $signed(10'sh17c) : $signed(_GEN_357); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_359 = 9'h159 == logLookUpAddr ? $signed(10'sh17c) : $signed(_GEN_358); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_360 = 9'h15a == logLookUpAddr ? $signed(10'sh17d) : $signed(_GEN_359); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_361 = 9'h15b == logLookUpAddr ? $signed(10'sh17e) : $signed(_GEN_360); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_362 = 9'h15c == logLookUpAddr ? $signed(10'sh17f) : $signed(_GEN_361); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_363 = 9'h15d == logLookUpAddr ? $signed(10'sh180) : $signed(_GEN_362); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_364 = 9'h15e == logLookUpAddr ? $signed(10'sh181) : $signed(_GEN_363); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_365 = 9'h15f == logLookUpAddr ? $signed(10'sh182) : $signed(_GEN_364); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_366 = 9'h160 == logLookUpAddr ? $signed(10'sh183) : $signed(_GEN_365); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_367 = 9'h161 == logLookUpAddr ? $signed(10'sh183) : $signed(_GEN_366); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_368 = 9'h162 == logLookUpAddr ? $signed(10'sh184) : $signed(_GEN_367); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_369 = 9'h163 == logLookUpAddr ? $signed(10'sh185) : $signed(_GEN_368); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_370 = 9'h164 == logLookUpAddr ? $signed(10'sh186) : $signed(_GEN_369); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_371 = 9'h165 == logLookUpAddr ? $signed(10'sh187) : $signed(_GEN_370); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_372 = 9'h166 == logLookUpAddr ? $signed(10'sh188) : $signed(_GEN_371); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_373 = 9'h167 == logLookUpAddr ? $signed(10'sh188) : $signed(_GEN_372); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_374 = 9'h168 == logLookUpAddr ? $signed(10'sh189) : $signed(_GEN_373); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_375 = 9'h169 == logLookUpAddr ? $signed(10'sh18a) : $signed(_GEN_374); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_376 = 9'h16a == logLookUpAddr ? $signed(10'sh18b) : $signed(_GEN_375); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_377 = 9'h16b == logLookUpAddr ? $signed(10'sh18c) : $signed(_GEN_376); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_378 = 9'h16c == logLookUpAddr ? $signed(10'sh18d) : $signed(_GEN_377); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_379 = 9'h16d == logLookUpAddr ? $signed(10'sh18e) : $signed(_GEN_378); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_380 = 9'h16e == logLookUpAddr ? $signed(10'sh18e) : $signed(_GEN_379); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_381 = 9'h16f == logLookUpAddr ? $signed(10'sh18f) : $signed(_GEN_380); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_382 = 9'h170 == logLookUpAddr ? $signed(10'sh190) : $signed(_GEN_381); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_383 = 9'h171 == logLookUpAddr ? $signed(10'sh191) : $signed(_GEN_382); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_384 = 9'h172 == logLookUpAddr ? $signed(10'sh192) : $signed(_GEN_383); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_385 = 9'h173 == logLookUpAddr ? $signed(10'sh193) : $signed(_GEN_384); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_386 = 9'h174 == logLookUpAddr ? $signed(10'sh193) : $signed(_GEN_385); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_387 = 9'h175 == logLookUpAddr ? $signed(10'sh194) : $signed(_GEN_386); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_388 = 9'h176 == logLookUpAddr ? $signed(10'sh195) : $signed(_GEN_387); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_389 = 9'h177 == logLookUpAddr ? $signed(10'sh196) : $signed(_GEN_388); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_390 = 9'h178 == logLookUpAddr ? $signed(10'sh197) : $signed(_GEN_389); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_391 = 9'h179 == logLookUpAddr ? $signed(10'sh198) : $signed(_GEN_390); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_392 = 9'h17a == logLookUpAddr ? $signed(10'sh198) : $signed(_GEN_391); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_393 = 9'h17b == logLookUpAddr ? $signed(10'sh199) : $signed(_GEN_392); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_394 = 9'h17c == logLookUpAddr ? $signed(10'sh19a) : $signed(_GEN_393); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_395 = 9'h17d == logLookUpAddr ? $signed(10'sh19b) : $signed(_GEN_394); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_396 = 9'h17e == logLookUpAddr ? $signed(10'sh19c) : $signed(_GEN_395); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_397 = 9'h17f == logLookUpAddr ? $signed(10'sh19d) : $signed(_GEN_396); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_398 = 9'h180 == logLookUpAddr ? $signed(10'sh19d) : $signed(_GEN_397); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_399 = 9'h181 == logLookUpAddr ? $signed(10'sh19e) : $signed(_GEN_398); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_400 = 9'h182 == logLookUpAddr ? $signed(10'sh19f) : $signed(_GEN_399); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_401 = 9'h183 == logLookUpAddr ? $signed(10'sh1a0) : $signed(_GEN_400); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_402 = 9'h184 == logLookUpAddr ? $signed(10'sh1a1) : $signed(_GEN_401); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_403 = 9'h185 == logLookUpAddr ? $signed(10'sh1a1) : $signed(_GEN_402); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_404 = 9'h186 == logLookUpAddr ? $signed(10'sh1a2) : $signed(_GEN_403); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_405 = 9'h187 == logLookUpAddr ? $signed(10'sh1a3) : $signed(_GEN_404); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_406 = 9'h188 == logLookUpAddr ? $signed(10'sh1a4) : $signed(_GEN_405); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_407 = 9'h189 == logLookUpAddr ? $signed(10'sh1a5) : $signed(_GEN_406); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_408 = 9'h18a == logLookUpAddr ? $signed(10'sh1a6) : $signed(_GEN_407); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_409 = 9'h18b == logLookUpAddr ? $signed(10'sh1a6) : $signed(_GEN_408); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_410 = 9'h18c == logLookUpAddr ? $signed(10'sh1a7) : $signed(_GEN_409); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_411 = 9'h18d == logLookUpAddr ? $signed(10'sh1a8) : $signed(_GEN_410); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_412 = 9'h18e == logLookUpAddr ? $signed(10'sh1a9) : $signed(_GEN_411); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_413 = 9'h18f == logLookUpAddr ? $signed(10'sh1aa) : $signed(_GEN_412); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_414 = 9'h190 == logLookUpAddr ? $signed(10'sh1aa) : $signed(_GEN_413); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_415 = 9'h191 == logLookUpAddr ? $signed(10'sh1ab) : $signed(_GEN_414); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_416 = 9'h192 == logLookUpAddr ? $signed(10'sh1ac) : $signed(_GEN_415); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_417 = 9'h193 == logLookUpAddr ? $signed(10'sh1ad) : $signed(_GEN_416); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_418 = 9'h194 == logLookUpAddr ? $signed(10'sh1ae) : $signed(_GEN_417); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_419 = 9'h195 == logLookUpAddr ? $signed(10'sh1ae) : $signed(_GEN_418); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_420 = 9'h196 == logLookUpAddr ? $signed(10'sh1af) : $signed(_GEN_419); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_421 = 9'h197 == logLookUpAddr ? $signed(10'sh1b0) : $signed(_GEN_420); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_422 = 9'h198 == logLookUpAddr ? $signed(10'sh1b1) : $signed(_GEN_421); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_423 = 9'h199 == logLookUpAddr ? $signed(10'sh1b2) : $signed(_GEN_422); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_424 = 9'h19a == logLookUpAddr ? $signed(10'sh1b2) : $signed(_GEN_423); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_425 = 9'h19b == logLookUpAddr ? $signed(10'sh1b3) : $signed(_GEN_424); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_426 = 9'h19c == logLookUpAddr ? $signed(10'sh1b4) : $signed(_GEN_425); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_427 = 9'h19d == logLookUpAddr ? $signed(10'sh1b5) : $signed(_GEN_426); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_428 = 9'h19e == logLookUpAddr ? $signed(10'sh1b6) : $signed(_GEN_427); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_429 = 9'h19f == logLookUpAddr ? $signed(10'sh1b6) : $signed(_GEN_428); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_430 = 9'h1a0 == logLookUpAddr ? $signed(10'sh1b7) : $signed(_GEN_429); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_431 = 9'h1a1 == logLookUpAddr ? $signed(10'sh1b8) : $signed(_GEN_430); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_432 = 9'h1a2 == logLookUpAddr ? $signed(10'sh1b9) : $signed(_GEN_431); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_433 = 9'h1a3 == logLookUpAddr ? $signed(10'sh1ba) : $signed(_GEN_432); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_434 = 9'h1a4 == logLookUpAddr ? $signed(10'sh1ba) : $signed(_GEN_433); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_435 = 9'h1a5 == logLookUpAddr ? $signed(10'sh1bb) : $signed(_GEN_434); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_436 = 9'h1a6 == logLookUpAddr ? $signed(10'sh1bc) : $signed(_GEN_435); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_437 = 9'h1a7 == logLookUpAddr ? $signed(10'sh1bd) : $signed(_GEN_436); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_438 = 9'h1a8 == logLookUpAddr ? $signed(10'sh1be) : $signed(_GEN_437); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_439 = 9'h1a9 == logLookUpAddr ? $signed(10'sh1be) : $signed(_GEN_438); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_440 = 9'h1aa == logLookUpAddr ? $signed(10'sh1bf) : $signed(_GEN_439); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_441 = 9'h1ab == logLookUpAddr ? $signed(10'sh1c0) : $signed(_GEN_440); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_442 = 9'h1ac == logLookUpAddr ? $signed(10'sh1c1) : $signed(_GEN_441); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_443 = 9'h1ad == logLookUpAddr ? $signed(10'sh1c2) : $signed(_GEN_442); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_444 = 9'h1ae == logLookUpAddr ? $signed(10'sh1c2) : $signed(_GEN_443); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_445 = 9'h1af == logLookUpAddr ? $signed(10'sh1c3) : $signed(_GEN_444); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_446 = 9'h1b0 == logLookUpAddr ? $signed(10'sh1c4) : $signed(_GEN_445); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_447 = 9'h1b1 == logLookUpAddr ? $signed(10'sh1c5) : $signed(_GEN_446); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_448 = 9'h1b2 == logLookUpAddr ? $signed(10'sh1c5) : $signed(_GEN_447); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_449 = 9'h1b3 == logLookUpAddr ? $signed(10'sh1c6) : $signed(_GEN_448); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_450 = 9'h1b4 == logLookUpAddr ? $signed(10'sh1c7) : $signed(_GEN_449); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_451 = 9'h1b5 == logLookUpAddr ? $signed(10'sh1c8) : $signed(_GEN_450); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_452 = 9'h1b6 == logLookUpAddr ? $signed(10'sh1c9) : $signed(_GEN_451); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_453 = 9'h1b7 == logLookUpAddr ? $signed(10'sh1c9) : $signed(_GEN_452); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_454 = 9'h1b8 == logLookUpAddr ? $signed(10'sh1ca) : $signed(_GEN_453); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_455 = 9'h1b9 == logLookUpAddr ? $signed(10'sh1cb) : $signed(_GEN_454); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_456 = 9'h1ba == logLookUpAddr ? $signed(10'sh1cc) : $signed(_GEN_455); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_457 = 9'h1bb == logLookUpAddr ? $signed(10'sh1cc) : $signed(_GEN_456); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_458 = 9'h1bc == logLookUpAddr ? $signed(10'sh1cd) : $signed(_GEN_457); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_459 = 9'h1bd == logLookUpAddr ? $signed(10'sh1ce) : $signed(_GEN_458); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_460 = 9'h1be == logLookUpAddr ? $signed(10'sh1cf) : $signed(_GEN_459); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_461 = 9'h1bf == logLookUpAddr ? $signed(10'sh1d0) : $signed(_GEN_460); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_462 = 9'h1c0 == logLookUpAddr ? $signed(10'sh1d0) : $signed(_GEN_461); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_463 = 9'h1c1 == logLookUpAddr ? $signed(10'sh1d1) : $signed(_GEN_462); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_464 = 9'h1c2 == logLookUpAddr ? $signed(10'sh1d2) : $signed(_GEN_463); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_465 = 9'h1c3 == logLookUpAddr ? $signed(10'sh1d3) : $signed(_GEN_464); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_466 = 9'h1c4 == logLookUpAddr ? $signed(10'sh1d3) : $signed(_GEN_465); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_467 = 9'h1c5 == logLookUpAddr ? $signed(10'sh1d4) : $signed(_GEN_466); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_468 = 9'h1c6 == logLookUpAddr ? $signed(10'sh1d5) : $signed(_GEN_467); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_469 = 9'h1c7 == logLookUpAddr ? $signed(10'sh1d6) : $signed(_GEN_468); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_470 = 9'h1c8 == logLookUpAddr ? $signed(10'sh1d6) : $signed(_GEN_469); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_471 = 9'h1c9 == logLookUpAddr ? $signed(10'sh1d7) : $signed(_GEN_470); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_472 = 9'h1ca == logLookUpAddr ? $signed(10'sh1d8) : $signed(_GEN_471); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_473 = 9'h1cb == logLookUpAddr ? $signed(10'sh1d9) : $signed(_GEN_472); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_474 = 9'h1cc == logLookUpAddr ? $signed(10'sh1da) : $signed(_GEN_473); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_475 = 9'h1cd == logLookUpAddr ? $signed(10'sh1da) : $signed(_GEN_474); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_476 = 9'h1ce == logLookUpAddr ? $signed(10'sh1db) : $signed(_GEN_475); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_477 = 9'h1cf == logLookUpAddr ? $signed(10'sh1dc) : $signed(_GEN_476); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_478 = 9'h1d0 == logLookUpAddr ? $signed(10'sh1dd) : $signed(_GEN_477); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_479 = 9'h1d1 == logLookUpAddr ? $signed(10'sh1dd) : $signed(_GEN_478); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_480 = 9'h1d2 == logLookUpAddr ? $signed(10'sh1de) : $signed(_GEN_479); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_481 = 9'h1d3 == logLookUpAddr ? $signed(10'sh1df) : $signed(_GEN_480); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_482 = 9'h1d4 == logLookUpAddr ? $signed(10'sh1e0) : $signed(_GEN_481); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_483 = 9'h1d5 == logLookUpAddr ? $signed(10'sh1e0) : $signed(_GEN_482); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_484 = 9'h1d6 == logLookUpAddr ? $signed(10'sh1e1) : $signed(_GEN_483); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_485 = 9'h1d7 == logLookUpAddr ? $signed(10'sh1e2) : $signed(_GEN_484); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_486 = 9'h1d8 == logLookUpAddr ? $signed(10'sh1e3) : $signed(_GEN_485); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_487 = 9'h1d9 == logLookUpAddr ? $signed(10'sh1e3) : $signed(_GEN_486); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_488 = 9'h1da == logLookUpAddr ? $signed(10'sh1e4) : $signed(_GEN_487); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_489 = 9'h1db == logLookUpAddr ? $signed(10'sh1e5) : $signed(_GEN_488); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_490 = 9'h1dc == logLookUpAddr ? $signed(10'sh1e6) : $signed(_GEN_489); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_491 = 9'h1dd == logLookUpAddr ? $signed(10'sh1e6) : $signed(_GEN_490); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_492 = 9'h1de == logLookUpAddr ? $signed(10'sh1e7) : $signed(_GEN_491); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_493 = 9'h1df == logLookUpAddr ? $signed(10'sh1e8) : $signed(_GEN_492); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_494 = 9'h1e0 == logLookUpAddr ? $signed(10'sh1e9) : $signed(_GEN_493); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_495 = 9'h1e1 == logLookUpAddr ? $signed(10'sh1e9) : $signed(_GEN_494); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_496 = 9'h1e2 == logLookUpAddr ? $signed(10'sh1ea) : $signed(_GEN_495); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_497 = 9'h1e3 == logLookUpAddr ? $signed(10'sh1eb) : $signed(_GEN_496); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_498 = 9'h1e4 == logLookUpAddr ? $signed(10'sh1ec) : $signed(_GEN_497); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_499 = 9'h1e5 == logLookUpAddr ? $signed(10'sh1ec) : $signed(_GEN_498); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_500 = 9'h1e6 == logLookUpAddr ? $signed(10'sh1ed) : $signed(_GEN_499); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_501 = 9'h1e7 == logLookUpAddr ? $signed(10'sh1ee) : $signed(_GEN_500); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_502 = 9'h1e8 == logLookUpAddr ? $signed(10'sh1ee) : $signed(_GEN_501); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_503 = 9'h1e9 == logLookUpAddr ? $signed(10'sh1ef) : $signed(_GEN_502); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_504 = 9'h1ea == logLookUpAddr ? $signed(10'sh1f0) : $signed(_GEN_503); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_505 = 9'h1eb == logLookUpAddr ? $signed(10'sh1f1) : $signed(_GEN_504); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_506 = 9'h1ec == logLookUpAddr ? $signed(10'sh1f1) : $signed(_GEN_505); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_507 = 9'h1ed == logLookUpAddr ? $signed(10'sh1f2) : $signed(_GEN_506); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_508 = 9'h1ee == logLookUpAddr ? $signed(10'sh1f3) : $signed(_GEN_507); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_509 = 9'h1ef == logLookUpAddr ? $signed(10'sh1f4) : $signed(_GEN_508); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_510 = 9'h1f0 == logLookUpAddr ? $signed(10'sh1f4) : $signed(_GEN_509); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_511 = 9'h1f1 == logLookUpAddr ? $signed(10'sh1f5) : $signed(_GEN_510); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_512 = 9'h1f2 == logLookUpAddr ? $signed(10'sh1f6) : $signed(_GEN_511); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_513 = 9'h1f3 == logLookUpAddr ? $signed(10'sh1f7) : $signed(_GEN_512); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_514 = 9'h1f4 == logLookUpAddr ? $signed(10'sh1f7) : $signed(_GEN_513); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_515 = 9'h1f5 == logLookUpAddr ? $signed(10'sh1f8) : $signed(_GEN_514); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_516 = 9'h1f6 == logLookUpAddr ? $signed(10'sh1f9) : $signed(_GEN_515); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_517 = 9'h1f7 == logLookUpAddr ? $signed(10'sh1f9) : $signed(_GEN_516); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_518 = 9'h1f8 == logLookUpAddr ? $signed(10'sh1fa) : $signed(_GEN_517); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_519 = 9'h1f9 == logLookUpAddr ? $signed(10'sh1fb) : $signed(_GEN_518); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_520 = 9'h1fa == logLookUpAddr ? $signed(10'sh1fc) : $signed(_GEN_519); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_521 = 9'h1fb == logLookUpAddr ? $signed(10'sh1fc) : $signed(_GEN_520); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_522 = 9'h1fc == logLookUpAddr ? $signed(10'sh1fd) : $signed(_GEN_521); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_523 = 9'h1fd == logLookUpAddr ? $signed(10'sh1fe) : $signed(_GEN_522); // @[LogMagMux.scala 136:11]
  wire [9:0] _GEN_524 = 9'h1fe == logLookUpAddr ? $signed(10'sh1ff) : $signed(_GEN_523); // @[LogMagMux.scala 136:11]
  wire [9:0] logFrac = 9'h1ff == logLookUpAddr ? $signed(10'sh1ff) : $signed(_GEN_524); // @[LogMagMux.scala 136:11]
  reg [4:0] _T_601; // @[Reg.scala 15:16]
  reg [31:0] _RAND_14;
  wire [13:0] _GEN_564 = {$signed(_T_601), 9'h0}; // @[LogMagMux.scala 141:91]
  wire [13:0] _GEN_565 = {{4{logFrac[9]}},logFrac}; // @[LogMagMux.scala 141:91]
  wire [13:0] _T_604 = $signed(_GEN_564) + $signed(_GEN_565); // @[LogMagMux.scala 141:91]
  wire [15:0] log2MagOut_imag = {{2{_T_604[13]}},_T_604}; // @[LogMagMux.scala 160:38]
  reg [1:0] _T_614; // @[Reg.scala 15:16]
  reg [31:0] _RAND_15;
  reg [1:0] _T_615; // @[Reg.scala 15:16]
  reg [31:0] _RAND_16;
  reg [1:0] _T_616; // @[Reg.scala 15:16]
  reg [31:0] _RAND_17;
  reg [1:0] _T_617; // @[Reg.scala 15:16]
  reg [31:0] _RAND_18;
  reg [15:0] _T_620_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_19;
  reg [15:0] _T_620_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_20;
  reg [15:0] _T_623_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_21;
  reg [15:0] _T_623_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_22;
  reg [15:0] _T_626_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_23;
  reg [15:0] _T_626_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_24;
  reg [15:0] _T_629_real; // @[Reg.scala 15:16]
  reg [31:0] _RAND_25;
  reg [15:0] _T_629_imag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_26;
  wire  _T_630 = 2'h3 == _T_617; // @[Mux.scala 68:19]
  wire [15:0] _T_633_real = _T_630 ? $signed(16'sh0) : $signed(io_in_bits_real); // @[Mux.scala 68:16]
  wire [15:0] _T_633_imag = _T_630 ? $signed(log2MagOut_imag) : $signed(io_in_bits_imag); // @[Mux.scala 68:16]
  wire  _T_634 = 2'h2 == _T_617; // @[Mux.scala 68:19]
  wire [15:0] _T_637_real = _T_634 ? $signed(16'sh0) : $signed(_T_633_real); // @[Mux.scala 68:16]
  wire [15:0] jplMagOut_imag = jplMag[15:0]; // @[LogMagMux.scala 151:23 LogMagMux.scala 154:18]
  wire [15:0] _T_637_imag = _T_634 ? $signed(jplMagOut_imag) : $signed(_T_633_imag); // @[Mux.scala 68:16]
  wire  _T_638 = 2'h1 == _T_617; // @[Mux.scala 68:19]
  wire [15:0] _T_641_real = _T_638 ? $signed(16'sh0) : $signed(_T_637_real); // @[Mux.scala 68:16]
  wire [32:0] _GEN_567 = _T_31[33:1]; // @[LogMagMux.scala 95:20 LogMagMux.scala 105:10]
  wire [15:0] magSqr = _GEN_567[15:0]; // @[LogMagMux.scala 95:20 LogMagMux.scala 105:10]
  wire [15:0] _T_641_imag = _T_638 ? $signed(magSqr) : $signed(_T_637_imag); // @[Mux.scala 68:16]
  wire  _T_642 = 2'h0 == _T_617; // @[Mux.scala 68:19]
  wire [15:0] output_mux_real = _T_642 ? $signed(_T_629_real) : $signed(_T_641_real); // @[Mux.scala 68:16]
  wire [15:0] output_mux_imag = _T_642 ? $signed(_T_629_imag) : $signed(_T_641_imag); // @[Mux.scala 68:16]
  wire  _T_645 = io_in_ready & io_in_valid; // @[Decoupled.scala 40:37]
  reg  initialInDone; // @[LogMagMux.scala 187:30]
  reg [31:0] _RAND_27;
  reg [2:0] _T_653; // @[LogMagMux.scala 190:24]
  reg [31:0] _RAND_28;
  wire [2:0] _T_656 = _T_653 + 3'h1; // @[LogMagMux.scala 193:22]
  wire  _T_657 = _T_653 == 3'h3; // @[LogMagMux.scala 196:18]
  wire  _T_659 = _T_657 & _T_645; // @[LogMagMux.scala 196:39]
  wire  _GEN_544 = _T_659 | initialInDone; // @[LogMagMux.scala 196:56]
  wire  _T_667 = ~initialInDone; // @[Skid.scala 29:30]
  wire  _T_668 = io_out_ready | _T_667; // @[Skid.scala 29:27]
  wire  skidInData_ready = _T_668; // @[LogMagMux.scala 205:24 Skid.scala 29:14]
  wire  skidInData_valid = io_in_valid; // @[LogMagMux.scala 205:24 LogMagMux.scala 207:20]
  wire  _T_662 = skidInData_ready & skidInData_valid; // @[Decoupled.scala 40:37]
  reg  _T_663; // @[Reg.scala 27:20]
  reg [31:0] _RAND_29;
  reg  _T_664; // @[Reg.scala 27:20]
  reg [31:0] _RAND_30;
  reg  _T_665; // @[Reg.scala 27:20]
  reg [31:0] _RAND_31;
  reg  _T_666; // @[Reg.scala 27:20]
  reg [31:0] _RAND_32;
  reg  _T_673; // @[Reg.scala 15:16]
  reg [31:0] _RAND_33;
  reg  _T_674; // @[Reg.scala 15:16]
  reg [31:0] _RAND_34;
  reg  _T_675; // @[Reg.scala 15:16]
  reg [31:0] _RAND_35;
  reg  _T_676; // @[Reg.scala 15:16]
  reg [31:0] _RAND_36;
  wire  _T_677 = _T_668 & io_in_valid; // @[Decoupled.scala 40:37]
  reg  _T_678; // @[Reg.scala 27:20]
  reg [31:0] _RAND_37;
  reg  _T_679; // @[Reg.scala 27:20]
  reg [31:0] _RAND_38;
  reg  _T_680; // @[Reg.scala 27:20]
  reg [31:0] _RAND_39;
  reg  _T_681; // @[Reg.scala 27:20]
  reg [31:0] _RAND_40;
  wire [15:0] skidInData_bits_real = output_mux_real; // @[LogMagMux.scala 205:24 LogMagMux.scala 206:19]
  wire [15:0] skidInData_bits_imag = output_mux_imag; // @[LogMagMux.scala 205:24 LogMagMux.scala 206:19]
  Queue_15 Queue ( // @[Skid.scala 21:23]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_real(Queue_io_enq_bits_real),
    .io_enq_bits_imag(Queue_io_enq_bits_imag),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_real(Queue_io_deq_bits_real),
    .io_deq_bits_imag(Queue_io_deq_bits_imag)
  );
  Queue_16 Queue_1 ( // @[Skid.scala 21:23]
    .clock(Queue_1_clock),
    .reset(Queue_1_reset),
    .io_enq_ready(Queue_1_io_enq_ready),
    .io_enq_valid(Queue_1_io_enq_valid),
    .io_enq_bits(Queue_1_io_enq_bits),
    .io_deq_ready(Queue_1_io_deq_ready),
    .io_deq_valid(Queue_1_io_deq_valid),
    .io_deq_bits(Queue_1_io_deq_bits)
  );
  assign io_in_ready = skidInData_ready; // @[LogMagMux.scala 210:15]
  assign io_out_valid = Queue_io_deq_valid; // @[Skid.scala 31:15]
  assign io_out_bits_real = Queue_io_deq_bits_real; // @[Skid.scala 32:14]
  assign io_out_bits_imag = Queue_io_deq_bits_imag; // @[Skid.scala 32:14]
  assign io_lastOut = Queue_1_io_deq_bits; // @[LogMagMux.scala 220:20]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = _T_666; // @[Skid.scala 25:24]
  assign Queue_io_enq_bits_real = output_mux_real; // @[LogMagMux.scala 211:52]
  assign Queue_io_enq_bits_imag = output_mux_imag; // @[LogMagMux.scala 211:52]
  assign Queue_io_deq_ready = io_out_ready; // @[Skid.scala 30:24]
  assign Queue_1_clock = clock;
  assign Queue_1_reset = reset;
  assign Queue_1_io_enq_valid = _T_681; // @[Skid.scala 25:24]
  assign Queue_1_io_enq_bits = _T_676; // @[LogMagMux.scala 219:59]
  assign Queue_1_io_deq_ready = io_out_ready; // @[Skid.scala 30:24]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_16 = _RAND_0[16:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  jplMagOp1 = _RAND_1[16:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  tmpOp2 = _RAND_2[16:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_20 = _RAND_3[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  jplMagOp2 = _RAND_4[17:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_23 = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_26 = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {2{`RANDOM}};
  _T_29 = _RAND_7[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {2{`RANDOM}};
  _T_30 = _RAND_8[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {2{`RANDOM}};
  _T_31 = _RAND_9[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_33 = _RAND_10[17:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  jplMag = _RAND_11[17:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  noLeadOne = _RAND_12[17:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  shiftNum = _RAND_13[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_601 = _RAND_14[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_614 = _RAND_15[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_615 = _RAND_16[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_616 = _RAND_17[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_617 = _RAND_18[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_620_real = _RAND_19[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_620_imag = _RAND_20[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_623_real = _RAND_21[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_623_imag = _RAND_22[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_626_real = _RAND_23[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_626_imag = _RAND_24[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_629_real = _RAND_25[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_629_imag = _RAND_26[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  initialInDone = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_653 = _RAND_28[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_663 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_664 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T_665 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _T_666 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _T_673 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _T_674 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _T_675 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _T_676 = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _T_678 = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _T_679 = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _T_680 = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _T_681 = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_16 <= $signed(u) + $signed(_GEN_559);
    jplMagOp1 <= _T_16;
    tmpOp2 <= $signed(u) - $signed(_GEN_560);
    _T_20 <= v[15:1];
    jplMagOp2 <= $signed(tmpOp2) + $signed(_GEN_561);
    _T_23 <= $signed(absInReal) * $signed(absInReal);
    _T_26 <= $signed(absInImag) * $signed(absInImag);
    _T_29 <= $signed(_T_24) + $signed(_T_27);
    _T_30 <= _T_29;
    _T_31 <= _T_30;
    if (_T_32) begin
      _T_33 <= {{1{jplMagOp1[16]}},jplMagOp1};
    end else begin
      _T_33 <= jplMagOp2;
    end
    jplMag <= _T_33;
    noLeadOne <= _T_589 - _T_590[17:0];
    shiftNum <= _T_596 - 5'h1;
    _T_601 <= logUInt - 5'h0;
    _T_614 <= io_sel;
    _T_615 <= _T_614;
    _T_616 <= _T_615;
    _T_617 <= _T_616;
    _T_620_real <= io_in_bits_real;
    _T_620_imag <= io_in_bits_imag;
    _T_623_real <= _T_620_real;
    _T_623_imag <= _T_620_imag;
    _T_626_real <= _T_623_real;
    _T_626_imag <= _T_623_imag;
    _T_629_real <= _T_626_real;
    _T_629_imag <= _T_626_imag;
    if (reset) begin
      initialInDone <= 1'h0;
    end else if (io_lastOut) begin
      initialInDone <= 1'h0;
    end else begin
      initialInDone <= _GEN_544;
    end
    if (reset) begin
      _T_653 <= 3'h0;
    end else if (io_lastOut) begin
      _T_653 <= 3'h0;
    end else if (_T_645) begin
      _T_653 <= _T_656;
    end
    if (reset) begin
      _T_663 <= 1'h0;
    end else begin
      _T_663 <= _T_662;
    end
    if (reset) begin
      _T_664 <= 1'h0;
    end else begin
      _T_664 <= _T_663;
    end
    if (reset) begin
      _T_665 <= 1'h0;
    end else begin
      _T_665 <= _T_664;
    end
    if (reset) begin
      _T_666 <= 1'h0;
    end else begin
      _T_666 <= _T_665;
    end
    _T_673 <= io_lastIn & _T_645;
    _T_674 <= _T_673;
    _T_675 <= _T_674;
    _T_676 <= _T_675;
    if (reset) begin
      _T_678 <= 1'h0;
    end else begin
      _T_678 <= _T_677;
    end
    if (reset) begin
      _T_679 <= 1'h0;
    end else begin
      _T_679 <= _T_678;
    end
    if (reset) begin
      _T_680 <= 1'h0;
    end else begin
      _T_680 <= _T_679;
    end
    if (reset) begin
      _T_681 <= 1'h0;
    end else begin
      _T_681 <= _T_680;
    end
  end
endmodule
module AXI4LogMagMuxBlock(
  input         clock,
  input         reset,
  output        auto_mem_in_aw_ready,
  input         auto_mem_in_aw_valid,
  input         auto_mem_in_aw_bits_id,
  input  [29:0] auto_mem_in_aw_bits_addr,
  output        auto_mem_in_w_ready,
  input         auto_mem_in_w_valid,
  input  [31:0] auto_mem_in_w_bits_data,
  input  [3:0]  auto_mem_in_w_bits_strb,
  input         auto_mem_in_b_ready,
  output        auto_mem_in_b_valid,
  output        auto_mem_in_b_bits_id,
  output        auto_mem_in_ar_ready,
  input         auto_mem_in_ar_valid,
  input         auto_mem_in_ar_bits_id,
  input  [29:0] auto_mem_in_ar_bits_addr,
  input  [2:0]  auto_mem_in_ar_bits_size,
  input         auto_mem_in_r_ready,
  output        auto_mem_in_r_valid,
  output        auto_mem_in_r_bits_id,
  output [31:0] auto_mem_in_r_bits_data,
  output        auto_stream_in_ready,
  input         auto_stream_in_valid,
  input  [31:0] auto_stream_in_bits_data,
  input         auto_stream_in_bits_last,
  input         auto_stream_out_ready,
  output        auto_stream_out_valid,
  output [31:0] auto_stream_out_bits_data,
  output        auto_stream_out_bits_last
);
  wire  logMagMux_clock; // @[LogMagMuxDspBlock.scala 27:27]
  wire  logMagMux_reset; // @[LogMagMuxDspBlock.scala 27:27]
  wire  logMagMux_io_in_ready; // @[LogMagMuxDspBlock.scala 27:27]
  wire  logMagMux_io_in_valid; // @[LogMagMuxDspBlock.scala 27:27]
  wire [15:0] logMagMux_io_in_bits_real; // @[LogMagMuxDspBlock.scala 27:27]
  wire [15:0] logMagMux_io_in_bits_imag; // @[LogMagMuxDspBlock.scala 27:27]
  wire  logMagMux_io_lastIn; // @[LogMagMuxDspBlock.scala 27:27]
  wire  logMagMux_io_out_ready; // @[LogMagMuxDspBlock.scala 27:27]
  wire  logMagMux_io_out_valid; // @[LogMagMuxDspBlock.scala 27:27]
  wire [15:0] logMagMux_io_out_bits_real; // @[LogMagMuxDspBlock.scala 27:27]
  wire [15:0] logMagMux_io_out_bits_imag; // @[LogMagMuxDspBlock.scala 27:27]
  wire [1:0] logMagMux_io_sel; // @[LogMagMuxDspBlock.scala 27:27]
  wire  logMagMux_io_lastOut; // @[LogMagMuxDspBlock.scala 27:27]
  wire  Queue_clock; // @[Decoupled.scala 296:21]
  wire  Queue_reset; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_bits_read; // @[Decoupled.scala 296:21]
  wire [31:0] Queue_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_bits_extra; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_bits_read; // @[Decoupled.scala 296:21]
  wire [31:0] Queue_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_bits_extra; // @[Decoupled.scala 296:21]
  reg [1:0] selReg; // @[LogMagMuxDspBlock.scala 29:33]
  reg [31:0] _RAND_0;
  wire  _T_2 = auto_mem_in_aw_valid & auto_mem_in_w_valid; // @[RegisterRouter.scala 40:39]
  wire  _T_3 = auto_mem_in_ar_valid | _T_2; // @[RegisterRouter.scala 40:26]
  wire  _T_4 = ~auto_mem_in_ar_valid; // @[RegisterRouter.scala 42:29]
  wire  _T_47_ready = Queue_io_enq_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 299:17]
  wire [29:0] _T_11 = auto_mem_in_ar_valid ? auto_mem_in_ar_bits_addr : auto_mem_in_aw_bits_addr; // @[RegisterRouter.scala 48:19]
  wire  _T_53 = _T_11[7:2] == 6'h0; // @[RegisterRouter.scala 59:16]
  wire  _T_5 = _T_47_ready & _T_4; // @[RegisterRouter.scala 42:26]
  wire [1:0] _T_14 = 2'h1 << auto_mem_in_ar_bits_size[0]; // @[OneHot.scala 65:12]
  wire [1:0] _T_16 = _T_14 | 2'h1; // @[Misc.scala 200:81]
  wire  _T_17 = auto_mem_in_ar_bits_size >= 3'h2; // @[Misc.scala 204:21]
  wire  _T_20 = ~auto_mem_in_ar_bits_addr[1]; // @[Misc.scala 209:20]
  wire  _T_22 = _T_16[1] & _T_20; // @[Misc.scala 213:38]
  wire  _T_23 = _T_17 | _T_22; // @[Misc.scala 213:29]
  wire  _T_25 = _T_16[1] & auto_mem_in_ar_bits_addr[1]; // @[Misc.scala 213:38]
  wire  _T_26 = _T_17 | _T_25; // @[Misc.scala 213:29]
  wire  _T_29 = ~auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 209:20]
  wire  _T_30 = _T_20 & _T_29; // @[Misc.scala 212:27]
  wire  _T_31 = _T_16[0] & _T_30; // @[Misc.scala 213:38]
  wire  _T_32 = _T_23 | _T_31; // @[Misc.scala 213:29]
  wire  _T_33 = _T_20 & auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  wire  _T_34 = _T_16[0] & _T_33; // @[Misc.scala 213:38]
  wire  _T_35 = _T_23 | _T_34; // @[Misc.scala 213:29]
  wire  _T_36 = auto_mem_in_ar_bits_addr[1] & _T_29; // @[Misc.scala 212:27]
  wire  _T_37 = _T_16[0] & _T_36; // @[Misc.scala 213:38]
  wire  _T_38 = _T_26 | _T_37; // @[Misc.scala 213:29]
  wire  _T_39 = auto_mem_in_ar_bits_addr[1] & auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  wire  _T_40 = _T_16[0] & _T_39; // @[Misc.scala 213:38]
  wire  _T_41 = _T_26 | _T_40; // @[Misc.scala 213:29]
  wire [3:0] _T_44 = {_T_41,_T_38,_T_35,_T_32}; // @[Cat.scala 29:58]
  wire [3:0] _T_46 = auto_mem_in_ar_valid ? _T_44 : auto_mem_in_w_bits_strb; // @[RegisterRouter.scala 54:25]
  wire [7:0] _T_63 = _T_46[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_65 = _T_46[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_67 = _T_46[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_69 = _T_46[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_72 = {_T_69,_T_67,_T_65,_T_63}; // @[Cat.scala 29:58]
  wire  _T_91 = _T_72[1:0] == 2'h3; // @[RegisterRouter.scala 59:16]
  wire  _T_117 = _T_3 & _T_47_ready; // @[RegisterRouter.scala 59:16]
  wire  _T_129 = _T_117 & _T_4; // @[RegisterRouter.scala 59:16]
  wire  _T_132 = _T_129 & _T_53; // @[RegisterRouter.scala 59:16]
  wire  _T_98 = _T_132 & _T_91; // @[RegisterRouter.scala 59:16]
  wire [1:0] _T_171 = _T_53 ? selReg : 2'h0; // @[RegisterRouter.scala 59:16]
  wire  _T_172_bits_read = Queue_io_deq_bits_read; // @[Decoupled.scala 317:19 Decoupled.scala 318:14]
  wire  _T_172_valid = Queue_io_deq_valid; // @[Decoupled.scala 317:19 Decoupled.scala 319:15]
  wire  _T_175 = ~_T_172_bits_read; // @[RegisterRouter.scala 65:29]
  LogMagMux logMagMux ( // @[LogMagMuxDspBlock.scala 27:27]
    .clock(logMagMux_clock),
    .reset(logMagMux_reset),
    .io_in_ready(logMagMux_io_in_ready),
    .io_in_valid(logMagMux_io_in_valid),
    .io_in_bits_real(logMagMux_io_in_bits_real),
    .io_in_bits_imag(logMagMux_io_in_bits_imag),
    .io_lastIn(logMagMux_io_lastIn),
    .io_out_ready(logMagMux_io_out_ready),
    .io_out_valid(logMagMux_io_out_valid),
    .io_out_bits_real(logMagMux_io_out_bits_real),
    .io_out_bits_imag(logMagMux_io_out_bits_imag),
    .io_sel(logMagMux_io_sel),
    .io_lastOut(logMagMux_io_lastOut)
  );
  Queue Queue ( // @[Decoupled.scala 296:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_read(Queue_io_enq_bits_read),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_extra(Queue_io_enq_bits_extra),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_read(Queue_io_deq_bits_read),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_extra(Queue_io_deq_bits_extra)
  );
  assign auto_mem_in_aw_ready = _T_5 & auto_mem_in_w_valid; // @[LazyModule.scala 173:31]
  assign auto_mem_in_w_ready = _T_5 & auto_mem_in_aw_valid; // @[LazyModule.scala 173:31]
  assign auto_mem_in_b_valid = _T_172_valid & _T_175; // @[LazyModule.scala 173:31]
  assign auto_mem_in_b_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_mem_in_ar_ready = Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_valid = _T_172_valid & _T_172_bits_read; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 173:31]
  assign auto_stream_in_ready = logMagMux_io_in_ready; // @[LazyModule.scala 173:31]
  assign auto_stream_out_valid = logMagMux_io_out_valid; // @[LazyModule.scala 173:49]
  assign auto_stream_out_bits_data = {logMagMux_io_out_bits_real,logMagMux_io_out_bits_imag}; // @[LazyModule.scala 173:49]
  assign auto_stream_out_bits_last = logMagMux_io_lastOut; // @[LazyModule.scala 173:49]
  assign logMagMux_clock = clock;
  assign logMagMux_reset = reset;
  assign logMagMux_io_in_valid = auto_stream_in_valid; // @[LogMagMuxDspBlock.scala 40:30]
  assign logMagMux_io_in_bits_real = auto_stream_in_bits_data[31:16]; // @[LogMagMuxDspBlock.scala 41:30]
  assign logMagMux_io_in_bits_imag = auto_stream_in_bits_data[15:0]; // @[LogMagMuxDspBlock.scala 41:30]
  assign logMagMux_io_lastIn = auto_stream_in_bits_last; // @[LogMagMuxDspBlock.scala 44:31]
  assign logMagMux_io_out_ready = auto_stream_out_ready; // @[LogMagMuxDspBlock.scala 49:28]
  assign logMagMux_io_sel = selReg; // @[LogMagMuxDspBlock.scala 35:22]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_mem_in_ar_valid | _T_2; // @[Decoupled.scala 297:22]
  assign Queue_io_enq_bits_read = auto_mem_in_ar_valid; // @[Decoupled.scala 298:21]
  assign Queue_io_enq_bits_data = {{30'd0}, _T_171}; // @[Decoupled.scala 298:21]
  assign Queue_io_enq_bits_extra = auto_mem_in_ar_valid ? auto_mem_in_ar_bits_id : auto_mem_in_aw_bits_id; // @[Decoupled.scala 298:21]
  assign Queue_io_deq_ready = _T_172_bits_read ? auto_mem_in_r_ready : auto_mem_in_b_ready; // @[Decoupled.scala 320:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  selReg = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      selReg <= 2'h0;
    end else if (_T_98) begin
      selReg <= auto_mem_in_w_bits_data[1:0];
    end
  end
endmodule
module AXI4Splitter_4(
  input         clock,
  input         reset,
  output        auto_mem_in_aw_ready,
  input         auto_mem_in_aw_valid,
  input         auto_mem_in_aw_bits_id,
  input  [29:0] auto_mem_in_aw_bits_addr,
  output        auto_mem_in_w_ready,
  input         auto_mem_in_w_valid,
  input  [31:0] auto_mem_in_w_bits_data,
  input  [3:0]  auto_mem_in_w_bits_strb,
  input         auto_mem_in_b_ready,
  output        auto_mem_in_b_valid,
  output        auto_mem_in_b_bits_id,
  output        auto_mem_in_ar_ready,
  input         auto_mem_in_ar_valid,
  input         auto_mem_in_ar_bits_id,
  input  [29:0] auto_mem_in_ar_bits_addr,
  input  [2:0]  auto_mem_in_ar_bits_size,
  input         auto_mem_in_r_ready,
  output        auto_mem_in_r_valid,
  output        auto_mem_in_r_bits_id,
  output [31:0] auto_mem_in_r_bits_data,
  output        auto_stream_in_ready,
  input         auto_stream_in_valid,
  input  [31:0] auto_stream_in_bits_data,
  input         auto_stream_in_bits_last,
  input         auto_stream_out_1_ready,
  output        auto_stream_out_1_valid,
  output [31:0] auto_stream_out_1_bits_data,
  output        auto_stream_out_1_bits_last,
  input         auto_stream_out_0_ready,
  output        auto_stream_out_0_valid,
  output [31:0] auto_stream_out_0_bits_data,
  output        auto_stream_out_0_bits_last
);
  wire  Queue_clock; // @[Decoupled.scala 296:21]
  wire  Queue_reset; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_bits_read; // @[Decoupled.scala 296:21]
  wire [31:0] Queue_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_bits_extra; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_bits_read; // @[Decoupled.scala 296:21]
  wire [31:0] Queue_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_bits_extra; // @[Decoupled.scala 296:21]
  reg [31:0] ctrlReg; // @[Splitter.scala 27:26]
  reg [31:0] _RAND_0;
  reg [31:0] maskReg; // @[Splitter.scala 28:26]
  reg [31:0] _RAND_1;
  wire  _T_4 = auto_mem_in_aw_valid & auto_mem_in_w_valid; // @[RegisterRouter.scala 40:39]
  wire  _T_5 = auto_mem_in_ar_valid | _T_4; // @[RegisterRouter.scala 40:26]
  wire  _T_6 = ~auto_mem_in_ar_valid; // @[RegisterRouter.scala 42:29]
  wire  _T_49_ready = Queue_io_enq_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 299:17]
  wire [29:0] _T_13 = auto_mem_in_ar_valid ? auto_mem_in_ar_bits_addr : auto_mem_in_aw_bits_addr; // @[RegisterRouter.scala 48:19]
  wire [1:0] _T_53 = _T_13[3:2] & 2'h2; // @[RegisterRouter.scala 59:16]
  wire  _T_55 = _T_53 == 2'h0; // @[RegisterRouter.scala 59:16]
  wire  _T_7 = _T_49_ready & _T_6; // @[RegisterRouter.scala 42:26]
  wire [1:0] _T_16 = 2'h1 << auto_mem_in_ar_bits_size[0]; // @[OneHot.scala 65:12]
  wire [1:0] _T_18 = _T_16 | 2'h1; // @[Misc.scala 200:81]
  wire  _T_19 = auto_mem_in_ar_bits_size >= 3'h2; // @[Misc.scala 204:21]
  wire  _T_22 = ~auto_mem_in_ar_bits_addr[1]; // @[Misc.scala 209:20]
  wire  _T_24 = _T_18[1] & _T_22; // @[Misc.scala 213:38]
  wire  _T_25 = _T_19 | _T_24; // @[Misc.scala 213:29]
  wire  _T_27 = _T_18[1] & auto_mem_in_ar_bits_addr[1]; // @[Misc.scala 213:38]
  wire  _T_28 = _T_19 | _T_27; // @[Misc.scala 213:29]
  wire  _T_31 = ~auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 209:20]
  wire  _T_32 = _T_22 & _T_31; // @[Misc.scala 212:27]
  wire  _T_33 = _T_18[0] & _T_32; // @[Misc.scala 213:38]
  wire  _T_34 = _T_25 | _T_33; // @[Misc.scala 213:29]
  wire  _T_35 = _T_22 & auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  wire  _T_36 = _T_18[0] & _T_35; // @[Misc.scala 213:38]
  wire  _T_37 = _T_25 | _T_36; // @[Misc.scala 213:29]
  wire  _T_38 = auto_mem_in_ar_bits_addr[1] & _T_31; // @[Misc.scala 212:27]
  wire  _T_39 = _T_18[0] & _T_38; // @[Misc.scala 213:38]
  wire  _T_40 = _T_28 | _T_39; // @[Misc.scala 213:29]
  wire  _T_41 = auto_mem_in_ar_bits_addr[1] & auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  wire  _T_42 = _T_18[0] & _T_41; // @[Misc.scala 213:38]
  wire  _T_43 = _T_28 | _T_42; // @[Misc.scala 213:29]
  wire [3:0] _T_46 = {_T_43,_T_40,_T_37,_T_34}; // @[Cat.scala 29:58]
  wire [3:0] _T_48 = auto_mem_in_ar_valid ? _T_46 : auto_mem_in_w_bits_strb; // @[RegisterRouter.scala 54:25]
  wire [7:0] _T_67 = _T_48[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_69 = _T_48[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_71 = _T_48[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_73 = _T_48[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_76 = {_T_73,_T_71,_T_69,_T_67}; // @[Cat.scala 29:58]
  wire  _T_95 = _T_76 == 32'hffffffff; // @[RegisterRouter.scala 59:16]
  wire  _T_148 = _T_5 & _T_49_ready; // @[RegisterRouter.scala 59:16]
  wire [1:0] _T_142 = 2'h1 << _T_13[2]; // @[OneHot.scala 58:35]
  wire  _T_165 = _T_148 & _T_6; // @[RegisterRouter.scala 59:16]
  wire  _T_172 = _T_165 & _T_142[1]; // @[RegisterRouter.scala 59:16]
  wire  _T_173 = _T_172 & _T_55; // @[RegisterRouter.scala 59:16]
  wire  _T_102 = _T_173 & _T_95; // @[RegisterRouter.scala 59:16]
  wire  _T_167 = _T_165 & _T_142[0]; // @[RegisterRouter.scala 59:16]
  wire  _T_168 = _T_167 & _T_55; // @[RegisterRouter.scala 59:16]
  wire  _T_125 = _T_168 & _T_95; // @[RegisterRouter.scala 59:16]
  wire  _GEN_11 = _T_13[2] ? _T_55 : _T_55; // @[MuxLiteral.scala 48:10]
  wire [31:0] _GEN_13 = _T_13[2] ? maskReg : ctrlReg; // @[MuxLiteral.scala 48:10]
  wire  _T_223_bits_read = Queue_io_deq_bits_read; // @[Decoupled.scala 317:19 Decoupled.scala 318:14]
  wire  _T_223_valid = Queue_io_deq_valid; // @[Decoupled.scala 317:19 Decoupled.scala 319:15]
  wire  _T_226 = ~_T_223_bits_read; // @[RegisterRouter.scala 65:29]
  wire  readyOR = auto_stream_out_0_ready | auto_stream_out_1_ready; // @[Splitter.scala 45:34]
  wire  readyAND = auto_stream_out_0_ready & auto_stream_out_1_ready; // @[Splitter.scala 46:34]
  wire  _T_229 = ctrlReg == 32'h0; // @[Splitter.scala 49:19]
  wire  _T_230 = ctrlReg == 32'h1; // @[Splitter.scala 52:24]
  wire  _GEN_14 = _T_230 & readyOR; // @[Splitter.scala 52:33]
  wire  _T_233 = ~maskReg[0]; // @[Splitter.scala 62:34]
  wire  _T_237 = ~maskReg[1]; // @[Splitter.scala 62:34]
  Queue Queue ( // @[Decoupled.scala 296:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_read(Queue_io_enq_bits_read),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_extra(Queue_io_enq_bits_extra),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_read(Queue_io_deq_bits_read),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_extra(Queue_io_deq_bits_extra)
  );
  assign auto_mem_in_aw_ready = _T_7 & auto_mem_in_w_valid; // @[LazyModule.scala 173:31]
  assign auto_mem_in_w_ready = _T_7 & auto_mem_in_aw_valid; // @[LazyModule.scala 173:31]
  assign auto_mem_in_b_valid = _T_223_valid & _T_226; // @[LazyModule.scala 173:31]
  assign auto_mem_in_b_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_mem_in_ar_ready = Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_valid = _T_223_valid & _T_223_bits_read; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 173:31]
  assign auto_stream_in_ready = _T_229 ? readyAND : _GEN_14; // @[LazyModule.scala 173:31]
  assign auto_stream_out_1_valid = auto_stream_in_valid & _T_237; // @[LazyModule.scala 173:49]
  assign auto_stream_out_1_bits_data = auto_stream_in_bits_data; // @[LazyModule.scala 173:49]
  assign auto_stream_out_1_bits_last = auto_stream_in_bits_last; // @[LazyModule.scala 173:49]
  assign auto_stream_out_0_valid = auto_stream_in_valid & _T_233; // @[LazyModule.scala 173:49]
  assign auto_stream_out_0_bits_data = auto_stream_in_bits_data; // @[LazyModule.scala 173:49]
  assign auto_stream_out_0_bits_last = auto_stream_in_bits_last; // @[LazyModule.scala 173:49]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_mem_in_ar_valid | _T_4; // @[Decoupled.scala 297:22]
  assign Queue_io_enq_bits_read = auto_mem_in_ar_valid; // @[Decoupled.scala 298:21]
  assign Queue_io_enq_bits_data = _GEN_11 ? _GEN_13 : 32'h0; // @[Decoupled.scala 298:21]
  assign Queue_io_enq_bits_extra = auto_mem_in_ar_valid ? auto_mem_in_ar_bits_id : auto_mem_in_aw_bits_id; // @[Decoupled.scala 298:21]
  assign Queue_io_deq_ready = _T_223_bits_read ? auto_mem_in_r_ready : auto_mem_in_b_ready; // @[Decoupled.scala 320:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ctrlReg = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  maskReg = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      ctrlReg <= 32'h0;
    end else if (_T_125) begin
      ctrlReg <= auto_mem_in_w_bits_data;
    end
    if (reset) begin
      maskReg <= 32'h0;
    end else if (_T_102) begin
      maskReg <= auto_mem_in_w_bits_data;
    end
  end
endmodule
module AXI4StreamMux_6(
  input         clock,
  input         reset,
  output        auto_register_in_aw_ready,
  input         auto_register_in_aw_valid,
  input         auto_register_in_aw_bits_id,
  input  [29:0] auto_register_in_aw_bits_addr,
  output        auto_register_in_w_ready,
  input         auto_register_in_w_valid,
  input  [31:0] auto_register_in_w_bits_data,
  input  [3:0]  auto_register_in_w_bits_strb,
  input         auto_register_in_b_ready,
  output        auto_register_in_b_valid,
  output        auto_register_in_b_bits_id,
  output        auto_register_in_ar_ready,
  input         auto_register_in_ar_valid,
  input         auto_register_in_ar_bits_id,
  input  [29:0] auto_register_in_ar_bits_addr,
  input  [2:0]  auto_register_in_ar_bits_size,
  input         auto_register_in_r_ready,
  output        auto_register_in_r_valid,
  output        auto_register_in_r_bits_id,
  output [31:0] auto_register_in_r_bits_data,
  output        auto_stream_in_2_ready,
  input         auto_stream_in_2_valid,
  input  [31:0] auto_stream_in_2_bits_data,
  input         auto_stream_in_2_bits_last,
  output        auto_stream_in_1_ready,
  input         auto_stream_in_1_valid,
  input  [31:0] auto_stream_in_1_bits_data,
  input         auto_stream_in_1_bits_last,
  output        auto_stream_in_0_ready,
  input         auto_stream_in_0_valid,
  input  [31:0] auto_stream_in_0_bits_data,
  input         auto_stream_in_0_bits_last,
  input         auto_stream_out_0_ready,
  output        auto_stream_out_0_valid,
  output [31:0] auto_stream_out_0_bits_data,
  output        auto_stream_out_0_bits_last
);
  wire  Queue_clock; // @[Decoupled.scala 296:21]
  wire  Queue_reset; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_bits_read; // @[Decoupled.scala 296:21]
  wire [31:0] Queue_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_bits_extra; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_bits_read; // @[Decoupled.scala 296:21]
  wire [31:0] Queue_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_bits_extra; // @[Decoupled.scala 296:21]
  reg [2:0] sels_0; // @[Mux.scala 32:23]
  reg [31:0] _RAND_0;
  reg [2:0] sels_1; // @[Mux.scala 32:23]
  reg [31:0] _RAND_1;
  wire  _T_3 = sels_0 == 3'h0; // @[Mux.scala 45:28]
  wire  _GEN_7 = _T_3 & auto_stream_in_0_valid; // @[Mux.scala 45:41]
  wire  _GEN_8 = _T_3 & auto_stream_out_0_ready; // @[Mux.scala 45:41]
  wire  _T_4 = sels_0 == 3'h1; // @[Mux.scala 45:28]
  wire  _GEN_12 = _T_4 ? auto_stream_in_1_bits_last : auto_stream_in_0_bits_last; // @[Mux.scala 45:41]
  wire [31:0] _GEN_15 = _T_4 ? auto_stream_in_1_bits_data : auto_stream_in_0_bits_data; // @[Mux.scala 45:41]
  wire  _GEN_16 = _T_4 ? auto_stream_in_1_valid : _GEN_7; // @[Mux.scala 45:41]
  wire  _GEN_17 = _T_4 & auto_stream_out_0_ready; // @[Mux.scala 45:41]
  wire  _T_5 = sels_0 == 3'h2; // @[Mux.scala 45:28]
  wire  _GEN_21 = _T_5 ? auto_stream_in_2_bits_last : _GEN_12; // @[Mux.scala 45:41]
  wire [31:0] _GEN_24 = _T_5 ? auto_stream_in_2_bits_data : _GEN_15; // @[Mux.scala 45:41]
  wire  _GEN_25 = _T_5 ? auto_stream_in_2_valid : _GEN_16; // @[Mux.scala 45:41]
  wire  _GEN_26 = _T_5 & auto_stream_out_0_ready; // @[Mux.scala 45:41]
  wire  _T_6 = sels_0 == 3'h3; // @[Mux.scala 45:28]
  wire  _GEN_30 = _T_6 ? 1'h0 : _GEN_21; // @[Mux.scala 45:41]
  wire [31:0] _GEN_33 = _T_6 ? 32'hffffffff : _GEN_24; // @[Mux.scala 45:41]
  wire  _GEN_34 = _T_6 | _GEN_25; // @[Mux.scala 45:41]
  wire  _T_7 = sels_0 == 3'h4; // @[Mux.scala 45:28]
  wire  _T_8 = sels_0 == sels_1; // @[Mux.scala 40:46]
  wire [2:0] _T_10 = _T_8 ? 3'h5 : sels_1; // @[Mux.scala 41:29]
  wire  _T_11 = _T_10 == 3'h0; // @[Mux.scala 45:28]
  wire  _T_12 = _T_10 == 3'h1; // @[Mux.scala 45:28]
  wire  _T_13 = _T_10 == 3'h2; // @[Mux.scala 45:28]
  wire  _T_17 = auto_register_in_aw_valid & auto_register_in_w_valid; // @[RegisterRouter.scala 40:39]
  wire  _T_18 = auto_register_in_ar_valid | _T_17; // @[RegisterRouter.scala 40:26]
  wire  _T_19 = ~auto_register_in_ar_valid; // @[RegisterRouter.scala 42:29]
  wire  _T_62_ready = Queue_io_enq_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 299:17]
  wire [29:0] _T_26 = auto_register_in_ar_valid ? auto_register_in_ar_bits_addr : auto_register_in_aw_bits_addr; // @[RegisterRouter.scala 48:19]
  wire [1:0] _T_66 = _T_26[3:2] & 2'h2; // @[RegisterRouter.scala 59:16]
  wire  _T_68 = _T_66 == 2'h0; // @[RegisterRouter.scala 59:16]
  wire  _T_20 = _T_62_ready & _T_19; // @[RegisterRouter.scala 42:26]
  wire [1:0] _T_29 = 2'h1 << auto_register_in_ar_bits_size[0]; // @[OneHot.scala 65:12]
  wire [1:0] _T_31 = _T_29 | 2'h1; // @[Misc.scala 200:81]
  wire  _T_32 = auto_register_in_ar_bits_size >= 3'h2; // @[Misc.scala 204:21]
  wire  _T_35 = ~auto_register_in_ar_bits_addr[1]; // @[Misc.scala 209:20]
  wire  _T_37 = _T_31[1] & _T_35; // @[Misc.scala 213:38]
  wire  _T_38 = _T_32 | _T_37; // @[Misc.scala 213:29]
  wire  _T_40 = _T_31[1] & auto_register_in_ar_bits_addr[1]; // @[Misc.scala 213:38]
  wire  _T_41 = _T_32 | _T_40; // @[Misc.scala 213:29]
  wire  _T_44 = ~auto_register_in_ar_bits_addr[0]; // @[Misc.scala 209:20]
  wire  _T_45 = _T_35 & _T_44; // @[Misc.scala 212:27]
  wire  _T_46 = _T_31[0] & _T_45; // @[Misc.scala 213:38]
  wire  _T_47 = _T_38 | _T_46; // @[Misc.scala 213:29]
  wire  _T_48 = _T_35 & auto_register_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  wire  _T_49 = _T_31[0] & _T_48; // @[Misc.scala 213:38]
  wire  _T_50 = _T_38 | _T_49; // @[Misc.scala 213:29]
  wire  _T_51 = auto_register_in_ar_bits_addr[1] & _T_44; // @[Misc.scala 212:27]
  wire  _T_52 = _T_31[0] & _T_51; // @[Misc.scala 213:38]
  wire  _T_53 = _T_41 | _T_52; // @[Misc.scala 213:29]
  wire  _T_54 = auto_register_in_ar_bits_addr[1] & auto_register_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  wire  _T_55 = _T_31[0] & _T_54; // @[Misc.scala 213:38]
  wire  _T_56 = _T_41 | _T_55; // @[Misc.scala 213:29]
  wire [3:0] _T_59 = {_T_56,_T_53,_T_50,_T_47}; // @[Cat.scala 29:58]
  wire [3:0] _T_61 = auto_register_in_ar_valid ? _T_59 : auto_register_in_w_bits_strb; // @[RegisterRouter.scala 54:25]
  wire [7:0] _T_80 = _T_61[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_82 = _T_61[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_84 = _T_61[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_86 = _T_61[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_89 = {_T_86,_T_84,_T_82,_T_80}; // @[Cat.scala 29:58]
  wire  _T_108 = _T_89[2:0] == 3'h7; // @[RegisterRouter.scala 59:16]
  wire  _T_161 = _T_18 & _T_62_ready; // @[RegisterRouter.scala 59:16]
  wire [1:0] _T_155 = 2'h1 << _T_26[2]; // @[OneHot.scala 58:35]
  wire  _T_178 = _T_161 & _T_19; // @[RegisterRouter.scala 59:16]
  wire  _T_185 = _T_178 & _T_155[1]; // @[RegisterRouter.scala 59:16]
  wire  _T_186 = _T_185 & _T_68; // @[RegisterRouter.scala 59:16]
  wire  _T_115 = _T_186 & _T_108; // @[RegisterRouter.scala 59:16]
  wire  _T_180 = _T_178 & _T_155[0]; // @[RegisterRouter.scala 59:16]
  wire  _T_181 = _T_180 & _T_68; // @[RegisterRouter.scala 59:16]
  wire  _T_138 = _T_181 & _T_108; // @[RegisterRouter.scala 59:16]
  wire  _GEN_101 = _T_26[2] ? _T_68 : _T_68; // @[MuxLiteral.scala 48:10]
  wire [2:0] _GEN_103 = _T_26[2] ? sels_1 : sels_0; // @[MuxLiteral.scala 48:10]
  wire [2:0] _T_235 = _GEN_101 ? _GEN_103 : 3'h0; // @[RegisterRouter.scala 59:16]
  wire  _T_236_bits_read = Queue_io_deq_bits_read; // @[Decoupled.scala 317:19 Decoupled.scala 318:14]
  wire  _T_236_valid = Queue_io_deq_valid; // @[Decoupled.scala 317:19 Decoupled.scala 319:15]
  wire  _T_239 = ~_T_236_bits_read; // @[RegisterRouter.scala 65:29]
  Queue Queue ( // @[Decoupled.scala 296:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_read(Queue_io_enq_bits_read),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_extra(Queue_io_enq_bits_extra),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_read(Queue_io_deq_bits_read),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_extra(Queue_io_deq_bits_extra)
  );
  assign auto_register_in_aw_ready = _T_20 & auto_register_in_w_valid; // @[LazyModule.scala 173:31]
  assign auto_register_in_w_ready = _T_20 & auto_register_in_aw_valid; // @[LazyModule.scala 173:31]
  assign auto_register_in_b_valid = _T_236_valid & _T_239; // @[LazyModule.scala 173:31]
  assign auto_register_in_b_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_register_in_ar_ready = Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_register_in_r_valid = _T_236_valid & _T_236_bits_read; // @[LazyModule.scala 173:31]
  assign auto_register_in_r_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_register_in_r_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 173:31]
  assign auto_stream_in_2_ready = _T_13 | _GEN_26; // @[LazyModule.scala 173:31]
  assign auto_stream_in_1_ready = _T_12 | _GEN_17; // @[LazyModule.scala 173:31]
  assign auto_stream_in_0_ready = _T_11 | _GEN_8; // @[LazyModule.scala 173:31]
  assign auto_stream_out_0_valid = _T_7 | _GEN_34; // @[LazyModule.scala 173:49]
  assign auto_stream_out_0_bits_data = _T_7 ? 32'h0 : _GEN_33; // @[LazyModule.scala 173:49]
  assign auto_stream_out_0_bits_last = _T_7 ? 1'h0 : _GEN_30; // @[LazyModule.scala 173:49]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_register_in_ar_valid | _T_17; // @[Decoupled.scala 297:22]
  assign Queue_io_enq_bits_read = auto_register_in_ar_valid; // @[Decoupled.scala 298:21]
  assign Queue_io_enq_bits_data = {{29'd0}, _T_235}; // @[Decoupled.scala 298:21]
  assign Queue_io_enq_bits_extra = auto_register_in_ar_valid ? auto_register_in_ar_bits_id : auto_register_in_aw_bits_id; // @[Decoupled.scala 298:21]
  assign Queue_io_deq_ready = _T_236_bits_read ? auto_register_in_r_ready : auto_register_in_b_ready; // @[Decoupled.scala 320:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  sels_0 = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  sels_1 = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      sels_0 <= 3'h5;
    end else if (_T_138) begin
      sels_0 <= auto_register_in_w_bits_data[2:0];
    end
    if (reset) begin
      sels_1 <= 3'h5;
    end else if (_T_115) begin
      sels_1 <= auto_register_in_w_bits_data[2:0];
    end
  end
endmodule
module AXI4StreamMux_7(
  input         clock,
  input         reset,
  output        auto_register_in_aw_ready,
  input         auto_register_in_aw_valid,
  input         auto_register_in_aw_bits_id,
  input  [29:0] auto_register_in_aw_bits_addr,
  output        auto_register_in_w_ready,
  input         auto_register_in_w_valid,
  input  [31:0] auto_register_in_w_bits_data,
  input  [3:0]  auto_register_in_w_bits_strb,
  input         auto_register_in_b_ready,
  output        auto_register_in_b_valid,
  output        auto_register_in_b_bits_id,
  output        auto_register_in_ar_ready,
  input         auto_register_in_ar_valid,
  input         auto_register_in_ar_bits_id,
  input  [29:0] auto_register_in_ar_bits_addr,
  input  [2:0]  auto_register_in_ar_bits_size,
  input         auto_register_in_r_ready,
  output        auto_register_in_r_valid,
  output        auto_register_in_r_bits_id,
  output [31:0] auto_register_in_r_bits_data,
  output        auto_stream_in_ready,
  input         auto_stream_in_valid,
  input  [31:0] auto_stream_in_bits_data,
  input         auto_stream_in_bits_last,
  input         auto_stream_out_1_ready,
  output        auto_stream_out_1_valid,
  output [31:0] auto_stream_out_1_bits_data,
  output        auto_stream_out_1_bits_last
);
  wire  Queue_clock; // @[Decoupled.scala 296:21]
  wire  Queue_reset; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_bits_read; // @[Decoupled.scala 296:21]
  wire [31:0] Queue_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_bits_extra; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_bits_read; // @[Decoupled.scala 296:21]
  wire [31:0] Queue_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_bits_extra; // @[Decoupled.scala 296:21]
  reg  sels_0; // @[Mux.scala 32:23]
  reg [31:0] _RAND_0;
  reg  sels_1; // @[Mux.scala 32:23]
  reg [31:0] _RAND_1;
  wire  _T_3 = ~sels_0; // @[Mux.scala 45:28]
  wire  _T_4 = sels_0 == sels_1; // @[Mux.scala 40:46]
  wire  _T_6 = _T_4 | sels_1; // @[Mux.scala 41:29]
  wire  _T_7 = ~_T_6; // @[Mux.scala 45:28]
  wire  _T_9 = auto_register_in_aw_valid & auto_register_in_w_valid; // @[RegisterRouter.scala 40:39]
  wire  _T_10 = auto_register_in_ar_valid | _T_9; // @[RegisterRouter.scala 40:26]
  wire  _T_11 = ~auto_register_in_ar_valid; // @[RegisterRouter.scala 42:29]
  wire  _T_54_ready = Queue_io_enq_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 299:17]
  wire [29:0] _T_18 = auto_register_in_ar_valid ? auto_register_in_ar_bits_addr : auto_register_in_aw_bits_addr; // @[RegisterRouter.scala 48:19]
  wire [1:0] _T_58 = _T_18[3:2] & 2'h2; // @[RegisterRouter.scala 59:16]
  wire  _T_60 = _T_58 == 2'h0; // @[RegisterRouter.scala 59:16]
  wire  _T_12 = _T_54_ready & _T_11; // @[RegisterRouter.scala 42:26]
  wire [1:0] _T_21 = 2'h1 << auto_register_in_ar_bits_size[0]; // @[OneHot.scala 65:12]
  wire [1:0] _T_23 = _T_21 | 2'h1; // @[Misc.scala 200:81]
  wire  _T_24 = auto_register_in_ar_bits_size >= 3'h2; // @[Misc.scala 204:21]
  wire  _T_27 = ~auto_register_in_ar_bits_addr[1]; // @[Misc.scala 209:20]
  wire  _T_29 = _T_23[1] & _T_27; // @[Misc.scala 213:38]
  wire  _T_30 = _T_24 | _T_29; // @[Misc.scala 213:29]
  wire  _T_32 = _T_23[1] & auto_register_in_ar_bits_addr[1]; // @[Misc.scala 213:38]
  wire  _T_33 = _T_24 | _T_32; // @[Misc.scala 213:29]
  wire  _T_36 = ~auto_register_in_ar_bits_addr[0]; // @[Misc.scala 209:20]
  wire  _T_37 = _T_27 & _T_36; // @[Misc.scala 212:27]
  wire  _T_38 = _T_23[0] & _T_37; // @[Misc.scala 213:38]
  wire  _T_39 = _T_30 | _T_38; // @[Misc.scala 213:29]
  wire  _T_40 = _T_27 & auto_register_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  wire  _T_41 = _T_23[0] & _T_40; // @[Misc.scala 213:38]
  wire  _T_42 = _T_30 | _T_41; // @[Misc.scala 213:29]
  wire  _T_43 = auto_register_in_ar_bits_addr[1] & _T_36; // @[Misc.scala 212:27]
  wire  _T_44 = _T_23[0] & _T_43; // @[Misc.scala 213:38]
  wire  _T_45 = _T_33 | _T_44; // @[Misc.scala 213:29]
  wire  _T_46 = auto_register_in_ar_bits_addr[1] & auto_register_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  wire  _T_47 = _T_23[0] & _T_46; // @[Misc.scala 213:38]
  wire  _T_48 = _T_33 | _T_47; // @[Misc.scala 213:29]
  wire [3:0] _T_51 = {_T_48,_T_45,_T_42,_T_39}; // @[Cat.scala 29:58]
  wire [3:0] _T_53 = auto_register_in_ar_valid ? _T_51 : auto_register_in_w_bits_strb; // @[RegisterRouter.scala 54:25]
  wire [7:0] _T_72 = _T_53[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_74 = _T_53[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_76 = _T_53[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_78 = _T_53[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_81 = {_T_78,_T_76,_T_74,_T_72}; // @[Cat.scala 29:58]
  wire  _T_153 = _T_10 & _T_54_ready; // @[RegisterRouter.scala 59:16]
  wire [1:0] _T_147 = 2'h1 << _T_18[2]; // @[OneHot.scala 58:35]
  wire  _T_170 = _T_153 & _T_11; // @[RegisterRouter.scala 59:16]
  wire  _T_177 = _T_170 & _T_147[1]; // @[RegisterRouter.scala 59:16]
  wire  _T_178 = _T_177 & _T_60; // @[RegisterRouter.scala 59:16]
  wire  _T_107 = _T_178 & _T_81[0]; // @[RegisterRouter.scala 59:16]
  wire  _GEN_18 = _T_107 ? auto_register_in_w_bits_data[0] : sels_1; // @[RegField.scala 134:88]
  wire  _T_172 = _T_170 & _T_147[0]; // @[RegisterRouter.scala 59:16]
  wire  _T_173 = _T_172 & _T_60; // @[RegisterRouter.scala 59:16]
  wire  _T_130 = _T_173 & _T_81[0]; // @[RegisterRouter.scala 59:16]
  wire  _GEN_19 = _T_130 ? auto_register_in_w_bits_data[0] : sels_0; // @[RegField.scala 134:88]
  wire  _GEN_29 = _T_18[2] ? _T_60 : _T_60; // @[MuxLiteral.scala 48:10]
  wire  _GEN_31 = _T_18[2] ? sels_1 : sels_0; // @[MuxLiteral.scala 48:10]
  wire  _T_227 = _GEN_29 & _GEN_31; // @[RegisterRouter.scala 59:16]
  wire  _T_228_bits_read = Queue_io_deq_bits_read; // @[Decoupled.scala 317:19 Decoupled.scala 318:14]
  wire  _T_228_valid = Queue_io_deq_valid; // @[Decoupled.scala 317:19 Decoupled.scala 319:15]
  wire  _T_231 = ~_T_228_bits_read; // @[RegisterRouter.scala 65:29]
  Queue Queue ( // @[Decoupled.scala 296:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_read(Queue_io_enq_bits_read),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_extra(Queue_io_enq_bits_extra),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_read(Queue_io_deq_bits_read),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_extra(Queue_io_deq_bits_extra)
  );
  assign auto_register_in_aw_ready = _T_12 & auto_register_in_w_valid; // @[LazyModule.scala 173:31]
  assign auto_register_in_w_ready = _T_12 & auto_register_in_aw_valid; // @[LazyModule.scala 173:31]
  assign auto_register_in_b_valid = _T_228_valid & _T_231; // @[LazyModule.scala 173:31]
  assign auto_register_in_b_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_register_in_ar_ready = Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_register_in_r_valid = _T_228_valid & _T_228_bits_read; // @[LazyModule.scala 173:31]
  assign auto_register_in_r_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_register_in_r_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 173:31]
  assign auto_stream_in_ready = _T_7 ? auto_stream_out_1_ready : _T_3; // @[LazyModule.scala 173:31]
  assign auto_stream_out_1_valid = _T_7 & auto_stream_in_valid; // @[LazyModule.scala 173:49]
  assign auto_stream_out_1_bits_data = auto_stream_in_bits_data; // @[LazyModule.scala 173:49]
  assign auto_stream_out_1_bits_last = auto_stream_in_bits_last; // @[LazyModule.scala 173:49]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_register_in_ar_valid | _T_9; // @[Decoupled.scala 297:22]
  assign Queue_io_enq_bits_read = auto_register_in_ar_valid; // @[Decoupled.scala 298:21]
  assign Queue_io_enq_bits_data = {{31'd0}, _T_227}; // @[Decoupled.scala 298:21]
  assign Queue_io_enq_bits_extra = auto_register_in_ar_valid ? auto_register_in_ar_bits_id : auto_register_in_aw_bits_id; // @[Decoupled.scala 298:21]
  assign Queue_io_deq_ready = _T_228_bits_read ? auto_register_in_r_ready : auto_register_in_b_ready; // @[Decoupled.scala 320:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  sels_0 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  sels_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    sels_0 <= reset | _GEN_19;
    sels_1 <= reset | _GEN_18;
  end
endmodule
module Accumulator(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [15:0] io_in_bits,
  input         io_lastIn,
  input  [7:0]  io_accDepthReg,
  input  [16:0] io_accWindowsReg,
  input         io_out_ready,
  output        io_out_valid,
  output [15:0] io_out_bits,
  output        io_lastOut
);
  reg [31:0] mem [0:127]; // @[Accumulator.scala 35:24]
  reg [31:0] _RAND_0;
  wire [31:0] mem__T_189_data; // @[Accumulator.scala 35:24]
  wire [6:0] mem__T_189_addr; // @[Accumulator.scala 35:24]
  wire [31:0] mem__T_235_data; // @[Accumulator.scala 35:24]
  wire [6:0] mem__T_235_addr; // @[Accumulator.scala 35:24]
  wire  mem__T_235_mask; // @[Accumulator.scala 35:24]
  wire  mem__T_235_en; // @[Accumulator.scala 35:24]
  reg  mem__T_189_en_pipe_0;
  reg [31:0] _RAND_1;
  reg [6:0] mem__T_189_addr_pipe_0;
  reg [31:0] _RAND_2;
  wire  readEn = io_in_ready & io_in_valid; // @[Decoupled.scala 40:37]
  reg  writeEn; // @[Accumulator.scala 38:24]
  reg [31:0] _RAND_3;
  reg [15:0] inDelayed; // @[Accumulator.scala 39:26]
  reg [31:0] _RAND_4;
  reg [15:0] cntWindows; // @[Accumulator.scala 40:27]
  reg [31:0] _RAND_5;
  reg [6:0] cntLoad; // @[Accumulator.scala 41:24]
  reg [31:0] _RAND_6;
  reg [6:0] cntAcc; // @[Accumulator.scala 42:23]
  reg [31:0] _RAND_7;
  reg [2:0] state; // @[Accumulator.scala 50:22]
  reg [31:0] _RAND_8;
  reg [2:0] statePrev; // @[Accumulator.scala 51:26]
  reg [31:0] _RAND_9;
  reg  last; // @[Accumulator.scala 53:21]
  reg [31:0] _RAND_10;
  wire  _T_3 = 3'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_7 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire [7:0] _T_9 = io_accDepthReg - 8'h1; // @[Accumulator.scala 66:40]
  wire [7:0] _GEN_34 = {{1'd0}, cntAcc}; // @[Accumulator.scala 66:20]
  wire  _T_10 = _GEN_34 == _T_9; // @[Accumulator.scala 66:20]
  wire  _T_12 = _T_10 & readEn; // @[Accumulator.scala 66:47]
  wire  _T_13 = _T_12 & io_lastIn; // @[Accumulator.scala 66:63]
  wire  _T_21 = 3'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_23 = readEn & io_lastIn; // @[Accumulator.scala 75:26]
  wire  _T_24 = ~io_out_ready; // @[Accumulator.scala 77:15]
  wire  _GEN_3 = _T_24 | last; // @[Accumulator.scala 77:30]
  wire [16:0] _T_26 = io_accWindowsReg - 17'h1; // @[Accumulator.scala 81:51]
  wire [16:0] _GEN_36 = {{1'd0}, cntWindows}; // @[Accumulator.scala 81:29]
  wire  _T_27 = _GEN_36 == _T_26; // @[Accumulator.scala 81:29]
  wire  _T_29 = _T_27 & readEn; // @[Accumulator.scala 81:58]
  wire  _T_33 = _T_29 & _T_10; // @[Accumulator.scala 81:72]
  wire  _T_36 = 3'h3 == state; // @[Conditional.scala 37:30]
  wire [7:0] _GEN_38 = {{1'd0}, cntLoad}; // @[Accumulator.scala 90:26]
  wire  _T_41 = _GEN_38 == _T_9; // @[Accumulator.scala 90:26]
  wire  _T_42 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  wire  _T_43 = _T_41 & _T_42; // @[Accumulator.scala 90:53]
  wire  _T_46 = _GEN_34 < _T_9; // @[Accumulator.scala 90:80]
  wire  _T_47 = _T_43 & _T_46; // @[Accumulator.scala 90:70]
  wire  _T_54 = _T_43 & readEn; // @[Accumulator.scala 93:70]
  wire  _T_58 = _T_54 & _T_10; // @[Accumulator.scala 93:86]
  wire  _T_61 = 3'h4 == state; // @[Conditional.scala 37:30]
  wire  _T_62 = state == 3'h3; // @[Accumulator.scala 105:30]
  wire  _T_63 = state == 3'h4; // @[Accumulator.scala 105:65]
  wire  loadingStates = _T_62 | _T_63; // @[Accumulator.scala 105:55]
  wire  _T_64 = state == 3'h1; // @[Accumulator.scala 106:34]
  wire  storingInitStates = _T_64 | _T_62; // @[Accumulator.scala 106:56]
  wire  _T_66 = state == 3'h2; // @[Accumulator.scala 107:26]
  wire  _T_67 = statePrev == 3'h1; // @[Accumulator.scala 107:62]
  wire  _T_68 = _T_66 & _T_67; // @[Accumulator.scala 107:49]
  wire  _T_69 = statePrev == 3'h3; // @[Accumulator.scala 107:98]
  wire  _T_71 = _T_69 & _T_64; // @[Accumulator.scala 107:122]
  wire  _T_72 = _T_68 | _T_71; // @[Accumulator.scala 107:84]
  wire  _T_75 = _T_69 & _T_66; // @[Accumulator.scala 107:191]
  wire  isTransit = _T_72 | _T_75; // @[Accumulator.scala 107:153]
  wire  isOnlyOneFrame = _T_63 & _T_67; // @[Accumulator.scala 108:47]
  reg  doNotScale; // @[Accumulator.scala 109:27]
  reg [31:0] _RAND_11;
  wire  _T_78 = statePrev == 3'h2; // @[Accumulator.scala 110:38]
  wire  isPrevStoreAndAcc = _T_78 & _T_62; // @[Accumulator.scala 110:62]
  wire  _GEN_19 = isOnlyOneFrame | doNotScale; // @[Accumulator.scala 116:24]
  wire  _T_88 = state == 3'h0; // @[Accumulator.scala 119:15]
  wire  _T_89 = storingInitStates | isTransit; // @[Accumulator.scala 123:28]
  wire  _T_90 = ~isPrevStoreAndAcc; // @[Accumulator.scala 123:45]
  wire  _T_91 = _T_89 & _T_90; // @[Accumulator.scala 123:42]
  wire  _T_92 = _T_91 | isOnlyOneFrame; // @[Accumulator.scala 123:64]
  wire [31:0] readVal = mem__T_189_data; // @[Accumulator.scala 43:21 Accumulator.scala 172:11]
  wire [31:0] _GEN_44 = {{16{inDelayed[15]}},inDelayed}; // @[FixedPointTypeClass.scala 20:58]
  wire [31:0] _T_95 = $signed(_GEN_44) + $signed(readVal); // @[FixedPointTypeClass.scala 20:58]
  wire [31:0] _GEN_21 = _T_92 ? $signed({{16{inDelayed[15]}},inDelayed}) : $signed(_T_95); // @[Accumulator.scala 123:83]
  wire [6:0] _T_98 = cntAcc + 7'h1; // @[Accumulator.scala 130:22]
  wire  _T_99 = loadingStates & io_out_ready; // @[Accumulator.scala 133:23]
  wire [6:0] _T_101 = cntLoad + 7'h1; // @[Accumulator.scala 134:24]
  wire [15:0] _T_111 = cntWindows + 16'h1; // @[Accumulator.scala 142:30]
  wire  _T_115 = _T_27 & _T_12; // @[Accumulator.scala 145:49]
  wire  _T_116 = last & io_out_ready; // @[Accumulator.scala 160:46]
  wire [6:0] loadAddress = _T_116 ? _T_101 : cntLoad; // @[Accumulator.scala 160:40]
  wire [6:0] readAddress = loadingStates ? loadAddress : cntAcc; // @[Accumulator.scala 167:24]
  wire  _T_195 = io_accWindowsReg[15:8] != 8'h0; // @[CircuitMath.scala 37:22]
  wire  _T_198 = io_accWindowsReg[15:12] != 4'h0; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_202 = io_accWindowsReg[14] ? 2'h2 : {{1'd0}, io_accWindowsReg[13]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_203 = io_accWindowsReg[15] ? 2'h3 : _T_202; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_207 = io_accWindowsReg[10] ? 2'h2 : {{1'd0}, io_accWindowsReg[9]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_208 = io_accWindowsReg[11] ? 2'h3 : _T_207; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_209 = _T_198 ? _T_203 : _T_208; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_210 = {_T_198,_T_209}; // @[Cat.scala 29:58]
  wire  _T_213 = io_accWindowsReg[7:4] != 4'h0; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_217 = io_accWindowsReg[6] ? 2'h2 : {{1'd0}, io_accWindowsReg[5]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_218 = io_accWindowsReg[7] ? 2'h3 : _T_217; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_222 = io_accWindowsReg[2] ? 2'h2 : {{1'd0}, io_accWindowsReg[1]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_223 = io_accWindowsReg[3] ? 2'h3 : _T_222; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_224 = _T_213 ? _T_218 : _T_223; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_225 = {_T_213,_T_224}; // @[Cat.scala 29:58]
  wire [2:0] _T_226 = _T_195 ? _T_210 : _T_225; // @[CircuitMath.scala 38:21]
  wire [3:0] _T_227 = {_T_195,_T_226}; // @[Cat.scala 29:58]
  wire [3:0] _T_228 = io_accWindowsReg[16] ? 4'h0 : _T_227; // @[CircuitMath.scala 38:21]
  wire [4:0] _T_229 = {io_accWindowsReg[16],_T_228}; // @[Cat.scala 29:58]
  wire [31:0] _T_230 = $signed(readVal) >>> _T_229; // @[FixedPointTypeClass.scala 118:51]
  wire [31:0] _T_231 = doNotScale ? $signed(readVal) : $signed(_T_230); // @[Accumulator.scala 178:17]
  reg [6:0] _T_232; // @[Accumulator.scala 184:22]
  reg [31:0] _RAND_12;
  wire [31:0] writeVal = _GEN_21; // @[Accumulator.scala 44:22 Accumulator.scala 124:14 Accumulator.scala 127:14]
  reg  _T_236; // @[Accumulator.scala 187:26]
  reg [31:0] _RAND_13;
  wire  _T_237 = state != 3'h0; // @[Accumulator.scala 187:51]
  reg [6:0] _T_239; // @[Accumulator.scala 188:27]
  reg [31:0] _RAND_14;
  wire [7:0] _GEN_47 = {{1'd0}, _T_239}; // @[Accumulator.scala 188:57]
  wire  _T_242 = _GEN_47 == _T_9; // @[Accumulator.scala 188:57]
  wire  _T_244 = _T_242 & _T_42; // @[Accumulator.scala 188:84]
  wire  _T_247 = ~loadingStates; // @[Accumulator.scala 193:22]
  wire  _T_248 = state != 3'h4; // @[Accumulator.scala 193:63]
  wire  _T_249 = io_out_ready & _T_248; // @[Accumulator.scala 193:54]
  assign mem__T_189_addr = mem__T_189_addr_pipe_0;
  assign mem__T_189_data = mem[mem__T_189_addr]; // @[Accumulator.scala 35:24]
  assign mem__T_235_data = writeVal;
  assign mem__T_235_addr = _T_232;
  assign mem__T_235_mask = 1'h1;
  assign mem__T_235_en = writeEn;
  assign io_in_ready = _T_247 | _T_249; // @[Accumulator.scala 193:18]
  assign io_out_valid = _T_236 & _T_237; // @[Accumulator.scala 187:16]
  assign io_out_bits = _T_231[15:0]; // @[Accumulator.scala 190:16]
  assign io_lastOut = _T_244 & _T_63; // @[Accumulator.scala 188:16]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    mem[initvar] = _RAND_0[31:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  mem__T_189_en_pipe_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  mem__T_189_addr_pipe_0 = _RAND_2[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  writeEn = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  inDelayed = _RAND_4[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  cntWindows = _RAND_5[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  cntLoad = _RAND_6[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  cntAcc = _RAND_7[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  state = _RAND_8[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  statePrev = _RAND_9[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  last = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  doNotScale = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_232 = _RAND_12[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_236 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_239 = _RAND_14[6:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(mem__T_235_en & mem__T_235_mask) begin
      mem[mem__T_235_addr] <= mem__T_235_data; // @[Accumulator.scala 35:24]
    end
    mem__T_189_en_pipe_0 <= 1'h1;
    if (loadingStates) begin
      if (_T_116) begin
        mem__T_189_addr_pipe_0 <= _T_101;
      end else begin
        mem__T_189_addr_pipe_0 <= cntLoad;
      end
    end else begin
      mem__T_189_addr_pipe_0 <= cntAcc;
    end
    if (reset) begin
      writeEn <= 1'h0;
    end else begin
      writeEn <= readEn;
    end
    inDelayed <= io_in_bits;
    if (reset) begin
      cntWindows <= 16'h0;
    end else if (_T_115) begin
      cntWindows <= 16'h0;
    end else if (_T_12) begin
      cntWindows <= _T_111;
    end
    if (reset) begin
      cntLoad <= 7'h0;
    end else if (_T_43) begin
      cntLoad <= 7'h0;
    end else if (_T_99) begin
      cntLoad <= _T_101;
    end else if (_T_99) begin
      cntLoad <= _T_101;
    end
    if (reset) begin
      cntAcc <= 7'h0;
    end else if (_T_12) begin
      cntAcc <= 7'h0;
    end else if (readEn) begin
      cntAcc <= _T_98;
    end
    if (reset) begin
      state <= 3'h0;
    end else if (_T_3) begin
      if (readEn) begin
        state <= 3'h1;
      end
    end else if (_T_7) begin
      if (_T_13) begin
        state <= 3'h4;
      end else if (_T_12) begin
        state <= 3'h2;
      end
    end else if (_T_21) begin
      if (_T_23) begin
        state <= 3'h4;
      end else if (_T_33) begin
        state <= 3'h3;
      end
    end else if (_T_36) begin
      if (_T_23) begin
        state <= 3'h4;
      end else if (_T_47) begin
        state <= 3'h1;
      end else if (_T_58) begin
        state <= 3'h2;
      end
    end else if (_T_61) begin
      if (io_lastOut) begin
        state <= 3'h0;
      end
    end
    if (reset) begin
      statePrev <= 3'h0;
    end else begin
      statePrev <= state;
    end
    if (reset) begin
      last <= 1'h0;
    end else if (_T_3) begin
      last <= 1'h0;
    end else if (!(_T_7)) begin
      if (_T_21) begin
        if (_T_23) begin
          last <= _GEN_3;
        end
      end
    end
    if (reset) begin
      doNotScale <= 1'h0;
    end else if (_T_88) begin
      doNotScale <= 1'h0;
    end else begin
      doNotScale <= _GEN_19;
    end
    _T_232 <= cntAcc;
    _T_236 <= _T_62 | _T_63;
    if (_T_116) begin
      _T_239 <= _T_101;
    end else begin
      _T_239 <= cntLoad;
    end
  end
endmodule
module AXI4AccumulatorBlock(
  input         clock,
  input         reset,
  output        auto_mem_in_aw_ready,
  input         auto_mem_in_aw_valid,
  input         auto_mem_in_aw_bits_id,
  input  [29:0] auto_mem_in_aw_bits_addr,
  output        auto_mem_in_w_ready,
  input         auto_mem_in_w_valid,
  input  [31:0] auto_mem_in_w_bits_data,
  input  [3:0]  auto_mem_in_w_bits_strb,
  input         auto_mem_in_b_ready,
  output        auto_mem_in_b_valid,
  output        auto_mem_in_b_bits_id,
  output        auto_mem_in_ar_ready,
  input         auto_mem_in_ar_valid,
  input         auto_mem_in_ar_bits_id,
  input  [29:0] auto_mem_in_ar_bits_addr,
  input  [2:0]  auto_mem_in_ar_bits_size,
  input         auto_mem_in_r_ready,
  output        auto_mem_in_r_valid,
  output        auto_mem_in_r_bits_id,
  output [31:0] auto_mem_in_r_bits_data,
  input         auto_master_out_ready,
  output        auto_master_out_valid,
  output [15:0] auto_master_out_bits_data,
  output        auto_master_out_bits_last,
  output        auto_slave_in_ready,
  input         auto_slave_in_valid,
  input  [31:0] auto_slave_in_bits_data,
  input         auto_slave_in_bits_last
);
  wire  acc_clock; // @[AccDspBlock.scala 39:21]
  wire  acc_reset; // @[AccDspBlock.scala 39:21]
  wire  acc_io_in_ready; // @[AccDspBlock.scala 39:21]
  wire  acc_io_in_valid; // @[AccDspBlock.scala 39:21]
  wire [15:0] acc_io_in_bits; // @[AccDspBlock.scala 39:21]
  wire  acc_io_lastIn; // @[AccDspBlock.scala 39:21]
  wire [7:0] acc_io_accDepthReg; // @[AccDspBlock.scala 39:21]
  wire [16:0] acc_io_accWindowsReg; // @[AccDspBlock.scala 39:21]
  wire  acc_io_out_ready; // @[AccDspBlock.scala 39:21]
  wire  acc_io_out_valid; // @[AccDspBlock.scala 39:21]
  wire [15:0] acc_io_out_bits; // @[AccDspBlock.scala 39:21]
  wire  acc_io_lastOut; // @[AccDspBlock.scala 39:21]
  wire  Queue_clock; // @[Decoupled.scala 296:21]
  wire  Queue_reset; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_bits_read; // @[Decoupled.scala 296:21]
  wire [31:0] Queue_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_bits_extra; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_bits_read; // @[Decoupled.scala 296:21]
  wire [31:0] Queue_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_bits_extra; // @[Decoupled.scala 296:21]
  reg [7:0] accDepth; // @[AccDspBlock.scala 42:34]
  reg [31:0] _RAND_0;
  reg [16:0] numWin; // @[AccDspBlock.scala 43:34]
  reg [31:0] _RAND_1;
  wire  _T_2 = auto_mem_in_aw_valid & auto_mem_in_w_valid; // @[RegisterRouter.scala 40:39]
  wire  _T_3 = auto_mem_in_ar_valid | _T_2; // @[RegisterRouter.scala 40:26]
  wire  _T_4 = ~auto_mem_in_ar_valid; // @[RegisterRouter.scala 42:29]
  wire  _T_47_ready = Queue_io_enq_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 299:17]
  wire [29:0] _T_11 = auto_mem_in_ar_valid ? auto_mem_in_ar_bits_addr : auto_mem_in_aw_bits_addr; // @[RegisterRouter.scala 48:19]
  wire [1:0] _T_51 = _T_11[3:2] & 2'h2; // @[RegisterRouter.scala 59:16]
  wire  _T_53 = _T_51 == 2'h0; // @[RegisterRouter.scala 59:16]
  wire  _T_5 = _T_47_ready & _T_4; // @[RegisterRouter.scala 42:26]
  wire [1:0] _T_14 = 2'h1 << auto_mem_in_ar_bits_size[0]; // @[OneHot.scala 65:12]
  wire [1:0] _T_16 = _T_14 | 2'h1; // @[Misc.scala 200:81]
  wire  _T_17 = auto_mem_in_ar_bits_size >= 3'h2; // @[Misc.scala 204:21]
  wire  _T_20 = ~auto_mem_in_ar_bits_addr[1]; // @[Misc.scala 209:20]
  wire  _T_22 = _T_16[1] & _T_20; // @[Misc.scala 213:38]
  wire  _T_23 = _T_17 | _T_22; // @[Misc.scala 213:29]
  wire  _T_25 = _T_16[1] & auto_mem_in_ar_bits_addr[1]; // @[Misc.scala 213:38]
  wire  _T_26 = _T_17 | _T_25; // @[Misc.scala 213:29]
  wire  _T_29 = ~auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 209:20]
  wire  _T_30 = _T_20 & _T_29; // @[Misc.scala 212:27]
  wire  _T_31 = _T_16[0] & _T_30; // @[Misc.scala 213:38]
  wire  _T_32 = _T_23 | _T_31; // @[Misc.scala 213:29]
  wire  _T_33 = _T_20 & auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  wire  _T_34 = _T_16[0] & _T_33; // @[Misc.scala 213:38]
  wire  _T_35 = _T_23 | _T_34; // @[Misc.scala 213:29]
  wire  _T_36 = auto_mem_in_ar_bits_addr[1] & _T_29; // @[Misc.scala 212:27]
  wire  _T_37 = _T_16[0] & _T_36; // @[Misc.scala 213:38]
  wire  _T_38 = _T_26 | _T_37; // @[Misc.scala 213:29]
  wire  _T_39 = auto_mem_in_ar_bits_addr[1] & auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  wire  _T_40 = _T_16[0] & _T_39; // @[Misc.scala 213:38]
  wire  _T_41 = _T_26 | _T_40; // @[Misc.scala 213:29]
  wire [3:0] _T_44 = {_T_41,_T_38,_T_35,_T_32}; // @[Cat.scala 29:58]
  wire [3:0] _T_46 = auto_mem_in_ar_valid ? _T_44 : auto_mem_in_w_bits_strb; // @[RegisterRouter.scala 54:25]
  wire [7:0] _T_65 = _T_46[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_67 = _T_46[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_69 = _T_46[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_71 = _T_46[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_74 = {_T_71,_T_69,_T_67,_T_65}; // @[Cat.scala 29:58]
  wire  _T_93 = _T_74[16:0] == 17'h1ffff; // @[RegisterRouter.scala 59:16]
  wire  _T_146 = _T_3 & _T_47_ready; // @[RegisterRouter.scala 59:16]
  wire [1:0] _T_140 = 2'h1 << _T_11[2]; // @[OneHot.scala 58:35]
  wire  _T_163 = _T_146 & _T_4; // @[RegisterRouter.scala 59:16]
  wire  _T_170 = _T_163 & _T_140[1]; // @[RegisterRouter.scala 59:16]
  wire  _T_171 = _T_170 & _T_53; // @[RegisterRouter.scala 59:16]
  wire  _T_100 = _T_171 & _T_93; // @[RegisterRouter.scala 59:16]
  wire  _T_116 = _T_74[7:0] == 8'hff; // @[RegisterRouter.scala 59:16]
  wire  _T_165 = _T_163 & _T_140[0]; // @[RegisterRouter.scala 59:16]
  wire  _T_166 = _T_165 & _T_53; // @[RegisterRouter.scala 59:16]
  wire  _T_123 = _T_166 & _T_116; // @[RegisterRouter.scala 59:16]
  wire  _GEN_11 = _T_11[2] ? _T_53 : _T_53; // @[MuxLiteral.scala 48:10]
  wire [16:0] _T_218_0 = {{9'd0}, accDepth}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [16:0] _GEN_13 = _T_11[2] ? numWin : _T_218_0; // @[MuxLiteral.scala 48:10]
  wire [16:0] _T_220 = _GEN_11 ? _GEN_13 : 17'h0; // @[RegisterRouter.scala 59:16]
  wire  _T_221_bits_read = Queue_io_deq_bits_read; // @[Decoupled.scala 317:19 Decoupled.scala 318:14]
  wire  _T_221_valid = Queue_io_deq_valid; // @[Decoupled.scala 317:19 Decoupled.scala 319:15]
  wire  _T_224 = ~_T_221_bits_read; // @[RegisterRouter.scala 65:29]
  wire [31:0] _T_228 = auto_slave_in_bits_data; // @[AccDspBlock.scala 63:48]
  Accumulator acc ( // @[AccDspBlock.scala 39:21]
    .clock(acc_clock),
    .reset(acc_reset),
    .io_in_ready(acc_io_in_ready),
    .io_in_valid(acc_io_in_valid),
    .io_in_bits(acc_io_in_bits),
    .io_lastIn(acc_io_lastIn),
    .io_accDepthReg(acc_io_accDepthReg),
    .io_accWindowsReg(acc_io_accWindowsReg),
    .io_out_ready(acc_io_out_ready),
    .io_out_valid(acc_io_out_valid),
    .io_out_bits(acc_io_out_bits),
    .io_lastOut(acc_io_lastOut)
  );
  Queue Queue ( // @[Decoupled.scala 296:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_read(Queue_io_enq_bits_read),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_extra(Queue_io_enq_bits_extra),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_read(Queue_io_deq_bits_read),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_extra(Queue_io_deq_bits_extra)
  );
  assign auto_mem_in_aw_ready = _T_5 & auto_mem_in_w_valid; // @[LazyModule.scala 173:31]
  assign auto_mem_in_w_ready = _T_5 & auto_mem_in_aw_valid; // @[LazyModule.scala 173:31]
  assign auto_mem_in_b_valid = _T_221_valid & _T_224; // @[LazyModule.scala 173:31]
  assign auto_mem_in_b_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_mem_in_ar_ready = Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_valid = _T_221_valid & _T_221_bits_read; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 173:31]
  assign auto_master_out_valid = acc_io_out_valid; // @[LazyModule.scala 173:49]
  assign auto_master_out_bits_data = acc_io_out_bits; // @[LazyModule.scala 173:49]
  assign auto_master_out_bits_last = acc_io_lastOut; // @[LazyModule.scala 173:49]
  assign auto_slave_in_ready = acc_io_in_ready; // @[LazyModule.scala 173:31]
  assign acc_clock = clock;
  assign acc_reset = reset;
  assign acc_io_in_valid = auto_slave_in_valid; // @[AccDspBlock.scala 61:24]
  assign acc_io_in_bits = _T_228[15:0]; // @[AccDspBlock.scala 63:24]
  assign acc_io_lastIn = auto_slave_in_bits_last; // @[AccDspBlock.scala 66:24]
  assign acc_io_accDepthReg = accDepth; // @[AccDspBlock.scala 45:26]
  assign acc_io_accWindowsReg = numWin; // @[AccDspBlock.scala 46:26]
  assign acc_io_out_ready = auto_master_out_ready; // @[AccDspBlock.scala 70:22]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_mem_in_ar_valid | _T_2; // @[Decoupled.scala 297:22]
  assign Queue_io_enq_bits_read = auto_mem_in_ar_valid; // @[Decoupled.scala 298:21]
  assign Queue_io_enq_bits_data = {{15'd0}, _T_220}; // @[Decoupled.scala 298:21]
  assign Queue_io_enq_bits_extra = auto_mem_in_ar_valid ? auto_mem_in_ar_bits_id : auto_mem_in_aw_bits_id; // @[Decoupled.scala 298:21]
  assign Queue_io_deq_ready = _T_221_bits_read ? auto_mem_in_r_ready : auto_mem_in_b_ready; // @[Decoupled.scala 320:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  accDepth = _RAND_0[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  numWin = _RAND_1[16:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      accDepth <= 8'h80;
    end else if (_T_123) begin
      accDepth <= auto_mem_in_w_bits_data[7:0];
    end
    if (reset) begin
      numWin <= 17'h10000;
    end else if (_T_100) begin
      numWin <= auto_mem_in_w_bits_data[16:0];
    end
  end
endmodule
module Queue_22(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [15:0] io_enq_bits_data,
  input         io_enq_bits_last,
  input         io_deq_ready,
  output        io_deq_valid,
  output [15:0] io_deq_bits_data,
  output        io_deq_bits_last
);
  reg [15:0] _T_data [0:127]; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_0;
  wire [15:0] _T_data__T_18_data; // @[Decoupled.scala 218:24]
  wire [6:0] _T_data__T_18_addr; // @[Decoupled.scala 218:24]
  wire [15:0] _T_data__T_10_data; // @[Decoupled.scala 218:24]
  wire [6:0] _T_data__T_10_addr; // @[Decoupled.scala 218:24]
  wire  _T_data__T_10_mask; // @[Decoupled.scala 218:24]
  wire  _T_data__T_10_en; // @[Decoupled.scala 218:24]
  reg  _T_last [0:127]; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_1;
  wire  _T_last__T_18_data; // @[Decoupled.scala 218:24]
  wire [6:0] _T_last__T_18_addr; // @[Decoupled.scala 218:24]
  wire  _T_last__T_10_data; // @[Decoupled.scala 218:24]
  wire [6:0] _T_last__T_10_addr; // @[Decoupled.scala 218:24]
  wire  _T_last__T_10_mask; // @[Decoupled.scala 218:24]
  wire  _T_last__T_10_en; // @[Decoupled.scala 218:24]
  reg [6:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_2;
  reg [6:0] value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_3;
  reg  _T_1; // @[Decoupled.scala 221:35]
  reg [31:0] _RAND_4;
  wire  _T_2 = value == value_1; // @[Decoupled.scala 223:41]
  wire  _T_3 = ~_T_1; // @[Decoupled.scala 224:36]
  wire  _T_4 = _T_2 & _T_3; // @[Decoupled.scala 224:33]
  wire  _T_5 = _T_2 & _T_1; // @[Decoupled.scala 225:32]
  wire  _T_6 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  _T_8 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire [6:0] _T_12 = value + 7'h1; // @[Counter.scala 39:22]
  wire [6:0] _T_14 = value_1 + 7'h1; // @[Counter.scala 39:22]
  wire  _T_15 = _T_6 != _T_8; // @[Decoupled.scala 236:16]
  assign _T_data__T_18_addr = value_1;
  assign _T_data__T_18_data = _T_data[_T_data__T_18_addr]; // @[Decoupled.scala 218:24]
  assign _T_data__T_10_data = io_enq_bits_data;
  assign _T_data__T_10_addr = value;
  assign _T_data__T_10_mask = 1'h1;
  assign _T_data__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_last__T_18_addr = value_1;
  assign _T_last__T_18_data = _T_last[_T_last__T_18_addr]; // @[Decoupled.scala 218:24]
  assign _T_last__T_10_data = io_enq_bits_last;
  assign _T_last__T_10_addr = value;
  assign _T_last__T_10_mask = 1'h1;
  assign _T_last__T_10_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~_T_5; // @[Decoupled.scala 241:16]
  assign io_deq_valid = ~_T_4; // @[Decoupled.scala 240:16]
  assign io_deq_bits_data = _T_data__T_18_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_last = _T_last__T_18_data; // @[Decoupled.scala 242:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    _T_data[initvar] = _RAND_0[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    _T_last[initvar] = _RAND_1[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  value = _RAND_2[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  value_1 = _RAND_3[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T_data__T_10_en & _T_data__T_10_mask) begin
      _T_data[_T_data__T_10_addr] <= _T_data__T_10_data; // @[Decoupled.scala 218:24]
    end
    if(_T_last__T_10_en & _T_last__T_10_mask) begin
      _T_last[_T_last__T_10_addr] <= _T_last__T_10_data; // @[Decoupled.scala 218:24]
    end
    if (reset) begin
      value <= 7'h0;
    end else if (_T_6) begin
      value <= _T_12;
    end
    if (reset) begin
      value_1 <= 7'h0;
    end else if (_T_8) begin
      value_1 <= _T_14;
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else if (_T_15) begin
      _T_1 <= _T_6;
    end
  end
endmodule
module Queue_23(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input         io_enq_bits_read,
  input  [9:0]  io_enq_bits_index,
  input  [31:0] io_enq_bits_data,
  input  [3:0]  io_enq_bits_mask,
  input         io_enq_bits_extra,
  input         io_deq_ready,
  output        io_deq_valid,
  output        io_deq_bits_read,
  output [9:0]  io_deq_bits_index,
  output [31:0] io_deq_bits_data,
  output [3:0]  io_deq_bits_mask,
  output        io_deq_bits_extra
);
  reg  _T_read [0:3]; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_0;
  wire  _T_read__T_18_data; // @[Decoupled.scala 218:24]
  wire [1:0] _T_read__T_18_addr; // @[Decoupled.scala 218:24]
  wire  _T_read__T_10_data; // @[Decoupled.scala 218:24]
  wire [1:0] _T_read__T_10_addr; // @[Decoupled.scala 218:24]
  wire  _T_read__T_10_mask; // @[Decoupled.scala 218:24]
  wire  _T_read__T_10_en; // @[Decoupled.scala 218:24]
  reg [9:0] _T_index [0:3]; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_1;
  wire [9:0] _T_index__T_18_data; // @[Decoupled.scala 218:24]
  wire [1:0] _T_index__T_18_addr; // @[Decoupled.scala 218:24]
  wire [9:0] _T_index__T_10_data; // @[Decoupled.scala 218:24]
  wire [1:0] _T_index__T_10_addr; // @[Decoupled.scala 218:24]
  wire  _T_index__T_10_mask; // @[Decoupled.scala 218:24]
  wire  _T_index__T_10_en; // @[Decoupled.scala 218:24]
  reg [31:0] _T_data [0:3]; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_2;
  wire [31:0] _T_data__T_18_data; // @[Decoupled.scala 218:24]
  wire [1:0] _T_data__T_18_addr; // @[Decoupled.scala 218:24]
  wire [31:0] _T_data__T_10_data; // @[Decoupled.scala 218:24]
  wire [1:0] _T_data__T_10_addr; // @[Decoupled.scala 218:24]
  wire  _T_data__T_10_mask; // @[Decoupled.scala 218:24]
  wire  _T_data__T_10_en; // @[Decoupled.scala 218:24]
  reg [3:0] _T_mask [0:3]; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_3;
  wire [3:0] _T_mask__T_18_data; // @[Decoupled.scala 218:24]
  wire [1:0] _T_mask__T_18_addr; // @[Decoupled.scala 218:24]
  wire [3:0] _T_mask__T_10_data; // @[Decoupled.scala 218:24]
  wire [1:0] _T_mask__T_10_addr; // @[Decoupled.scala 218:24]
  wire  _T_mask__T_10_mask; // @[Decoupled.scala 218:24]
  wire  _T_mask__T_10_en; // @[Decoupled.scala 218:24]
  reg  _T_extra [0:3]; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_4;
  wire  _T_extra__T_18_data; // @[Decoupled.scala 218:24]
  wire [1:0] _T_extra__T_18_addr; // @[Decoupled.scala 218:24]
  wire  _T_extra__T_10_data; // @[Decoupled.scala 218:24]
  wire [1:0] _T_extra__T_10_addr; // @[Decoupled.scala 218:24]
  wire  _T_extra__T_10_mask; // @[Decoupled.scala 218:24]
  wire  _T_extra__T_10_en; // @[Decoupled.scala 218:24]
  reg [1:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  reg [1:0] value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_6;
  reg  _T_1; // @[Decoupled.scala 221:35]
  reg [31:0] _RAND_7;
  wire  _T_2 = value == value_1; // @[Decoupled.scala 223:41]
  wire  _T_3 = ~_T_1; // @[Decoupled.scala 224:36]
  wire  _T_4 = _T_2 & _T_3; // @[Decoupled.scala 224:33]
  wire  _T_5 = _T_2 & _T_1; // @[Decoupled.scala 225:32]
  wire  _T_6 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  _T_8 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire [1:0] _T_12 = value + 2'h1; // @[Counter.scala 39:22]
  wire [1:0] _T_14 = value_1 + 2'h1; // @[Counter.scala 39:22]
  wire  _T_15 = _T_6 != _T_8; // @[Decoupled.scala 236:16]
  assign _T_read__T_18_addr = value_1;
  assign _T_read__T_18_data = _T_read[_T_read__T_18_addr]; // @[Decoupled.scala 218:24]
  assign _T_read__T_10_data = io_enq_bits_read;
  assign _T_read__T_10_addr = value;
  assign _T_read__T_10_mask = 1'h1;
  assign _T_read__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_index__T_18_addr = value_1;
  assign _T_index__T_18_data = _T_index[_T_index__T_18_addr]; // @[Decoupled.scala 218:24]
  assign _T_index__T_10_data = io_enq_bits_index;
  assign _T_index__T_10_addr = value;
  assign _T_index__T_10_mask = 1'h1;
  assign _T_index__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_data__T_18_addr = value_1;
  assign _T_data__T_18_data = _T_data[_T_data__T_18_addr]; // @[Decoupled.scala 218:24]
  assign _T_data__T_10_data = io_enq_bits_data;
  assign _T_data__T_10_addr = value;
  assign _T_data__T_10_mask = 1'h1;
  assign _T_data__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_mask__T_18_addr = value_1;
  assign _T_mask__T_18_data = _T_mask[_T_mask__T_18_addr]; // @[Decoupled.scala 218:24]
  assign _T_mask__T_10_data = io_enq_bits_mask;
  assign _T_mask__T_10_addr = value;
  assign _T_mask__T_10_mask = 1'h1;
  assign _T_mask__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_extra__T_18_addr = value_1;
  assign _T_extra__T_18_data = _T_extra[_T_extra__T_18_addr]; // @[Decoupled.scala 218:24]
  assign _T_extra__T_10_data = io_enq_bits_extra;
  assign _T_extra__T_10_addr = value;
  assign _T_extra__T_10_mask = 1'h1;
  assign _T_extra__T_10_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~_T_5; // @[Decoupled.scala 241:16]
  assign io_deq_valid = ~_T_4; // @[Decoupled.scala 240:16]
  assign io_deq_bits_read = _T_read__T_18_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_index = _T_index__T_18_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_data = _T_data__T_18_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_mask = _T_mask__T_18_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_extra = _T_extra__T_18_data; // @[Decoupled.scala 242:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    _T_read[initvar] = _RAND_0[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    _T_index[initvar] = _RAND_1[9:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    _T_data[initvar] = _RAND_2[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    _T_mask[initvar] = _RAND_3[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_4 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    _T_extra[initvar] = _RAND_4[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  value_1 = _RAND_6[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_1 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T_read__T_10_en & _T_read__T_10_mask) begin
      _T_read[_T_read__T_10_addr] <= _T_read__T_10_data; // @[Decoupled.scala 218:24]
    end
    if(_T_index__T_10_en & _T_index__T_10_mask) begin
      _T_index[_T_index__T_10_addr] <= _T_index__T_10_data; // @[Decoupled.scala 218:24]
    end
    if(_T_data__T_10_en & _T_data__T_10_mask) begin
      _T_data[_T_data__T_10_addr] <= _T_data__T_10_data; // @[Decoupled.scala 218:24]
    end
    if(_T_mask__T_10_en & _T_mask__T_10_mask) begin
      _T_mask[_T_mask__T_10_addr] <= _T_mask__T_10_data; // @[Decoupled.scala 218:24]
    end
    if(_T_extra__T_10_en & _T_extra__T_10_mask) begin
      _T_extra[_T_extra__T_10_addr] <= _T_extra__T_10_data; // @[Decoupled.scala 218:24]
    end
    if (reset) begin
      value <= 2'h0;
    end else if (_T_6) begin
      value <= _T_12;
    end
    if (reset) begin
      value_1 <= 2'h0;
    end else if (_T_8) begin
      value_1 <= _T_14;
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else if (_T_15) begin
      _T_1 <= _T_6;
    end
  end
endmodule
module AXI4DspQueueBlock(
  input         clock,
  input         reset,
  output        auto_stream_in_ready,
  input         auto_stream_in_valid,
  input  [15:0] auto_stream_in_bits_data,
  input         auto_stream_in_bits_last,
  input         auto_stream_out_ready,
  output        auto_stream_out_valid,
  output [15:0] auto_stream_out_bits_data,
  output        auto_stream_out_bits_last,
  output        auto_in_aw_ready,
  input         auto_in_aw_valid,
  input         auto_in_aw_bits_id,
  input  [29:0] auto_in_aw_bits_addr,
  output        auto_in_w_ready,
  input         auto_in_w_valid,
  input  [31:0] auto_in_w_bits_data,
  input  [3:0]  auto_in_w_bits_strb,
  input         auto_in_b_ready,
  output        auto_in_b_valid,
  output        auto_in_b_bits_id,
  output        auto_in_ar_ready,
  input         auto_in_ar_valid,
  input         auto_in_ar_bits_id,
  input  [29:0] auto_in_ar_bits_addr,
  input  [2:0]  auto_in_ar_bits_size,
  input         auto_in_r_ready,
  output        auto_in_r_valid,
  output        auto_in_r_bits_id,
  output [31:0] auto_in_r_bits_data
);
  wire  queuedStream_clock; // @[Decoupled.scala 296:21]
  wire  queuedStream_reset; // @[Decoupled.scala 296:21]
  wire  queuedStream_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  queuedStream_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [15:0] queuedStream_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire  queuedStream_io_enq_bits_last; // @[Decoupled.scala 296:21]
  wire  queuedStream_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  queuedStream_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [15:0] queuedStream_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire  queuedStream_io_deq_bits_last; // @[Decoupled.scala 296:21]
  wire  Queue_clock; // @[Decoupled.scala 296:21]
  wire  Queue_reset; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_bits_read; // @[Decoupled.scala 296:21]
  wire [9:0] Queue_io_enq_bits_index; // @[Decoupled.scala 296:21]
  wire [31:0] Queue_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire [3:0] Queue_io_enq_bits_mask; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_bits_extra; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_bits_read; // @[Decoupled.scala 296:21]
  wire [9:0] Queue_io_deq_bits_index; // @[Decoupled.scala 296:21]
  wire [31:0] Queue_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire [3:0] Queue_io_deq_bits_mask; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_bits_extra; // @[Decoupled.scala 296:21]
  wire  Queue_1_clock; // @[Decoupled.scala 296:21]
  wire  Queue_1_reset; // @[Decoupled.scala 296:21]
  wire  Queue_1_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  Queue_1_io_enq_valid; // @[Decoupled.scala 296:21]
  wire  Queue_1_io_enq_bits_read; // @[Decoupled.scala 296:21]
  wire [31:0] Queue_1_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire  Queue_1_io_enq_bits_extra; // @[Decoupled.scala 296:21]
  wire  Queue_1_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  Queue_1_io_deq_valid; // @[Decoupled.scala 296:21]
  wire  Queue_1_io_deq_bits_read; // @[Decoupled.scala 296:21]
  wire [31:0] Queue_1_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire  Queue_1_io_deq_bits_extra; // @[Decoupled.scala 296:21]
  wire  _T_53_ready = Queue_1_io_enq_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 299:17]
  wire  _T_154 = Queue_io_deq_valid & _T_53_ready; // @[RegisterRouter.scala 59:16]
  wire  _T_155 = ~Queue_io_deq_bits_read; // @[RegisterRouter.scala 59:16]
  wire  _T_156 = _T_154 & _T_155; // @[RegisterRouter.scala 59:16]
  wire [9:0] _T_57 = Queue_io_deq_bits_index; // @[RegisterRouter.scala 59:16]
  wire  _T_59 = _T_57 == 10'h0; // @[RegisterRouter.scala 59:16]
  wire  _T_159 = _T_156 & _T_59; // @[RegisterRouter.scala 59:16]
  wire [7:0] _T_90 = Queue_io_deq_bits_mask[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_88 = Queue_io_deq_bits_mask[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_86 = Queue_io_deq_bits_mask[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_84 = Queue_io_deq_bits_mask[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_93 = {_T_90,_T_88,_T_86,_T_84}; // @[Cat.scala 29:58]
  wire  _T_101 = _T_93 == 32'hffffffff; // @[RegisterRouter.scala 59:16]
  wire  _T_105 = _T_159 & _T_101; // @[RegisterRouter.scala 59:16]
  wire [31:0] _T_106 = Queue_io_deq_bits_data; // @[RegisterRouter.scala 59:16]
  wire [31:0] queueThreshold = _T_105 ? _T_106 : 32'h80; // @[RegField.scala 134:88]
  wire  _T_8 = auto_in_aw_valid & auto_in_w_valid; // @[RegisterRouter.scala 40:39]
  wire  _T_10 = ~auto_in_ar_valid; // @[RegisterRouter.scala 42:29]
  wire  _T_54_ready = Queue_io_enq_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 299:17]
  wire [29:0] _T_17 = auto_in_ar_valid ? auto_in_ar_bits_addr : auto_in_aw_bits_addr; // @[RegisterRouter.scala 48:19]
  wire  _T_11 = _T_54_ready & _T_10; // @[RegisterRouter.scala 42:26]
  wire [1:0] _T_20 = 2'h1 << auto_in_ar_bits_size[0]; // @[OneHot.scala 65:12]
  wire [1:0] _T_22 = _T_20 | 2'h1; // @[Misc.scala 200:81]
  wire  _T_23 = auto_in_ar_bits_size >= 3'h2; // @[Misc.scala 204:21]
  wire  _T_26 = ~auto_in_ar_bits_addr[1]; // @[Misc.scala 209:20]
  wire  _T_28 = _T_22[1] & _T_26; // @[Misc.scala 213:38]
  wire  _T_29 = _T_23 | _T_28; // @[Misc.scala 213:29]
  wire  _T_31 = _T_22[1] & auto_in_ar_bits_addr[1]; // @[Misc.scala 213:38]
  wire  _T_32 = _T_23 | _T_31; // @[Misc.scala 213:29]
  wire  _T_35 = ~auto_in_ar_bits_addr[0]; // @[Misc.scala 209:20]
  wire  _T_36 = _T_26 & _T_35; // @[Misc.scala 212:27]
  wire  _T_37 = _T_22[0] & _T_36; // @[Misc.scala 213:38]
  wire  _T_38 = _T_29 | _T_37; // @[Misc.scala 213:29]
  wire  _T_39 = _T_26 & auto_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  wire  _T_40 = _T_22[0] & _T_39; // @[Misc.scala 213:38]
  wire  _T_41 = _T_29 | _T_40; // @[Misc.scala 213:29]
  wire  _T_42 = auto_in_ar_bits_addr[1] & _T_35; // @[Misc.scala 212:27]
  wire  _T_43 = _T_22[0] & _T_42; // @[Misc.scala 213:38]
  wire  _T_44 = _T_32 | _T_43; // @[Misc.scala 213:29]
  wire  _T_45 = auto_in_ar_bits_addr[1] & auto_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  wire  _T_46 = _T_22[0] & _T_45; // @[Misc.scala 213:38]
  wire  _T_47 = _T_32 | _T_46; // @[Misc.scala 213:29]
  wire [3:0] _T_50 = {_T_47,_T_44,_T_41,_T_38}; // @[Cat.scala 29:58]
  wire  _T_178_bits_read = Queue_1_io_deq_bits_read; // @[Decoupled.scala 317:19 Decoupled.scala 318:14]
  wire  _T_178_valid = Queue_1_io_deq_valid; // @[Decoupled.scala 317:19 Decoupled.scala 319:15]
  wire  _T_181 = ~_T_178_bits_read; // @[RegisterRouter.scala 65:29]
  Queue_22 queuedStream ( // @[Decoupled.scala 296:21]
    .clock(queuedStream_clock),
    .reset(queuedStream_reset),
    .io_enq_ready(queuedStream_io_enq_ready),
    .io_enq_valid(queuedStream_io_enq_valid),
    .io_enq_bits_data(queuedStream_io_enq_bits_data),
    .io_enq_bits_last(queuedStream_io_enq_bits_last),
    .io_deq_ready(queuedStream_io_deq_ready),
    .io_deq_valid(queuedStream_io_deq_valid),
    .io_deq_bits_data(queuedStream_io_deq_bits_data),
    .io_deq_bits_last(queuedStream_io_deq_bits_last)
  );
  Queue_23 Queue ( // @[Decoupled.scala 296:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_read(Queue_io_enq_bits_read),
    .io_enq_bits_index(Queue_io_enq_bits_index),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_mask(Queue_io_enq_bits_mask),
    .io_enq_bits_extra(Queue_io_enq_bits_extra),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_read(Queue_io_deq_bits_read),
    .io_deq_bits_index(Queue_io_deq_bits_index),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_mask(Queue_io_deq_bits_mask),
    .io_deq_bits_extra(Queue_io_deq_bits_extra)
  );
  Queue Queue_1 ( // @[Decoupled.scala 296:21]
    .clock(Queue_1_clock),
    .reset(Queue_1_reset),
    .io_enq_ready(Queue_1_io_enq_ready),
    .io_enq_valid(Queue_1_io_enq_valid),
    .io_enq_bits_read(Queue_1_io_enq_bits_read),
    .io_enq_bits_data(Queue_1_io_enq_bits_data),
    .io_enq_bits_extra(Queue_1_io_enq_bits_extra),
    .io_deq_ready(Queue_1_io_deq_ready),
    .io_deq_valid(Queue_1_io_deq_valid),
    .io_deq_bits_read(Queue_1_io_deq_bits_read),
    .io_deq_bits_data(Queue_1_io_deq_bits_data),
    .io_deq_bits_extra(Queue_1_io_deq_bits_extra)
  );
  assign auto_stream_in_ready = queuedStream_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_stream_out_valid = queuedStream_io_deq_valid; // @[LazyModule.scala 173:49]
  assign auto_stream_out_bits_data = queuedStream_io_deq_bits_data; // @[LazyModule.scala 173:49]
  assign auto_stream_out_bits_last = queuedStream_io_deq_bits_last; // @[LazyModule.scala 173:49]
  assign auto_in_aw_ready = _T_11 & auto_in_w_valid; // @[LazyModule.scala 173:31]
  assign auto_in_w_ready = _T_11 & auto_in_aw_valid; // @[LazyModule.scala 173:31]
  assign auto_in_b_valid = _T_178_valid & _T_181; // @[LazyModule.scala 173:31]
  assign auto_in_b_bits_id = Queue_1_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_in_ar_ready = Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_in_r_valid = _T_178_valid & _T_178_bits_read; // @[LazyModule.scala 173:31]
  assign auto_in_r_bits_id = Queue_1_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_in_r_bits_data = Queue_1_io_deq_bits_data; // @[LazyModule.scala 173:31]
  assign queuedStream_clock = clock;
  assign queuedStream_reset = reset;
  assign queuedStream_io_enq_valid = auto_stream_in_valid; // @[Decoupled.scala 297:22]
  assign queuedStream_io_enq_bits_data = auto_stream_in_bits_data; // @[Decoupled.scala 298:21]
  assign queuedStream_io_enq_bits_last = auto_stream_in_bits_last; // @[Decoupled.scala 298:21]
  assign queuedStream_io_deq_ready = auto_stream_out_ready; // @[DspQueueBlock.scala 25:13]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_in_ar_valid | _T_8; // @[Decoupled.scala 297:22]
  assign Queue_io_enq_bits_read = auto_in_ar_valid; // @[Decoupled.scala 298:21]
  assign Queue_io_enq_bits_index = _T_17[11:2]; // @[Decoupled.scala 298:21]
  assign Queue_io_enq_bits_data = auto_in_w_bits_data; // @[Decoupled.scala 298:21]
  assign Queue_io_enq_bits_mask = auto_in_ar_valid ? _T_50 : auto_in_w_bits_strb; // @[Decoupled.scala 298:21]
  assign Queue_io_enq_bits_extra = auto_in_ar_valid ? auto_in_ar_bits_id : auto_in_aw_bits_id; // @[Decoupled.scala 298:21]
  assign Queue_io_deq_ready = Queue_1_io_enq_ready; // @[RegisterRouter.scala 59:16]
  assign Queue_1_clock = clock;
  assign Queue_1_reset = reset;
  assign Queue_1_io_enq_valid = Queue_io_deq_valid; // @[Decoupled.scala 297:22]
  assign Queue_1_io_enq_bits_read = Queue_io_deq_bits_read; // @[Decoupled.scala 298:21]
  assign Queue_1_io_enq_bits_data = _T_59 ? queueThreshold : 32'h0; // @[Decoupled.scala 298:21]
  assign Queue_1_io_enq_bits_extra = Queue_io_deq_bits_extra; // @[Decoupled.scala 298:21]
  assign Queue_1_io_deq_ready = _T_178_bits_read ? auto_in_r_ready : auto_in_b_ready; // @[Decoupled.scala 320:15]
endmodule
module AXI4Xbar_1(
  input         clock,
  input         reset,
  output        auto_in_aw_ready,
  input         auto_in_aw_valid,
  input         auto_in_aw_bits_id,
  input  [29:0] auto_in_aw_bits_addr,
  input  [2:0]  auto_in_aw_bits_size,
  output        auto_in_w_ready,
  input         auto_in_w_valid,
  input  [31:0] auto_in_w_bits_data,
  input  [3:0]  auto_in_w_bits_strb,
  input         auto_in_w_bits_last,
  input         auto_in_b_ready,
  output        auto_in_b_valid,
  output [1:0]  auto_in_b_bits_resp,
  output        auto_in_ar_ready,
  input         auto_in_ar_valid,
  input         auto_in_ar_bits_id,
  input  [29:0] auto_in_ar_bits_addr,
  input  [2:0]  auto_in_ar_bits_size,
  input         auto_in_r_ready,
  output        auto_in_r_valid,
  output [31:0] auto_in_r_bits_data,
  output [1:0]  auto_in_r_bits_resp,
  output        auto_in_r_bits_last,
  input         auto_out_1_aw_ready,
  output        auto_out_1_aw_valid,
  output        auto_out_1_aw_bits_id,
  output [29:0] auto_out_1_aw_bits_addr,
  output [2:0]  auto_out_1_aw_bits_size,
  input         auto_out_1_w_ready,
  output        auto_out_1_w_valid,
  output [31:0] auto_out_1_w_bits_data,
  output [3:0]  auto_out_1_w_bits_strb,
  output        auto_out_1_w_bits_last,
  output        auto_out_1_b_ready,
  input         auto_out_1_b_valid,
  input         auto_out_1_b_bits_id,
  input  [1:0]  auto_out_1_b_bits_resp,
  input         auto_out_1_ar_ready,
  output        auto_out_1_ar_valid,
  output        auto_out_1_ar_bits_id,
  output [29:0] auto_out_1_ar_bits_addr,
  output [2:0]  auto_out_1_ar_bits_size,
  output        auto_out_1_r_ready,
  input         auto_out_1_r_valid,
  input         auto_out_1_r_bits_id,
  input  [31:0] auto_out_1_r_bits_data,
  input  [1:0]  auto_out_1_r_bits_resp,
  input         auto_out_1_r_bits_last,
  input         auto_out_0_aw_ready,
  output        auto_out_0_aw_valid,
  output        auto_out_0_aw_bits_id,
  output [29:0] auto_out_0_aw_bits_addr,
  output [2:0]  auto_out_0_aw_bits_size,
  input         auto_out_0_w_ready,
  output        auto_out_0_w_valid,
  output [31:0] auto_out_0_w_bits_data,
  output [3:0]  auto_out_0_w_bits_strb,
  output        auto_out_0_w_bits_last,
  output        auto_out_0_b_ready,
  input         auto_out_0_b_valid,
  input         auto_out_0_b_bits_id,
  input  [1:0]  auto_out_0_b_bits_resp,
  input         auto_out_0_ar_ready,
  output        auto_out_0_ar_valid,
  output        auto_out_0_ar_bits_id,
  output [29:0] auto_out_0_ar_bits_addr,
  output [2:0]  auto_out_0_ar_bits_size,
  output        auto_out_0_r_ready,
  input         auto_out_0_r_valid,
  input         auto_out_0_r_bits_id,
  input  [31:0] auto_out_0_r_bits_data,
  input  [1:0]  auto_out_0_r_bits_resp,
  input         auto_out_0_r_bits_last
);
  wire  awIn_0_clock; // @[Xbar.scala 55:47]
  wire  awIn_0_reset; // @[Xbar.scala 55:47]
  wire  awIn_0_io_enq_ready; // @[Xbar.scala 55:47]
  wire  awIn_0_io_enq_valid; // @[Xbar.scala 55:47]
  wire [1:0] awIn_0_io_enq_bits; // @[Xbar.scala 55:47]
  wire  awIn_0_io_deq_ready; // @[Xbar.scala 55:47]
  wire  awIn_0_io_deq_valid; // @[Xbar.scala 55:47]
  wire [1:0] awIn_0_io_deq_bits; // @[Xbar.scala 55:47]
  wire [30:0] _T_1 = {1'b0,$signed(auto_in_ar_bits_addr)}; // @[Parameters.scala 137:49]
  wire [30:0] _T_3 = $signed(_T_1) & 31'sh1000; // @[Parameters.scala 137:52]
  wire  requestARIO_0_0 = $signed(_T_3) == 31'sh0; // @[Parameters.scala 137:67]
  wire [29:0] _T_5 = auto_in_ar_bits_addr ^ 30'h1000; // @[Parameters.scala 137:31]
  wire [30:0] _T_6 = {1'b0,$signed(_T_5)}; // @[Parameters.scala 137:49]
  wire [30:0] _T_8 = $signed(_T_6) & 31'sh1000; // @[Parameters.scala 137:52]
  wire  requestARIO_0_1 = $signed(_T_8) == 31'sh0; // @[Parameters.scala 137:67]
  wire [30:0] _T_11 = {1'b0,$signed(auto_in_aw_bits_addr)}; // @[Parameters.scala 137:49]
  wire [30:0] _T_13 = $signed(_T_11) & 31'sh1000; // @[Parameters.scala 137:52]
  wire  requestAWIO_0_0 = $signed(_T_13) == 31'sh0; // @[Parameters.scala 137:67]
  wire [29:0] _T_15 = auto_in_aw_bits_addr ^ 30'h1000; // @[Parameters.scala 137:31]
  wire [30:0] _T_16 = {1'b0,$signed(_T_15)}; // @[Parameters.scala 137:49]
  wire [30:0] _T_18 = $signed(_T_16) & 31'sh1000; // @[Parameters.scala 137:52]
  wire  requestAWIO_0_1 = $signed(_T_18) == 31'sh0; // @[Parameters.scala 137:67]
  wire  requestROI_0_0 = ~auto_out_0_r_bits_id; // @[Parameters.scala 47:9]
  wire  requestROI_1_0 = ~auto_out_1_r_bits_id; // @[Parameters.scala 47:9]
  wire  requestBOI_0_0 = ~auto_out_0_b_bits_id; // @[Parameters.scala 47:9]
  wire  requestBOI_1_0 = ~auto_out_1_b_bits_id; // @[Parameters.scala 47:9]
  wire [1:0] _T_20 = {requestAWIO_0_1,requestAWIO_0_0}; // @[Xbar.scala 64:75]
  wire  requestWIO_0_0 = awIn_0_io_deq_bits[0]; // @[Xbar.scala 65:73]
  wire  requestWIO_0_1 = awIn_0_io_deq_bits[1]; // @[Xbar.scala 65:73]
  wire [1:0] _T_27 = {requestARIO_0_1,requestARIO_0_0}; // @[Xbar.scala 93:45]
  wire  _T_108 = requestARIO_0_0 & auto_out_0_ar_ready; // @[Mux.scala 27:72]
  wire  _T_109 = requestARIO_0_1 & auto_out_1_ar_ready; // @[Mux.scala 27:72]
  wire  in_0_ar_ready = _T_108 | _T_109; // @[Mux.scala 27:72]
  reg [2:0] _T_36; // @[Xbar.scala 104:34]
  reg [31:0] _RAND_0;
  wire  _T_55 = _T_36 == 3'h0; // @[Xbar.scala 112:22]
  reg  _T_37; // @[Xbar.scala 105:29]
  reg [31:0] _RAND_1;
  wire  _T_54 = _T_37 == _T_27[1]; // @[Xbar.scala 111:75]
  wire  _T_56 = _T_55 | _T_54; // @[Xbar.scala 112:34]
  wire  _T_57 = _T_36 != 3'h7; // @[Xbar.scala 112:80]
  wire  _T_59 = _T_56 & _T_57; // @[Xbar.scala 112:48]
  wire  io_in_0_ar_ready = in_0_ar_ready & _T_59; // @[Xbar.scala 130:45]
  wire  _T_31 = io_in_0_ar_ready & auto_in_ar_valid; // @[Decoupled.scala 40:37]
  reg  _T_222; // @[Xbar.scala 242:23]
  reg [31:0] _RAND_2;
  wire  _T_127 = auto_out_0_r_valid & requestROI_0_0; // @[Xbar.scala 222:40]
  wire  _T_129 = auto_out_1_r_valid & requestROI_1_0; // @[Xbar.scala 222:40]
  wire  _T_223 = _T_127 | _T_129; // @[Xbar.scala 246:36]
  reg  _T_278_0; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_3;
  wire  _T_284 = _T_278_0 & _T_127; // @[Mux.scala 27:72]
  reg  _T_278_1; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_4;
  wire  _T_285 = _T_278_1 & _T_129; // @[Mux.scala 27:72]
  wire  _T_286 = _T_284 | _T_285; // @[Mux.scala 27:72]
  wire  in_0_r_valid = _T_222 ? _T_223 : _T_286; // @[Xbar.scala 278:22]
  wire  _T_33 = auto_in_r_ready & in_0_r_valid; // @[Decoupled.scala 40:37]
  wire [1:0] _T_224 = {_T_129,_T_127}; // @[Cat.scala 29:58]
  reg [1:0] _T_231; // @[Arbiter.scala 20:23]
  reg [31:0] _RAND_5;
  wire [1:0] _T_232 = ~_T_231; // @[Arbiter.scala 21:30]
  wire [1:0] _T_233 = _T_224 & _T_232; // @[Arbiter.scala 21:28]
  wire [3:0] _T_234 = {_T_233,_T_129,_T_127}; // @[Cat.scala 29:58]
  wire [3:0] _GEN_18 = {{1'd0}, _T_234[3:1]}; // @[package.scala 208:43]
  wire [3:0] _T_236 = _T_234 | _GEN_18; // @[package.scala 208:43]
  wire [3:0] _T_239 = {_T_231, 2'h0}; // @[Arbiter.scala 22:66]
  wire [3:0] _GEN_19 = {{1'd0}, _T_236[3:1]}; // @[Arbiter.scala 22:58]
  wire [3:0] _T_240 = _GEN_19 | _T_239; // @[Arbiter.scala 22:58]
  wire [1:0] _T_243 = _T_240[3:2] & _T_240[1:0]; // @[Arbiter.scala 23:39]
  wire [1:0] _T_244 = ~_T_243; // @[Arbiter.scala 23:18]
  wire  _T_256 = _T_244[0] & _T_127; // @[Xbar.scala 250:63]
  wire  _T_279_0 = _T_222 ? _T_256 : _T_278_0; // @[Xbar.scala 262:23]
  wire [35:0] _T_291 = {auto_out_0_r_bits_id,auto_out_0_r_bits_data,auto_out_0_r_bits_resp,auto_out_0_r_bits_last}; // @[Mux.scala 27:72]
  wire [35:0] _T_292 = _T_279_0 ? _T_291 : 36'h0; // @[Mux.scala 27:72]
  wire  _T_257 = _T_244[1] & _T_129; // @[Xbar.scala 250:63]
  wire  _T_279_1 = _T_222 ? _T_257 : _T_278_1; // @[Xbar.scala 262:23]
  wire [35:0] _T_295 = {auto_out_1_r_bits_id,auto_out_1_r_bits_data,auto_out_1_r_bits_resp,auto_out_1_r_bits_last}; // @[Mux.scala 27:72]
  wire [35:0] _T_296 = _T_279_1 ? _T_295 : 36'h0; // @[Mux.scala 27:72]
  wire [35:0] _T_297 = _T_292 | _T_296; // @[Mux.scala 27:72]
  wire  in_0_r_bits_last = _T_297[0]; // @[Mux.scala 27:72]
  wire  _T_35 = _T_33 & in_0_r_bits_last; // @[Xbar.scala 120:45]
  wire [2:0] _GEN_20 = {{2'd0}, _T_31}; // @[Xbar.scala 106:30]
  wire [2:0] _T_39 = _T_36 + _GEN_20; // @[Xbar.scala 106:30]
  wire [2:0] _GEN_21 = {{2'd0}, _T_35}; // @[Xbar.scala 106:48]
  wire [2:0] _T_41 = _T_39 - _GEN_21; // @[Xbar.scala 106:48]
  wire  _T_42 = ~_T_35; // @[Xbar.scala 107:23]
  wire  _T_43 = _T_36 != 3'h0; // @[Xbar.scala 107:43]
  wire  _T_44 = _T_42 | _T_43; // @[Xbar.scala 107:34]
  wire  _T_46 = _T_44 | reset; // @[Xbar.scala 107:22]
  wire  _T_47 = ~_T_46; // @[Xbar.scala 107:22]
  wire  _T_48 = ~_T_31; // @[Xbar.scala 108:23]
  wire  _T_50 = _T_48 | _T_57; // @[Xbar.scala 108:34]
  wire  _T_52 = _T_50 | reset; // @[Xbar.scala 108:22]
  wire  _T_53 = ~_T_52; // @[Xbar.scala 108:22]
  wire  _T_115 = requestAWIO_0_0 & auto_out_0_aw_ready; // @[Mux.scala 27:72]
  wire  _T_116 = requestAWIO_0_1 & auto_out_1_aw_ready; // @[Mux.scala 27:72]
  wire  in_0_aw_ready = _T_115 | _T_116; // @[Mux.scala 27:72]
  reg  _T_90; // @[Xbar.scala 137:30]
  reg [31:0] _RAND_6;
  wire  _T_94 = _T_90 | awIn_0_io_enq_ready; // @[Xbar.scala 139:57]
  wire  _T_95 = in_0_aw_ready & _T_94; // @[Xbar.scala 139:45]
  reg [2:0] _T_64; // @[Xbar.scala 104:34]
  reg [31:0] _RAND_7;
  wire  _T_83 = _T_64 == 3'h0; // @[Xbar.scala 112:22]
  reg  _T_65; // @[Xbar.scala 105:29]
  reg [31:0] _RAND_8;
  wire  _T_82 = _T_65 == _T_20[1]; // @[Xbar.scala 111:75]
  wire  _T_84 = _T_83 | _T_82; // @[Xbar.scala 112:34]
  wire  _T_85 = _T_64 != 3'h7; // @[Xbar.scala 112:80]
  wire  _T_87 = _T_84 & _T_85; // @[Xbar.scala 112:48]
  wire  io_in_0_aw_ready = _T_95 & _T_87; // @[Xbar.scala 139:82]
  wire  _T_60 = io_in_0_aw_ready & auto_in_aw_valid; // @[Decoupled.scala 40:37]
  reg  _T_304; // @[Xbar.scala 242:23]
  reg [31:0] _RAND_9;
  wire  _T_131 = auto_out_0_b_valid & requestBOI_0_0; // @[Xbar.scala 222:40]
  wire  _T_133 = auto_out_1_b_valid & requestBOI_1_0; // @[Xbar.scala 222:40]
  wire  _T_305 = _T_131 | _T_133; // @[Xbar.scala 246:36]
  reg  _T_360_0; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_10;
  wire  _T_366 = _T_360_0 & _T_131; // @[Mux.scala 27:72]
  reg  _T_360_1; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_11;
  wire  _T_367 = _T_360_1 & _T_133; // @[Mux.scala 27:72]
  wire  _T_368 = _T_366 | _T_367; // @[Mux.scala 27:72]
  wire  in_0_b_valid = _T_304 ? _T_305 : _T_368; // @[Xbar.scala 278:22]
  wire  _T_62 = auto_in_b_ready & in_0_b_valid; // @[Decoupled.scala 40:37]
  wire [2:0] _GEN_22 = {{2'd0}, _T_60}; // @[Xbar.scala 106:30]
  wire [2:0] _T_67 = _T_64 + _GEN_22; // @[Xbar.scala 106:30]
  wire [2:0] _GEN_23 = {{2'd0}, _T_62}; // @[Xbar.scala 106:48]
  wire [2:0] _T_69 = _T_67 - _GEN_23; // @[Xbar.scala 106:48]
  wire  _T_70 = ~_T_62; // @[Xbar.scala 107:23]
  wire  _T_71 = _T_64 != 3'h0; // @[Xbar.scala 107:43]
  wire  _T_72 = _T_70 | _T_71; // @[Xbar.scala 107:34]
  wire  _T_74 = _T_72 | reset; // @[Xbar.scala 107:22]
  wire  _T_75 = ~_T_74; // @[Xbar.scala 107:22]
  wire  _T_76 = ~_T_60; // @[Xbar.scala 108:23]
  wire  _T_78 = _T_76 | _T_85; // @[Xbar.scala 108:34]
  wire  _T_80 = _T_78 | reset; // @[Xbar.scala 108:22]
  wire  _T_81 = ~_T_80; // @[Xbar.scala 108:22]
  wire  in_0_ar_valid = auto_in_ar_valid & _T_59; // @[Xbar.scala 129:45]
  wire  _T_92 = auto_in_aw_valid & _T_94; // @[Xbar.scala 138:45]
  wire  in_0_aw_valid = _T_92 & _T_87; // @[Xbar.scala 138:82]
  wire  _T_97 = ~_T_90; // @[Xbar.scala 140:54]
  wire  _T_99 = awIn_0_io_enq_ready & awIn_0_io_enq_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_2 = _T_99 | _T_90; // @[Xbar.scala 141:38]
  wire  _T_100 = in_0_aw_ready & in_0_aw_valid; // @[Decoupled.scala 40:37]
  wire  in_0_w_valid = auto_in_w_valid & awIn_0_io_deq_valid; // @[Xbar.scala 145:43]
  wire  _T_122 = requestWIO_0_0 & auto_out_0_w_ready; // @[Mux.scala 27:72]
  wire  _T_123 = requestWIO_0_1 & auto_out_1_w_ready; // @[Mux.scala 27:72]
  wire  in_0_w_ready = _T_122 | _T_123; // @[Mux.scala 27:72]
  wire  _T_103 = auto_in_w_valid & auto_in_w_bits_last; // @[Xbar.scala 147:50]
  wire  out_0_ar_valid = in_0_ar_valid & requestARIO_0_0; // @[Xbar.scala 222:40]
  wire  out_1_ar_valid = in_0_ar_valid & requestARIO_0_1; // @[Xbar.scala 222:40]
  wire  out_0_aw_valid = in_0_aw_valid & requestAWIO_0_0; // @[Xbar.scala 222:40]
  wire  out_1_aw_valid = in_0_aw_valid & requestAWIO_0_1; // @[Xbar.scala 222:40]
  wire  _T_140 = ~out_0_aw_valid; // @[Xbar.scala 256:60]
  wire  _T_146 = _T_140 | out_0_aw_valid; // @[Xbar.scala 258:23]
  wire  _T_148 = _T_146 | reset; // @[Xbar.scala 258:12]
  wire  _T_149 = ~_T_148; // @[Xbar.scala 258:12]
  wire  _T_161 = ~out_0_ar_valid; // @[Xbar.scala 256:60]
  wire  _T_167 = _T_161 | out_0_ar_valid; // @[Xbar.scala 258:23]
  wire  _T_169 = _T_167 | reset; // @[Xbar.scala 258:12]
  wire  _T_170 = ~_T_169; // @[Xbar.scala 258:12]
  wire  _T_184 = ~out_1_aw_valid; // @[Xbar.scala 256:60]
  wire  _T_190 = _T_184 | out_1_aw_valid; // @[Xbar.scala 258:23]
  wire  _T_192 = _T_190 | reset; // @[Xbar.scala 258:12]
  wire  _T_193 = ~_T_192; // @[Xbar.scala 258:12]
  wire  _T_205 = ~out_1_ar_valid; // @[Xbar.scala 256:60]
  wire  _T_211 = _T_205 | out_1_ar_valid; // @[Xbar.scala 258:23]
  wire  _T_213 = _T_211 | reset; // @[Xbar.scala 258:12]
  wire  _T_214 = ~_T_213; // @[Xbar.scala 258:12]
  wire  _T_245 = _T_224 != 2'h0; // @[Arbiter.scala 24:27]
  wire  _T_246 = _T_222 & _T_245; // @[Arbiter.scala 24:18]
  wire [1:0] _T_247 = _T_244 & _T_224; // @[Arbiter.scala 25:29]
  wire [2:0] _T_248 = {_T_247, 1'h0}; // @[package.scala 199:48]
  wire [1:0] _T_250 = _T_247 | _T_248[1:0]; // @[package.scala 199:43]
  wire  _T_260 = _T_256 | _T_257; // @[Xbar.scala 255:50]
  wire  _T_262 = ~_T_256; // @[Xbar.scala 256:60]
  wire  _T_265 = ~_T_257; // @[Xbar.scala 256:60]
  wire  _T_266 = _T_262 | _T_265; // @[Xbar.scala 256:57]
  wire  _T_269 = _T_266 | reset; // @[Xbar.scala 256:11]
  wire  _T_270 = ~_T_269; // @[Xbar.scala 256:11]
  wire  _T_271 = ~_T_223; // @[Xbar.scala 258:13]
  wire  _T_273 = _T_271 | _T_260; // @[Xbar.scala 258:23]
  wire  _T_275 = _T_273 | reset; // @[Xbar.scala 258:12]
  wire  _T_276 = ~_T_275; // @[Xbar.scala 258:12]
  wire  _GEN_13 = _T_223 ? 1'h0 : _T_222; // @[Xbar.scala 266:21]
  wire  _GEN_14 = _T_33 | _GEN_13; // @[Xbar.scala 267:24]
  wire  _T_281_0 = _T_222 ? _T_244[0] : _T_278_0; // @[Xbar.scala 270:24]
  wire  _T_281_1 = _T_222 ? _T_244[1] : _T_278_1; // @[Xbar.scala 270:24]
  wire [1:0] _T_306 = {_T_133,_T_131}; // @[Cat.scala 29:58]
  reg [1:0] _T_313; // @[Arbiter.scala 20:23]
  reg [31:0] _RAND_12;
  wire [1:0] _T_314 = ~_T_313; // @[Arbiter.scala 21:30]
  wire [1:0] _T_315 = _T_306 & _T_314; // @[Arbiter.scala 21:28]
  wire [3:0] _T_316 = {_T_315,_T_133,_T_131}; // @[Cat.scala 29:58]
  wire [3:0] _GEN_24 = {{1'd0}, _T_316[3:1]}; // @[package.scala 208:43]
  wire [3:0] _T_318 = _T_316 | _GEN_24; // @[package.scala 208:43]
  wire [3:0] _T_321 = {_T_313, 2'h0}; // @[Arbiter.scala 22:66]
  wire [3:0] _GEN_25 = {{1'd0}, _T_318[3:1]}; // @[Arbiter.scala 22:58]
  wire [3:0] _T_322 = _GEN_25 | _T_321; // @[Arbiter.scala 22:58]
  wire [1:0] _T_325 = _T_322[3:2] & _T_322[1:0]; // @[Arbiter.scala 23:39]
  wire [1:0] _T_326 = ~_T_325; // @[Arbiter.scala 23:18]
  wire  _T_327 = _T_306 != 2'h0; // @[Arbiter.scala 24:27]
  wire  _T_328 = _T_304 & _T_327; // @[Arbiter.scala 24:18]
  wire [1:0] _T_329 = _T_326 & _T_306; // @[Arbiter.scala 25:29]
  wire [2:0] _T_330 = {_T_329, 1'h0}; // @[package.scala 199:48]
  wire [1:0] _T_332 = _T_329 | _T_330[1:0]; // @[package.scala 199:43]
  wire  _T_338 = _T_326[0] & _T_131; // @[Xbar.scala 250:63]
  wire  _T_339 = _T_326[1] & _T_133; // @[Xbar.scala 250:63]
  wire  _T_342 = _T_338 | _T_339; // @[Xbar.scala 255:50]
  wire  _T_344 = ~_T_338; // @[Xbar.scala 256:60]
  wire  _T_347 = ~_T_339; // @[Xbar.scala 256:60]
  wire  _T_348 = _T_344 | _T_347; // @[Xbar.scala 256:57]
  wire  _T_351 = _T_348 | reset; // @[Xbar.scala 256:11]
  wire  _T_352 = ~_T_351; // @[Xbar.scala 256:11]
  wire  _T_353 = ~_T_305; // @[Xbar.scala 258:13]
  wire  _T_355 = _T_353 | _T_342; // @[Xbar.scala 258:23]
  wire  _T_357 = _T_355 | reset; // @[Xbar.scala 258:12]
  wire  _T_358 = ~_T_357; // @[Xbar.scala 258:12]
  wire  _T_361_0 = _T_304 ? _T_338 : _T_360_0; // @[Xbar.scala 262:23]
  wire  _T_361_1 = _T_304 ? _T_339 : _T_360_1; // @[Xbar.scala 262:23]
  wire  _GEN_16 = _T_305 ? 1'h0 : _T_304; // @[Xbar.scala 266:21]
  wire  _GEN_17 = _T_62 | _GEN_16; // @[Xbar.scala 267:24]
  wire  _T_363_0 = _T_304 ? _T_326[0] : _T_360_0; // @[Xbar.scala 270:24]
  wire  _T_363_1 = _T_304 ? _T_326[1] : _T_360_1; // @[Xbar.scala 270:24]
  wire [2:0] _T_371 = {auto_out_0_b_bits_id,auto_out_0_b_bits_resp}; // @[Mux.scala 27:72]
  wire [2:0] _T_372 = _T_361_0 ? _T_371 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_373 = {auto_out_1_b_bits_id,auto_out_1_b_bits_resp}; // @[Mux.scala 27:72]
  wire [2:0] _T_374 = _T_361_1 ? _T_373 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_375 = _T_372 | _T_374; // @[Mux.scala 27:72]
  QueueCompatibility awIn_0 ( // @[Xbar.scala 55:47]
    .clock(awIn_0_clock),
    .reset(awIn_0_reset),
    .io_enq_ready(awIn_0_io_enq_ready),
    .io_enq_valid(awIn_0_io_enq_valid),
    .io_enq_bits(awIn_0_io_enq_bits),
    .io_deq_ready(awIn_0_io_deq_ready),
    .io_deq_valid(awIn_0_io_deq_valid),
    .io_deq_bits(awIn_0_io_deq_bits)
  );
  assign auto_in_aw_ready = _T_95 & _T_87; // @[LazyModule.scala 173:31]
  assign auto_in_w_ready = in_0_w_ready & awIn_0_io_deq_valid; // @[LazyModule.scala 173:31]
  assign auto_in_b_valid = _T_304 ? _T_305 : _T_368; // @[LazyModule.scala 173:31]
  assign auto_in_b_bits_resp = _T_375[1:0]; // @[LazyModule.scala 173:31]
  assign auto_in_ar_ready = in_0_ar_ready & _T_59; // @[LazyModule.scala 173:31]
  assign auto_in_r_valid = _T_222 ? _T_223 : _T_286; // @[LazyModule.scala 173:31]
  assign auto_in_r_bits_data = _T_297[34:3]; // @[LazyModule.scala 173:31]
  assign auto_in_r_bits_resp = _T_297[2:1]; // @[LazyModule.scala 173:31]
  assign auto_in_r_bits_last = _T_297[0]; // @[LazyModule.scala 173:31]
  assign auto_out_1_aw_valid = in_0_aw_valid & requestAWIO_0_1; // @[LazyModule.scala 173:49]
  assign auto_out_1_aw_bits_id = auto_in_aw_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_1_aw_bits_addr = auto_in_aw_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_1_aw_bits_size = auto_in_aw_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_1_w_valid = in_0_w_valid & requestWIO_0_1; // @[LazyModule.scala 173:49]
  assign auto_out_1_w_bits_data = auto_in_w_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_1_w_bits_strb = auto_in_w_bits_strb; // @[LazyModule.scala 173:49]
  assign auto_out_1_w_bits_last = auto_in_w_bits_last; // @[LazyModule.scala 173:49]
  assign auto_out_1_b_ready = auto_in_b_ready & _T_363_1; // @[LazyModule.scala 173:49]
  assign auto_out_1_ar_valid = in_0_ar_valid & requestARIO_0_1; // @[LazyModule.scala 173:49]
  assign auto_out_1_ar_bits_id = auto_in_ar_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_1_ar_bits_addr = auto_in_ar_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_1_ar_bits_size = auto_in_ar_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_1_r_ready = auto_in_r_ready & _T_281_1; // @[LazyModule.scala 173:49]
  assign auto_out_0_aw_valid = in_0_aw_valid & requestAWIO_0_0; // @[LazyModule.scala 173:49]
  assign auto_out_0_aw_bits_id = auto_in_aw_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_0_aw_bits_addr = auto_in_aw_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_0_aw_bits_size = auto_in_aw_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_0_w_valid = in_0_w_valid & requestWIO_0_0; // @[LazyModule.scala 173:49]
  assign auto_out_0_w_bits_data = auto_in_w_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_0_w_bits_strb = auto_in_w_bits_strb; // @[LazyModule.scala 173:49]
  assign auto_out_0_w_bits_last = auto_in_w_bits_last; // @[LazyModule.scala 173:49]
  assign auto_out_0_b_ready = auto_in_b_ready & _T_363_0; // @[LazyModule.scala 173:49]
  assign auto_out_0_ar_valid = in_0_ar_valid & requestARIO_0_0; // @[LazyModule.scala 173:49]
  assign auto_out_0_ar_bits_id = auto_in_ar_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_0_ar_bits_addr = auto_in_ar_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_0_ar_bits_size = auto_in_ar_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_0_r_ready = auto_in_r_ready & _T_281_0; // @[LazyModule.scala 173:49]
  assign awIn_0_clock = clock;
  assign awIn_0_reset = reset;
  assign awIn_0_io_enq_valid = auto_in_aw_valid & _T_97; // @[Xbar.scala 140:30]
  assign awIn_0_io_enq_bits = {requestAWIO_0_1,requestAWIO_0_0}; // @[Xbar.scala 64:57]
  assign awIn_0_io_deq_ready = _T_103 & in_0_w_ready; // @[Xbar.scala 147:30]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_36 = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_37 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_222 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_278_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_278_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_231 = _RAND_5[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_90 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_64 = _RAND_7[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_65 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_304 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_360_0 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_360_1 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_313 = _RAND_12[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      _T_36 <= 3'h0;
    end else begin
      _T_36 <= _T_41;
    end
    if (_T_31) begin
      _T_37 <= _T_27[1];
    end
    _T_222 <= reset | _GEN_14;
    if (reset) begin
      _T_278_0 <= 1'h0;
    end else if (_T_222) begin
      _T_278_0 <= _T_256;
    end
    if (reset) begin
      _T_278_1 <= 1'h0;
    end else if (_T_222) begin
      _T_278_1 <= _T_257;
    end
    if (reset) begin
      _T_231 <= 2'h3;
    end else if (_T_246) begin
      _T_231 <= _T_250;
    end
    if (reset) begin
      _T_90 <= 1'h0;
    end else if (_T_100) begin
      _T_90 <= 1'h0;
    end else begin
      _T_90 <= _GEN_2;
    end
    if (reset) begin
      _T_64 <= 3'h0;
    end else begin
      _T_64 <= _T_69;
    end
    if (_T_60) begin
      _T_65 <= _T_20[1];
    end
    _T_304 <= reset | _GEN_17;
    if (reset) begin
      _T_360_0 <= 1'h0;
    end else if (_T_304) begin
      _T_360_0 <= _T_338;
    end
    if (reset) begin
      _T_360_1 <= 1'h0;
    end else if (_T_304) begin
      _T_360_1 <= _T_339;
    end
    if (reset) begin
      _T_313 <= 2'h3;
    end else if (_T_328) begin
      _T_313 <= _T_332;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_47) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:107 assert (!resp_fire || count =/= UInt(0))\n"); // @[Xbar.scala 107:22]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_47) begin
          $fatal; // @[Xbar.scala 107:22]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_53) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:108 assert (!req_fire  || count =/= UInt(flight))\n"); // @[Xbar.scala 108:22]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_53) begin
          $fatal; // @[Xbar.scala 108:22]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_75) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:107 assert (!resp_fire || count =/= UInt(0))\n"); // @[Xbar.scala 107:22]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_75) begin
          $fatal; // @[Xbar.scala 107:22]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_81) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:108 assert (!req_fire  || count =/= UInt(flight))\n"); // @[Xbar.scala 108:22]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_81) begin
          $fatal; // @[Xbar.scala 108:22]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_149) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_149) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_170) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_170) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_193) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_193) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_214) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_214) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_270) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:256 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n"); // @[Xbar.scala 256:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_270) begin
          $fatal; // @[Xbar.scala 256:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_276) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_276) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_352) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:256 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n"); // @[Xbar.scala 256:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_352) begin
          $fatal; // @[Xbar.scala 256:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_358) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_358) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module Queue_25(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input         io_enq_bits_id,
  input  [29:0] io_enq_bits_addr,
  input  [2:0]  io_enq_bits_size,
  input         io_deq_ready,
  output        io_deq_valid,
  output        io_deq_bits_id,
  output [29:0] io_deq_bits_addr,
  output [2:0]  io_deq_bits_size
);
  reg  _T_id [0:1]; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_0;
  wire  _T_id__T_18_data; // @[Decoupled.scala 218:24]
  wire  _T_id__T_18_addr; // @[Decoupled.scala 218:24]
  wire  _T_id__T_10_data; // @[Decoupled.scala 218:24]
  wire  _T_id__T_10_addr; // @[Decoupled.scala 218:24]
  wire  _T_id__T_10_mask; // @[Decoupled.scala 218:24]
  wire  _T_id__T_10_en; // @[Decoupled.scala 218:24]
  reg [29:0] _T_addr [0:1]; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_1;
  wire [29:0] _T_addr__T_18_data; // @[Decoupled.scala 218:24]
  wire  _T_addr__T_18_addr; // @[Decoupled.scala 218:24]
  wire [29:0] _T_addr__T_10_data; // @[Decoupled.scala 218:24]
  wire  _T_addr__T_10_addr; // @[Decoupled.scala 218:24]
  wire  _T_addr__T_10_mask; // @[Decoupled.scala 218:24]
  wire  _T_addr__T_10_en; // @[Decoupled.scala 218:24]
  reg [2:0] _T_size [0:1]; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_2;
  wire [2:0] _T_size__T_18_data; // @[Decoupled.scala 218:24]
  wire  _T_size__T_18_addr; // @[Decoupled.scala 218:24]
  wire [2:0] _T_size__T_10_data; // @[Decoupled.scala 218:24]
  wire  _T_size__T_10_addr; // @[Decoupled.scala 218:24]
  wire  _T_size__T_10_mask; // @[Decoupled.scala 218:24]
  wire  _T_size__T_10_en; // @[Decoupled.scala 218:24]
  reg  value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_3;
  reg  value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_4;
  reg  _T_1; // @[Decoupled.scala 221:35]
  reg [31:0] _RAND_5;
  wire  _T_2 = value == value_1; // @[Decoupled.scala 223:41]
  wire  _T_3 = ~_T_1; // @[Decoupled.scala 224:36]
  wire  _T_4 = _T_2 & _T_3; // @[Decoupled.scala 224:33]
  wire  _T_5 = _T_2 & _T_1; // @[Decoupled.scala 225:32]
  wire  _T_6 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  _T_8 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire  _T_12 = value + 1'h1; // @[Counter.scala 39:22]
  wire  _T_14 = value_1 + 1'h1; // @[Counter.scala 39:22]
  wire  _T_15 = _T_6 != _T_8; // @[Decoupled.scala 236:16]
  assign _T_id__T_18_addr = value_1;
  assign _T_id__T_18_data = _T_id[_T_id__T_18_addr]; // @[Decoupled.scala 218:24]
  assign _T_id__T_10_data = io_enq_bits_id;
  assign _T_id__T_10_addr = value;
  assign _T_id__T_10_mask = 1'h1;
  assign _T_id__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_addr__T_18_addr = value_1;
  assign _T_addr__T_18_data = _T_addr[_T_addr__T_18_addr]; // @[Decoupled.scala 218:24]
  assign _T_addr__T_10_data = io_enq_bits_addr;
  assign _T_addr__T_10_addr = value;
  assign _T_addr__T_10_mask = 1'h1;
  assign _T_addr__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_size__T_18_addr = value_1;
  assign _T_size__T_18_data = _T_size[_T_size__T_18_addr]; // @[Decoupled.scala 218:24]
  assign _T_size__T_10_data = io_enq_bits_size;
  assign _T_size__T_10_addr = value;
  assign _T_size__T_10_mask = 1'h1;
  assign _T_size__T_10_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~_T_5; // @[Decoupled.scala 241:16]
  assign io_deq_valid = ~_T_4; // @[Decoupled.scala 240:16]
  assign io_deq_bits_id = _T_id__T_18_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_addr = _T_addr__T_18_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_size = _T_size__T_18_data; // @[Decoupled.scala 242:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_id[initvar] = _RAND_0[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_addr[initvar] = _RAND_1[29:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_size[initvar] = _RAND_2[2:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  value = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  value_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_1 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T_id__T_10_en & _T_id__T_10_mask) begin
      _T_id[_T_id__T_10_addr] <= _T_id__T_10_data; // @[Decoupled.scala 218:24]
    end
    if(_T_addr__T_10_en & _T_addr__T_10_mask) begin
      _T_addr[_T_addr__T_10_addr] <= _T_addr__T_10_data; // @[Decoupled.scala 218:24]
    end
    if(_T_size__T_10_en & _T_size__T_10_mask) begin
      _T_size[_T_size__T_10_addr] <= _T_size__T_10_data; // @[Decoupled.scala 218:24]
    end
    if (reset) begin
      value <= 1'h0;
    end else if (_T_6) begin
      value <= _T_12;
    end
    if (reset) begin
      value_1 <= 1'h0;
    end else if (_T_8) begin
      value_1 <= _T_14;
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else if (_T_15) begin
      _T_1 <= _T_6;
    end
  end
endmodule
module Queue_26(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [31:0] io_enq_bits_data,
  input  [3:0]  io_enq_bits_strb,
  input         io_enq_bits_last,
  input         io_deq_ready,
  output        io_deq_valid,
  output [31:0] io_deq_bits_data,
  output [3:0]  io_deq_bits_strb,
  output        io_deq_bits_last
);
  reg [31:0] _T_data [0:1]; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_0;
  wire [31:0] _T_data__T_18_data; // @[Decoupled.scala 218:24]
  wire  _T_data__T_18_addr; // @[Decoupled.scala 218:24]
  wire [31:0] _T_data__T_10_data; // @[Decoupled.scala 218:24]
  wire  _T_data__T_10_addr; // @[Decoupled.scala 218:24]
  wire  _T_data__T_10_mask; // @[Decoupled.scala 218:24]
  wire  _T_data__T_10_en; // @[Decoupled.scala 218:24]
  reg [3:0] _T_strb [0:1]; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_1;
  wire [3:0] _T_strb__T_18_data; // @[Decoupled.scala 218:24]
  wire  _T_strb__T_18_addr; // @[Decoupled.scala 218:24]
  wire [3:0] _T_strb__T_10_data; // @[Decoupled.scala 218:24]
  wire  _T_strb__T_10_addr; // @[Decoupled.scala 218:24]
  wire  _T_strb__T_10_mask; // @[Decoupled.scala 218:24]
  wire  _T_strb__T_10_en; // @[Decoupled.scala 218:24]
  reg  _T_last [0:1]; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_2;
  wire  _T_last__T_18_data; // @[Decoupled.scala 218:24]
  wire  _T_last__T_18_addr; // @[Decoupled.scala 218:24]
  wire  _T_last__T_10_data; // @[Decoupled.scala 218:24]
  wire  _T_last__T_10_addr; // @[Decoupled.scala 218:24]
  wire  _T_last__T_10_mask; // @[Decoupled.scala 218:24]
  wire  _T_last__T_10_en; // @[Decoupled.scala 218:24]
  reg  value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_3;
  reg  value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_4;
  reg  _T_1; // @[Decoupled.scala 221:35]
  reg [31:0] _RAND_5;
  wire  _T_2 = value == value_1; // @[Decoupled.scala 223:41]
  wire  _T_3 = ~_T_1; // @[Decoupled.scala 224:36]
  wire  _T_4 = _T_2 & _T_3; // @[Decoupled.scala 224:33]
  wire  _T_5 = _T_2 & _T_1; // @[Decoupled.scala 225:32]
  wire  _T_6 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  _T_8 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire  _T_12 = value + 1'h1; // @[Counter.scala 39:22]
  wire  _T_14 = value_1 + 1'h1; // @[Counter.scala 39:22]
  wire  _T_15 = _T_6 != _T_8; // @[Decoupled.scala 236:16]
  assign _T_data__T_18_addr = value_1;
  assign _T_data__T_18_data = _T_data[_T_data__T_18_addr]; // @[Decoupled.scala 218:24]
  assign _T_data__T_10_data = io_enq_bits_data;
  assign _T_data__T_10_addr = value;
  assign _T_data__T_10_mask = 1'h1;
  assign _T_data__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_strb__T_18_addr = value_1;
  assign _T_strb__T_18_data = _T_strb[_T_strb__T_18_addr]; // @[Decoupled.scala 218:24]
  assign _T_strb__T_10_data = io_enq_bits_strb;
  assign _T_strb__T_10_addr = value;
  assign _T_strb__T_10_mask = 1'h1;
  assign _T_strb__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_last__T_18_addr = value_1;
  assign _T_last__T_18_data = _T_last[_T_last__T_18_addr]; // @[Decoupled.scala 218:24]
  assign _T_last__T_10_data = io_enq_bits_last;
  assign _T_last__T_10_addr = value;
  assign _T_last__T_10_mask = 1'h1;
  assign _T_last__T_10_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~_T_5; // @[Decoupled.scala 241:16]
  assign io_deq_valid = ~_T_4; // @[Decoupled.scala 240:16]
  assign io_deq_bits_data = _T_data__T_18_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_strb = _T_strb__T_18_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_last = _T_last__T_18_data; // @[Decoupled.scala 242:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_data[initvar] = _RAND_0[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_strb[initvar] = _RAND_1[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_last[initvar] = _RAND_2[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  value = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  value_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_1 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T_data__T_10_en & _T_data__T_10_mask) begin
      _T_data[_T_data__T_10_addr] <= _T_data__T_10_data; // @[Decoupled.scala 218:24]
    end
    if(_T_strb__T_10_en & _T_strb__T_10_mask) begin
      _T_strb[_T_strb__T_10_addr] <= _T_strb__T_10_data; // @[Decoupled.scala 218:24]
    end
    if(_T_last__T_10_en & _T_last__T_10_mask) begin
      _T_last[_T_last__T_10_addr] <= _T_last__T_10_data; // @[Decoupled.scala 218:24]
    end
    if (reset) begin
      value <= 1'h0;
    end else if (_T_6) begin
      value <= _T_12;
    end
    if (reset) begin
      value_1 <= 1'h0;
    end else if (_T_8) begin
      value_1 <= _T_14;
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else if (_T_15) begin
      _T_1 <= _T_6;
    end
  end
endmodule
module Queue_27(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input        io_enq_bits_id,
  input  [1:0] io_enq_bits_resp,
  input        io_deq_ready,
  output       io_deq_valid,
  output       io_deq_bits_id,
  output [1:0] io_deq_bits_resp
);
  reg  _T_id [0:1]; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_0;
  wire  _T_id__T_18_data; // @[Decoupled.scala 218:24]
  wire  _T_id__T_18_addr; // @[Decoupled.scala 218:24]
  wire  _T_id__T_10_data; // @[Decoupled.scala 218:24]
  wire  _T_id__T_10_addr; // @[Decoupled.scala 218:24]
  wire  _T_id__T_10_mask; // @[Decoupled.scala 218:24]
  wire  _T_id__T_10_en; // @[Decoupled.scala 218:24]
  reg [1:0] _T_resp [0:1]; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_1;
  wire [1:0] _T_resp__T_18_data; // @[Decoupled.scala 218:24]
  wire  _T_resp__T_18_addr; // @[Decoupled.scala 218:24]
  wire [1:0] _T_resp__T_10_data; // @[Decoupled.scala 218:24]
  wire  _T_resp__T_10_addr; // @[Decoupled.scala 218:24]
  wire  _T_resp__T_10_mask; // @[Decoupled.scala 218:24]
  wire  _T_resp__T_10_en; // @[Decoupled.scala 218:24]
  reg  value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_2;
  reg  value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_3;
  reg  _T_1; // @[Decoupled.scala 221:35]
  reg [31:0] _RAND_4;
  wire  _T_2 = value == value_1; // @[Decoupled.scala 223:41]
  wire  _T_3 = ~_T_1; // @[Decoupled.scala 224:36]
  wire  _T_4 = _T_2 & _T_3; // @[Decoupled.scala 224:33]
  wire  _T_5 = _T_2 & _T_1; // @[Decoupled.scala 225:32]
  wire  _T_6 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  _T_8 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire  _T_12 = value + 1'h1; // @[Counter.scala 39:22]
  wire  _T_14 = value_1 + 1'h1; // @[Counter.scala 39:22]
  wire  _T_15 = _T_6 != _T_8; // @[Decoupled.scala 236:16]
  assign _T_id__T_18_addr = value_1;
  assign _T_id__T_18_data = _T_id[_T_id__T_18_addr]; // @[Decoupled.scala 218:24]
  assign _T_id__T_10_data = io_enq_bits_id;
  assign _T_id__T_10_addr = value;
  assign _T_id__T_10_mask = 1'h1;
  assign _T_id__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_resp__T_18_addr = value_1;
  assign _T_resp__T_18_data = _T_resp[_T_resp__T_18_addr]; // @[Decoupled.scala 218:24]
  assign _T_resp__T_10_data = io_enq_bits_resp;
  assign _T_resp__T_10_addr = value;
  assign _T_resp__T_10_mask = 1'h1;
  assign _T_resp__T_10_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~_T_5; // @[Decoupled.scala 241:16]
  assign io_deq_valid = ~_T_4; // @[Decoupled.scala 240:16]
  assign io_deq_bits_id = _T_id__T_18_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_resp = _T_resp__T_18_data; // @[Decoupled.scala 242:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_id[initvar] = _RAND_0[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_resp[initvar] = _RAND_1[1:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  value = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  value_1 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T_id__T_10_en & _T_id__T_10_mask) begin
      _T_id[_T_id__T_10_addr] <= _T_id__T_10_data; // @[Decoupled.scala 218:24]
    end
    if(_T_resp__T_10_en & _T_resp__T_10_mask) begin
      _T_resp[_T_resp__T_10_addr] <= _T_resp__T_10_data; // @[Decoupled.scala 218:24]
    end
    if (reset) begin
      value <= 1'h0;
    end else if (_T_6) begin
      value <= _T_12;
    end
    if (reset) begin
      value_1 <= 1'h0;
    end else if (_T_8) begin
      value_1 <= _T_14;
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else if (_T_15) begin
      _T_1 <= _T_6;
    end
  end
endmodule
module Queue_29(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input         io_enq_bits_id,
  input  [31:0] io_enq_bits_data,
  input  [1:0]  io_enq_bits_resp,
  input         io_enq_bits_last,
  input         io_deq_ready,
  output        io_deq_valid,
  output        io_deq_bits_id,
  output [31:0] io_deq_bits_data,
  output [1:0]  io_deq_bits_resp,
  output        io_deq_bits_last
);
  reg  _T_id [0:1]; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_0;
  wire  _T_id__T_18_data; // @[Decoupled.scala 218:24]
  wire  _T_id__T_18_addr; // @[Decoupled.scala 218:24]
  wire  _T_id__T_10_data; // @[Decoupled.scala 218:24]
  wire  _T_id__T_10_addr; // @[Decoupled.scala 218:24]
  wire  _T_id__T_10_mask; // @[Decoupled.scala 218:24]
  wire  _T_id__T_10_en; // @[Decoupled.scala 218:24]
  reg [31:0] _T_data [0:1]; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_1;
  wire [31:0] _T_data__T_18_data; // @[Decoupled.scala 218:24]
  wire  _T_data__T_18_addr; // @[Decoupled.scala 218:24]
  wire [31:0] _T_data__T_10_data; // @[Decoupled.scala 218:24]
  wire  _T_data__T_10_addr; // @[Decoupled.scala 218:24]
  wire  _T_data__T_10_mask; // @[Decoupled.scala 218:24]
  wire  _T_data__T_10_en; // @[Decoupled.scala 218:24]
  reg [1:0] _T_resp [0:1]; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_2;
  wire [1:0] _T_resp__T_18_data; // @[Decoupled.scala 218:24]
  wire  _T_resp__T_18_addr; // @[Decoupled.scala 218:24]
  wire [1:0] _T_resp__T_10_data; // @[Decoupled.scala 218:24]
  wire  _T_resp__T_10_addr; // @[Decoupled.scala 218:24]
  wire  _T_resp__T_10_mask; // @[Decoupled.scala 218:24]
  wire  _T_resp__T_10_en; // @[Decoupled.scala 218:24]
  reg  _T_last [0:1]; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_3;
  wire  _T_last__T_18_data; // @[Decoupled.scala 218:24]
  wire  _T_last__T_18_addr; // @[Decoupled.scala 218:24]
  wire  _T_last__T_10_data; // @[Decoupled.scala 218:24]
  wire  _T_last__T_10_addr; // @[Decoupled.scala 218:24]
  wire  _T_last__T_10_mask; // @[Decoupled.scala 218:24]
  wire  _T_last__T_10_en; // @[Decoupled.scala 218:24]
  reg  value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_4;
  reg  value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  reg  _T_1; // @[Decoupled.scala 221:35]
  reg [31:0] _RAND_6;
  wire  _T_2 = value == value_1; // @[Decoupled.scala 223:41]
  wire  _T_3 = ~_T_1; // @[Decoupled.scala 224:36]
  wire  _T_4 = _T_2 & _T_3; // @[Decoupled.scala 224:33]
  wire  _T_5 = _T_2 & _T_1; // @[Decoupled.scala 225:32]
  wire  _T_6 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  _T_8 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire  _T_12 = value + 1'h1; // @[Counter.scala 39:22]
  wire  _T_14 = value_1 + 1'h1; // @[Counter.scala 39:22]
  wire  _T_15 = _T_6 != _T_8; // @[Decoupled.scala 236:16]
  assign _T_id__T_18_addr = value_1;
  assign _T_id__T_18_data = _T_id[_T_id__T_18_addr]; // @[Decoupled.scala 218:24]
  assign _T_id__T_10_data = io_enq_bits_id;
  assign _T_id__T_10_addr = value;
  assign _T_id__T_10_mask = 1'h1;
  assign _T_id__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_data__T_18_addr = value_1;
  assign _T_data__T_18_data = _T_data[_T_data__T_18_addr]; // @[Decoupled.scala 218:24]
  assign _T_data__T_10_data = io_enq_bits_data;
  assign _T_data__T_10_addr = value;
  assign _T_data__T_10_mask = 1'h1;
  assign _T_data__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_resp__T_18_addr = value_1;
  assign _T_resp__T_18_data = _T_resp[_T_resp__T_18_addr]; // @[Decoupled.scala 218:24]
  assign _T_resp__T_10_data = io_enq_bits_resp;
  assign _T_resp__T_10_addr = value;
  assign _T_resp__T_10_mask = 1'h1;
  assign _T_resp__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_last__T_18_addr = value_1;
  assign _T_last__T_18_data = _T_last[_T_last__T_18_addr]; // @[Decoupled.scala 218:24]
  assign _T_last__T_10_data = io_enq_bits_last;
  assign _T_last__T_10_addr = value;
  assign _T_last__T_10_mask = 1'h1;
  assign _T_last__T_10_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~_T_5; // @[Decoupled.scala 241:16]
  assign io_deq_valid = ~_T_4; // @[Decoupled.scala 240:16]
  assign io_deq_bits_id = _T_id__T_18_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_data = _T_data__T_18_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_resp = _T_resp__T_18_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_last = _T_last__T_18_data; // @[Decoupled.scala 242:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_id[initvar] = _RAND_0[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_data[initvar] = _RAND_1[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_resp[initvar] = _RAND_2[1:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_last[initvar] = _RAND_3[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  value = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value_1 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_1 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T_id__T_10_en & _T_id__T_10_mask) begin
      _T_id[_T_id__T_10_addr] <= _T_id__T_10_data; // @[Decoupled.scala 218:24]
    end
    if(_T_data__T_10_en & _T_data__T_10_mask) begin
      _T_data[_T_data__T_10_addr] <= _T_data__T_10_data; // @[Decoupled.scala 218:24]
    end
    if(_T_resp__T_10_en & _T_resp__T_10_mask) begin
      _T_resp[_T_resp__T_10_addr] <= _T_resp__T_10_data; // @[Decoupled.scala 218:24]
    end
    if(_T_last__T_10_en & _T_last__T_10_mask) begin
      _T_last[_T_last__T_10_addr] <= _T_last__T_10_data; // @[Decoupled.scala 218:24]
    end
    if (reset) begin
      value <= 1'h0;
    end else if (_T_6) begin
      value <= _T_12;
    end
    if (reset) begin
      value_1 <= 1'h0;
    end else if (_T_8) begin
      value_1 <= _T_14;
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else if (_T_15) begin
      _T_1 <= _T_6;
    end
  end
endmodule
module AXI4Buffer(
  input         clock,
  input         reset,
  output        auto_in_aw_ready,
  input         auto_in_aw_valid,
  input         auto_in_aw_bits_id,
  input  [29:0] auto_in_aw_bits_addr,
  input  [2:0]  auto_in_aw_bits_size,
  output        auto_in_w_ready,
  input         auto_in_w_valid,
  input  [31:0] auto_in_w_bits_data,
  input  [3:0]  auto_in_w_bits_strb,
  input         auto_in_w_bits_last,
  input         auto_in_b_ready,
  output        auto_in_b_valid,
  output        auto_in_b_bits_id,
  output [1:0]  auto_in_b_bits_resp,
  output        auto_in_ar_ready,
  input         auto_in_ar_valid,
  input         auto_in_ar_bits_id,
  input  [29:0] auto_in_ar_bits_addr,
  input  [2:0]  auto_in_ar_bits_size,
  input         auto_in_r_ready,
  output        auto_in_r_valid,
  output        auto_in_r_bits_id,
  output [31:0] auto_in_r_bits_data,
  output [1:0]  auto_in_r_bits_resp,
  output        auto_in_r_bits_last,
  input         auto_out_aw_ready,
  output        auto_out_aw_valid,
  output        auto_out_aw_bits_id,
  output [29:0] auto_out_aw_bits_addr,
  input         auto_out_w_ready,
  output        auto_out_w_valid,
  output [31:0] auto_out_w_bits_data,
  output [3:0]  auto_out_w_bits_strb,
  output        auto_out_w_bits_last,
  output        auto_out_b_ready,
  input         auto_out_b_valid,
  input         auto_out_b_bits_id,
  input  [1:0]  auto_out_b_bits_resp,
  input         auto_out_ar_ready,
  output        auto_out_ar_valid,
  output        auto_out_ar_bits_id,
  output [29:0] auto_out_ar_bits_addr,
  output [2:0]  auto_out_ar_bits_size,
  output        auto_out_r_ready,
  input         auto_out_r_valid,
  input         auto_out_r_bits_id,
  input  [31:0] auto_out_r_bits_data,
  input  [1:0]  auto_out_r_bits_resp,
  input         auto_out_r_bits_last
);
  wire  Queue_clock; // @[Decoupled.scala 296:21]
  wire  Queue_reset; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_bits_id; // @[Decoupled.scala 296:21]
  wire [29:0] Queue_io_enq_bits_addr; // @[Decoupled.scala 296:21]
  wire [2:0] Queue_io_enq_bits_size; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_bits_id; // @[Decoupled.scala 296:21]
  wire [29:0] Queue_io_deq_bits_addr; // @[Decoupled.scala 296:21]
  wire [2:0] Queue_io_deq_bits_size; // @[Decoupled.scala 296:21]
  wire  Queue_1_clock; // @[Decoupled.scala 296:21]
  wire  Queue_1_reset; // @[Decoupled.scala 296:21]
  wire  Queue_1_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  Queue_1_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [31:0] Queue_1_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire [3:0] Queue_1_io_enq_bits_strb; // @[Decoupled.scala 296:21]
  wire  Queue_1_io_enq_bits_last; // @[Decoupled.scala 296:21]
  wire  Queue_1_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  Queue_1_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [31:0] Queue_1_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire [3:0] Queue_1_io_deq_bits_strb; // @[Decoupled.scala 296:21]
  wire  Queue_1_io_deq_bits_last; // @[Decoupled.scala 296:21]
  wire  Queue_2_clock; // @[Decoupled.scala 296:21]
  wire  Queue_2_reset; // @[Decoupled.scala 296:21]
  wire  Queue_2_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  Queue_2_io_enq_valid; // @[Decoupled.scala 296:21]
  wire  Queue_2_io_enq_bits_id; // @[Decoupled.scala 296:21]
  wire [1:0] Queue_2_io_enq_bits_resp; // @[Decoupled.scala 296:21]
  wire  Queue_2_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  Queue_2_io_deq_valid; // @[Decoupled.scala 296:21]
  wire  Queue_2_io_deq_bits_id; // @[Decoupled.scala 296:21]
  wire [1:0] Queue_2_io_deq_bits_resp; // @[Decoupled.scala 296:21]
  wire  Queue_3_clock; // @[Decoupled.scala 296:21]
  wire  Queue_3_reset; // @[Decoupled.scala 296:21]
  wire  Queue_3_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  Queue_3_io_enq_valid; // @[Decoupled.scala 296:21]
  wire  Queue_3_io_enq_bits_id; // @[Decoupled.scala 296:21]
  wire [29:0] Queue_3_io_enq_bits_addr; // @[Decoupled.scala 296:21]
  wire [2:0] Queue_3_io_enq_bits_size; // @[Decoupled.scala 296:21]
  wire  Queue_3_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  Queue_3_io_deq_valid; // @[Decoupled.scala 296:21]
  wire  Queue_3_io_deq_bits_id; // @[Decoupled.scala 296:21]
  wire [29:0] Queue_3_io_deq_bits_addr; // @[Decoupled.scala 296:21]
  wire [2:0] Queue_3_io_deq_bits_size; // @[Decoupled.scala 296:21]
  wire  Queue_4_clock; // @[Decoupled.scala 296:21]
  wire  Queue_4_reset; // @[Decoupled.scala 296:21]
  wire  Queue_4_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  Queue_4_io_enq_valid; // @[Decoupled.scala 296:21]
  wire  Queue_4_io_enq_bits_id; // @[Decoupled.scala 296:21]
  wire [31:0] Queue_4_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] Queue_4_io_enq_bits_resp; // @[Decoupled.scala 296:21]
  wire  Queue_4_io_enq_bits_last; // @[Decoupled.scala 296:21]
  wire  Queue_4_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  Queue_4_io_deq_valid; // @[Decoupled.scala 296:21]
  wire  Queue_4_io_deq_bits_id; // @[Decoupled.scala 296:21]
  wire [31:0] Queue_4_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] Queue_4_io_deq_bits_resp; // @[Decoupled.scala 296:21]
  wire  Queue_4_io_deq_bits_last; // @[Decoupled.scala 296:21]
  Queue_25 Queue ( // @[Decoupled.scala 296:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_id(Queue_io_enq_bits_id),
    .io_enq_bits_addr(Queue_io_enq_bits_addr),
    .io_enq_bits_size(Queue_io_enq_bits_size),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_id(Queue_io_deq_bits_id),
    .io_deq_bits_addr(Queue_io_deq_bits_addr),
    .io_deq_bits_size(Queue_io_deq_bits_size)
  );
  Queue_26 Queue_1 ( // @[Decoupled.scala 296:21]
    .clock(Queue_1_clock),
    .reset(Queue_1_reset),
    .io_enq_ready(Queue_1_io_enq_ready),
    .io_enq_valid(Queue_1_io_enq_valid),
    .io_enq_bits_data(Queue_1_io_enq_bits_data),
    .io_enq_bits_strb(Queue_1_io_enq_bits_strb),
    .io_enq_bits_last(Queue_1_io_enq_bits_last),
    .io_deq_ready(Queue_1_io_deq_ready),
    .io_deq_valid(Queue_1_io_deq_valid),
    .io_deq_bits_data(Queue_1_io_deq_bits_data),
    .io_deq_bits_strb(Queue_1_io_deq_bits_strb),
    .io_deq_bits_last(Queue_1_io_deq_bits_last)
  );
  Queue_27 Queue_2 ( // @[Decoupled.scala 296:21]
    .clock(Queue_2_clock),
    .reset(Queue_2_reset),
    .io_enq_ready(Queue_2_io_enq_ready),
    .io_enq_valid(Queue_2_io_enq_valid),
    .io_enq_bits_id(Queue_2_io_enq_bits_id),
    .io_enq_bits_resp(Queue_2_io_enq_bits_resp),
    .io_deq_ready(Queue_2_io_deq_ready),
    .io_deq_valid(Queue_2_io_deq_valid),
    .io_deq_bits_id(Queue_2_io_deq_bits_id),
    .io_deq_bits_resp(Queue_2_io_deq_bits_resp)
  );
  Queue_25 Queue_3 ( // @[Decoupled.scala 296:21]
    .clock(Queue_3_clock),
    .reset(Queue_3_reset),
    .io_enq_ready(Queue_3_io_enq_ready),
    .io_enq_valid(Queue_3_io_enq_valid),
    .io_enq_bits_id(Queue_3_io_enq_bits_id),
    .io_enq_bits_addr(Queue_3_io_enq_bits_addr),
    .io_enq_bits_size(Queue_3_io_enq_bits_size),
    .io_deq_ready(Queue_3_io_deq_ready),
    .io_deq_valid(Queue_3_io_deq_valid),
    .io_deq_bits_id(Queue_3_io_deq_bits_id),
    .io_deq_bits_addr(Queue_3_io_deq_bits_addr),
    .io_deq_bits_size(Queue_3_io_deq_bits_size)
  );
  Queue_29 Queue_4 ( // @[Decoupled.scala 296:21]
    .clock(Queue_4_clock),
    .reset(Queue_4_reset),
    .io_enq_ready(Queue_4_io_enq_ready),
    .io_enq_valid(Queue_4_io_enq_valid),
    .io_enq_bits_id(Queue_4_io_enq_bits_id),
    .io_enq_bits_data(Queue_4_io_enq_bits_data),
    .io_enq_bits_resp(Queue_4_io_enq_bits_resp),
    .io_enq_bits_last(Queue_4_io_enq_bits_last),
    .io_deq_ready(Queue_4_io_deq_ready),
    .io_deq_valid(Queue_4_io_deq_valid),
    .io_deq_bits_id(Queue_4_io_deq_bits_id),
    .io_deq_bits_data(Queue_4_io_deq_bits_data),
    .io_deq_bits_resp(Queue_4_io_deq_bits_resp),
    .io_deq_bits_last(Queue_4_io_deq_bits_last)
  );
  assign auto_in_aw_ready = Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_in_w_ready = Queue_1_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_in_b_valid = Queue_2_io_deq_valid; // @[LazyModule.scala 173:31]
  assign auto_in_b_bits_id = Queue_2_io_deq_bits_id; // @[LazyModule.scala 173:31]
  assign auto_in_b_bits_resp = Queue_2_io_deq_bits_resp; // @[LazyModule.scala 173:31]
  assign auto_in_ar_ready = Queue_3_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_in_r_valid = Queue_4_io_deq_valid; // @[LazyModule.scala 173:31]
  assign auto_in_r_bits_id = Queue_4_io_deq_bits_id; // @[LazyModule.scala 173:31]
  assign auto_in_r_bits_data = Queue_4_io_deq_bits_data; // @[LazyModule.scala 173:31]
  assign auto_in_r_bits_resp = Queue_4_io_deq_bits_resp; // @[LazyModule.scala 173:31]
  assign auto_in_r_bits_last = Queue_4_io_deq_bits_last; // @[LazyModule.scala 173:31]
  assign auto_out_aw_valid = Queue_io_deq_valid; // @[LazyModule.scala 173:49]
  assign auto_out_aw_bits_id = Queue_io_deq_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_aw_bits_addr = Queue_io_deq_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_w_valid = Queue_1_io_deq_valid; // @[LazyModule.scala 173:49]
  assign auto_out_w_bits_data = Queue_1_io_deq_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_w_bits_strb = Queue_1_io_deq_bits_strb; // @[LazyModule.scala 173:49]
  assign auto_out_w_bits_last = Queue_1_io_deq_bits_last; // @[LazyModule.scala 173:49]
  assign auto_out_b_ready = Queue_2_io_enq_ready; // @[LazyModule.scala 173:49]
  assign auto_out_ar_valid = Queue_3_io_deq_valid; // @[LazyModule.scala 173:49]
  assign auto_out_ar_bits_id = Queue_3_io_deq_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_ar_bits_addr = Queue_3_io_deq_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_ar_bits_size = Queue_3_io_deq_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_r_ready = Queue_4_io_enq_ready; // @[LazyModule.scala 173:49]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_in_aw_valid; // @[Decoupled.scala 297:22]
  assign Queue_io_enq_bits_id = auto_in_aw_bits_id; // @[Decoupled.scala 298:21]
  assign Queue_io_enq_bits_addr = auto_in_aw_bits_addr; // @[Decoupled.scala 298:21]
  assign Queue_io_enq_bits_size = auto_in_aw_bits_size; // @[Decoupled.scala 298:21]
  assign Queue_io_deq_ready = auto_out_aw_ready; // @[Decoupled.scala 320:15]
  assign Queue_1_clock = clock;
  assign Queue_1_reset = reset;
  assign Queue_1_io_enq_valid = auto_in_w_valid; // @[Decoupled.scala 297:22]
  assign Queue_1_io_enq_bits_data = auto_in_w_bits_data; // @[Decoupled.scala 298:21]
  assign Queue_1_io_enq_bits_strb = auto_in_w_bits_strb; // @[Decoupled.scala 298:21]
  assign Queue_1_io_enq_bits_last = auto_in_w_bits_last; // @[Decoupled.scala 298:21]
  assign Queue_1_io_deq_ready = auto_out_w_ready; // @[Decoupled.scala 320:15]
  assign Queue_2_clock = clock;
  assign Queue_2_reset = reset;
  assign Queue_2_io_enq_valid = auto_out_b_valid; // @[Decoupled.scala 297:22]
  assign Queue_2_io_enq_bits_id = auto_out_b_bits_id; // @[Decoupled.scala 298:21]
  assign Queue_2_io_enq_bits_resp = auto_out_b_bits_resp; // @[Decoupled.scala 298:21]
  assign Queue_2_io_deq_ready = auto_in_b_ready; // @[Decoupled.scala 320:15]
  assign Queue_3_clock = clock;
  assign Queue_3_reset = reset;
  assign Queue_3_io_enq_valid = auto_in_ar_valid; // @[Decoupled.scala 297:22]
  assign Queue_3_io_enq_bits_id = auto_in_ar_bits_id; // @[Decoupled.scala 298:21]
  assign Queue_3_io_enq_bits_addr = auto_in_ar_bits_addr; // @[Decoupled.scala 298:21]
  assign Queue_3_io_enq_bits_size = auto_in_ar_bits_size; // @[Decoupled.scala 298:21]
  assign Queue_3_io_deq_ready = auto_out_ar_ready; // @[Decoupled.scala 320:15]
  assign Queue_4_clock = clock;
  assign Queue_4_reset = reset;
  assign Queue_4_io_enq_valid = auto_out_r_valid; // @[Decoupled.scala 297:22]
  assign Queue_4_io_enq_bits_id = auto_out_r_bits_id; // @[Decoupled.scala 298:21]
  assign Queue_4_io_enq_bits_data = auto_out_r_bits_data; // @[Decoupled.scala 298:21]
  assign Queue_4_io_enq_bits_resp = auto_out_r_bits_resp; // @[Decoupled.scala 298:21]
  assign Queue_4_io_enq_bits_last = auto_out_r_bits_last; // @[Decoupled.scala 298:21]
  assign Queue_4_io_deq_ready = auto_in_r_ready; // @[Decoupled.scala 320:15]
endmodule
module AccumulatorChain(
  input         clock,
  input         reset,
  output        auto_bus_in_aw_ready,
  input         auto_bus_in_aw_valid,
  input         auto_bus_in_aw_bits_id,
  input  [29:0] auto_bus_in_aw_bits_addr,
  input  [2:0]  auto_bus_in_aw_bits_size,
  output        auto_bus_in_w_ready,
  input         auto_bus_in_w_valid,
  input  [31:0] auto_bus_in_w_bits_data,
  input  [3:0]  auto_bus_in_w_bits_strb,
  input         auto_bus_in_w_bits_last,
  input         auto_bus_in_b_ready,
  output        auto_bus_in_b_valid,
  output [1:0]  auto_bus_in_b_bits_resp,
  output        auto_bus_in_ar_ready,
  input         auto_bus_in_ar_valid,
  input         auto_bus_in_ar_bits_id,
  input  [29:0] auto_bus_in_ar_bits_addr,
  input  [2:0]  auto_bus_in_ar_bits_size,
  input         auto_bus_in_r_ready,
  output        auto_bus_in_r_valid,
  output [31:0] auto_bus_in_r_bits_data,
  output [1:0]  auto_bus_in_r_bits_resp,
  output        auto_bus_in_r_bits_last,
  input         auto_dspQueue_stream_out_ready,
  output        auto_dspQueue_stream_out_valid,
  output [15:0] auto_dspQueue_stream_out_bits_data,
  output        auto_dspQueue_stream_out_bits_last,
  output        auto_accumulator_slave_in_ready,
  input         auto_accumulator_slave_in_valid,
  input  [31:0] auto_accumulator_slave_in_bits_data,
  input         auto_accumulator_slave_in_bits_last
);
  wire  accumulator_clock; // @[AccChain.scala 27:30]
  wire  accumulator_reset; // @[AccChain.scala 27:30]
  wire  accumulator_auto_mem_in_aw_ready; // @[AccChain.scala 27:30]
  wire  accumulator_auto_mem_in_aw_valid; // @[AccChain.scala 27:30]
  wire  accumulator_auto_mem_in_aw_bits_id; // @[AccChain.scala 27:30]
  wire [29:0] accumulator_auto_mem_in_aw_bits_addr; // @[AccChain.scala 27:30]
  wire  accumulator_auto_mem_in_w_ready; // @[AccChain.scala 27:30]
  wire  accumulator_auto_mem_in_w_valid; // @[AccChain.scala 27:30]
  wire [31:0] accumulator_auto_mem_in_w_bits_data; // @[AccChain.scala 27:30]
  wire [3:0] accumulator_auto_mem_in_w_bits_strb; // @[AccChain.scala 27:30]
  wire  accumulator_auto_mem_in_b_ready; // @[AccChain.scala 27:30]
  wire  accumulator_auto_mem_in_b_valid; // @[AccChain.scala 27:30]
  wire  accumulator_auto_mem_in_b_bits_id; // @[AccChain.scala 27:30]
  wire  accumulator_auto_mem_in_ar_ready; // @[AccChain.scala 27:30]
  wire  accumulator_auto_mem_in_ar_valid; // @[AccChain.scala 27:30]
  wire  accumulator_auto_mem_in_ar_bits_id; // @[AccChain.scala 27:30]
  wire [29:0] accumulator_auto_mem_in_ar_bits_addr; // @[AccChain.scala 27:30]
  wire [2:0] accumulator_auto_mem_in_ar_bits_size; // @[AccChain.scala 27:30]
  wire  accumulator_auto_mem_in_r_ready; // @[AccChain.scala 27:30]
  wire  accumulator_auto_mem_in_r_valid; // @[AccChain.scala 27:30]
  wire  accumulator_auto_mem_in_r_bits_id; // @[AccChain.scala 27:30]
  wire [31:0] accumulator_auto_mem_in_r_bits_data; // @[AccChain.scala 27:30]
  wire  accumulator_auto_master_out_ready; // @[AccChain.scala 27:30]
  wire  accumulator_auto_master_out_valid; // @[AccChain.scala 27:30]
  wire [15:0] accumulator_auto_master_out_bits_data; // @[AccChain.scala 27:30]
  wire  accumulator_auto_master_out_bits_last; // @[AccChain.scala 27:30]
  wire  accumulator_auto_slave_in_ready; // @[AccChain.scala 27:30]
  wire  accumulator_auto_slave_in_valid; // @[AccChain.scala 27:30]
  wire [31:0] accumulator_auto_slave_in_bits_data; // @[AccChain.scala 27:30]
  wire  accumulator_auto_slave_in_bits_last; // @[AccChain.scala 27:30]
  wire  dspQueue_clock; // @[AccChain.scala 29:27]
  wire  dspQueue_reset; // @[AccChain.scala 29:27]
  wire  dspQueue_auto_stream_in_ready; // @[AccChain.scala 29:27]
  wire  dspQueue_auto_stream_in_valid; // @[AccChain.scala 29:27]
  wire [15:0] dspQueue_auto_stream_in_bits_data; // @[AccChain.scala 29:27]
  wire  dspQueue_auto_stream_in_bits_last; // @[AccChain.scala 29:27]
  wire  dspQueue_auto_stream_out_ready; // @[AccChain.scala 29:27]
  wire  dspQueue_auto_stream_out_valid; // @[AccChain.scala 29:27]
  wire [15:0] dspQueue_auto_stream_out_bits_data; // @[AccChain.scala 29:27]
  wire  dspQueue_auto_stream_out_bits_last; // @[AccChain.scala 29:27]
  wire  dspQueue_auto_in_aw_ready; // @[AccChain.scala 29:27]
  wire  dspQueue_auto_in_aw_valid; // @[AccChain.scala 29:27]
  wire  dspQueue_auto_in_aw_bits_id; // @[AccChain.scala 29:27]
  wire [29:0] dspQueue_auto_in_aw_bits_addr; // @[AccChain.scala 29:27]
  wire  dspQueue_auto_in_w_ready; // @[AccChain.scala 29:27]
  wire  dspQueue_auto_in_w_valid; // @[AccChain.scala 29:27]
  wire [31:0] dspQueue_auto_in_w_bits_data; // @[AccChain.scala 29:27]
  wire [3:0] dspQueue_auto_in_w_bits_strb; // @[AccChain.scala 29:27]
  wire  dspQueue_auto_in_b_ready; // @[AccChain.scala 29:27]
  wire  dspQueue_auto_in_b_valid; // @[AccChain.scala 29:27]
  wire  dspQueue_auto_in_b_bits_id; // @[AccChain.scala 29:27]
  wire  dspQueue_auto_in_ar_ready; // @[AccChain.scala 29:27]
  wire  dspQueue_auto_in_ar_valid; // @[AccChain.scala 29:27]
  wire  dspQueue_auto_in_ar_bits_id; // @[AccChain.scala 29:27]
  wire [29:0] dspQueue_auto_in_ar_bits_addr; // @[AccChain.scala 29:27]
  wire [2:0] dspQueue_auto_in_ar_bits_size; // @[AccChain.scala 29:27]
  wire  dspQueue_auto_in_r_ready; // @[AccChain.scala 29:27]
  wire  dspQueue_auto_in_r_valid; // @[AccChain.scala 29:27]
  wire  dspQueue_auto_in_r_bits_id; // @[AccChain.scala 29:27]
  wire [31:0] dspQueue_auto_in_r_bits_data; // @[AccChain.scala 29:27]
  wire  bus_clock; // @[AccChain.scala 44:23]
  wire  bus_reset; // @[AccChain.scala 44:23]
  wire  bus_auto_in_aw_ready; // @[AccChain.scala 44:23]
  wire  bus_auto_in_aw_valid; // @[AccChain.scala 44:23]
  wire  bus_auto_in_aw_bits_id; // @[AccChain.scala 44:23]
  wire [29:0] bus_auto_in_aw_bits_addr; // @[AccChain.scala 44:23]
  wire [2:0] bus_auto_in_aw_bits_size; // @[AccChain.scala 44:23]
  wire  bus_auto_in_w_ready; // @[AccChain.scala 44:23]
  wire  bus_auto_in_w_valid; // @[AccChain.scala 44:23]
  wire [31:0] bus_auto_in_w_bits_data; // @[AccChain.scala 44:23]
  wire [3:0] bus_auto_in_w_bits_strb; // @[AccChain.scala 44:23]
  wire  bus_auto_in_w_bits_last; // @[AccChain.scala 44:23]
  wire  bus_auto_in_b_ready; // @[AccChain.scala 44:23]
  wire  bus_auto_in_b_valid; // @[AccChain.scala 44:23]
  wire [1:0] bus_auto_in_b_bits_resp; // @[AccChain.scala 44:23]
  wire  bus_auto_in_ar_ready; // @[AccChain.scala 44:23]
  wire  bus_auto_in_ar_valid; // @[AccChain.scala 44:23]
  wire  bus_auto_in_ar_bits_id; // @[AccChain.scala 44:23]
  wire [29:0] bus_auto_in_ar_bits_addr; // @[AccChain.scala 44:23]
  wire [2:0] bus_auto_in_ar_bits_size; // @[AccChain.scala 44:23]
  wire  bus_auto_in_r_ready; // @[AccChain.scala 44:23]
  wire  bus_auto_in_r_valid; // @[AccChain.scala 44:23]
  wire [31:0] bus_auto_in_r_bits_data; // @[AccChain.scala 44:23]
  wire [1:0] bus_auto_in_r_bits_resp; // @[AccChain.scala 44:23]
  wire  bus_auto_in_r_bits_last; // @[AccChain.scala 44:23]
  wire  bus_auto_out_1_aw_ready; // @[AccChain.scala 44:23]
  wire  bus_auto_out_1_aw_valid; // @[AccChain.scala 44:23]
  wire  bus_auto_out_1_aw_bits_id; // @[AccChain.scala 44:23]
  wire [29:0] bus_auto_out_1_aw_bits_addr; // @[AccChain.scala 44:23]
  wire [2:0] bus_auto_out_1_aw_bits_size; // @[AccChain.scala 44:23]
  wire  bus_auto_out_1_w_ready; // @[AccChain.scala 44:23]
  wire  bus_auto_out_1_w_valid; // @[AccChain.scala 44:23]
  wire [31:0] bus_auto_out_1_w_bits_data; // @[AccChain.scala 44:23]
  wire [3:0] bus_auto_out_1_w_bits_strb; // @[AccChain.scala 44:23]
  wire  bus_auto_out_1_w_bits_last; // @[AccChain.scala 44:23]
  wire  bus_auto_out_1_b_ready; // @[AccChain.scala 44:23]
  wire  bus_auto_out_1_b_valid; // @[AccChain.scala 44:23]
  wire  bus_auto_out_1_b_bits_id; // @[AccChain.scala 44:23]
  wire [1:0] bus_auto_out_1_b_bits_resp; // @[AccChain.scala 44:23]
  wire  bus_auto_out_1_ar_ready; // @[AccChain.scala 44:23]
  wire  bus_auto_out_1_ar_valid; // @[AccChain.scala 44:23]
  wire  bus_auto_out_1_ar_bits_id; // @[AccChain.scala 44:23]
  wire [29:0] bus_auto_out_1_ar_bits_addr; // @[AccChain.scala 44:23]
  wire [2:0] bus_auto_out_1_ar_bits_size; // @[AccChain.scala 44:23]
  wire  bus_auto_out_1_r_ready; // @[AccChain.scala 44:23]
  wire  bus_auto_out_1_r_valid; // @[AccChain.scala 44:23]
  wire  bus_auto_out_1_r_bits_id; // @[AccChain.scala 44:23]
  wire [31:0] bus_auto_out_1_r_bits_data; // @[AccChain.scala 44:23]
  wire [1:0] bus_auto_out_1_r_bits_resp; // @[AccChain.scala 44:23]
  wire  bus_auto_out_1_r_bits_last; // @[AccChain.scala 44:23]
  wire  bus_auto_out_0_aw_ready; // @[AccChain.scala 44:23]
  wire  bus_auto_out_0_aw_valid; // @[AccChain.scala 44:23]
  wire  bus_auto_out_0_aw_bits_id; // @[AccChain.scala 44:23]
  wire [29:0] bus_auto_out_0_aw_bits_addr; // @[AccChain.scala 44:23]
  wire [2:0] bus_auto_out_0_aw_bits_size; // @[AccChain.scala 44:23]
  wire  bus_auto_out_0_w_ready; // @[AccChain.scala 44:23]
  wire  bus_auto_out_0_w_valid; // @[AccChain.scala 44:23]
  wire [31:0] bus_auto_out_0_w_bits_data; // @[AccChain.scala 44:23]
  wire [3:0] bus_auto_out_0_w_bits_strb; // @[AccChain.scala 44:23]
  wire  bus_auto_out_0_w_bits_last; // @[AccChain.scala 44:23]
  wire  bus_auto_out_0_b_ready; // @[AccChain.scala 44:23]
  wire  bus_auto_out_0_b_valid; // @[AccChain.scala 44:23]
  wire  bus_auto_out_0_b_bits_id; // @[AccChain.scala 44:23]
  wire [1:0] bus_auto_out_0_b_bits_resp; // @[AccChain.scala 44:23]
  wire  bus_auto_out_0_ar_ready; // @[AccChain.scala 44:23]
  wire  bus_auto_out_0_ar_valid; // @[AccChain.scala 44:23]
  wire  bus_auto_out_0_ar_bits_id; // @[AccChain.scala 44:23]
  wire [29:0] bus_auto_out_0_ar_bits_addr; // @[AccChain.scala 44:23]
  wire [2:0] bus_auto_out_0_ar_bits_size; // @[AccChain.scala 44:23]
  wire  bus_auto_out_0_r_ready; // @[AccChain.scala 44:23]
  wire  bus_auto_out_0_r_valid; // @[AccChain.scala 44:23]
  wire  bus_auto_out_0_r_bits_id; // @[AccChain.scala 44:23]
  wire [31:0] bus_auto_out_0_r_bits_data; // @[AccChain.scala 44:23]
  wire [1:0] bus_auto_out_0_r_bits_resp; // @[AccChain.scala 44:23]
  wire  bus_auto_out_0_r_bits_last; // @[AccChain.scala 44:23]
  wire  axi4buf_clock; // @[Buffer.scala 58:29]
  wire  axi4buf_reset; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_in_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_in_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_in_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_auto_in_aw_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_auto_in_aw_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_in_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_in_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_auto_in_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_auto_in_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_in_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_in_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_in_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_in_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_auto_in_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_in_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_in_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_in_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_auto_in_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_auto_in_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_in_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_in_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_in_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_auto_in_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_auto_in_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_in_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_out_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_out_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_out_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_auto_out_aw_bits_addr; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_out_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_out_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_auto_out_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_auto_out_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_out_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_out_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_out_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_out_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_auto_out_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_out_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_out_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_out_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_auto_out_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_auto_out_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_out_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_out_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_out_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_auto_out_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_auto_out_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_out_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_1_clock; // @[Buffer.scala 58:29]
  wire  axi4buf_1_reset; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_in_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_in_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_in_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_1_auto_in_aw_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_1_auto_in_aw_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_in_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_in_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_1_auto_in_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_1_auto_in_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_in_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_in_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_in_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_in_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_1_auto_in_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_in_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_in_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_in_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_1_auto_in_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_1_auto_in_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_in_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_in_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_in_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_1_auto_in_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_1_auto_in_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_in_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_out_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_out_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_out_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_1_auto_out_aw_bits_addr; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_out_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_out_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_1_auto_out_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_1_auto_out_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_out_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_out_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_out_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_out_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_1_auto_out_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_out_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_out_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_out_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_1_auto_out_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_1_auto_out_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_out_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_out_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_out_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_1_auto_out_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_1_auto_out_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_out_r_bits_last; // @[Buffer.scala 58:29]
  AXI4AccumulatorBlock accumulator ( // @[AccChain.scala 27:30]
    .clock(accumulator_clock),
    .reset(accumulator_reset),
    .auto_mem_in_aw_ready(accumulator_auto_mem_in_aw_ready),
    .auto_mem_in_aw_valid(accumulator_auto_mem_in_aw_valid),
    .auto_mem_in_aw_bits_id(accumulator_auto_mem_in_aw_bits_id),
    .auto_mem_in_aw_bits_addr(accumulator_auto_mem_in_aw_bits_addr),
    .auto_mem_in_w_ready(accumulator_auto_mem_in_w_ready),
    .auto_mem_in_w_valid(accumulator_auto_mem_in_w_valid),
    .auto_mem_in_w_bits_data(accumulator_auto_mem_in_w_bits_data),
    .auto_mem_in_w_bits_strb(accumulator_auto_mem_in_w_bits_strb),
    .auto_mem_in_b_ready(accumulator_auto_mem_in_b_ready),
    .auto_mem_in_b_valid(accumulator_auto_mem_in_b_valid),
    .auto_mem_in_b_bits_id(accumulator_auto_mem_in_b_bits_id),
    .auto_mem_in_ar_ready(accumulator_auto_mem_in_ar_ready),
    .auto_mem_in_ar_valid(accumulator_auto_mem_in_ar_valid),
    .auto_mem_in_ar_bits_id(accumulator_auto_mem_in_ar_bits_id),
    .auto_mem_in_ar_bits_addr(accumulator_auto_mem_in_ar_bits_addr),
    .auto_mem_in_ar_bits_size(accumulator_auto_mem_in_ar_bits_size),
    .auto_mem_in_r_ready(accumulator_auto_mem_in_r_ready),
    .auto_mem_in_r_valid(accumulator_auto_mem_in_r_valid),
    .auto_mem_in_r_bits_id(accumulator_auto_mem_in_r_bits_id),
    .auto_mem_in_r_bits_data(accumulator_auto_mem_in_r_bits_data),
    .auto_master_out_ready(accumulator_auto_master_out_ready),
    .auto_master_out_valid(accumulator_auto_master_out_valid),
    .auto_master_out_bits_data(accumulator_auto_master_out_bits_data),
    .auto_master_out_bits_last(accumulator_auto_master_out_bits_last),
    .auto_slave_in_ready(accumulator_auto_slave_in_ready),
    .auto_slave_in_valid(accumulator_auto_slave_in_valid),
    .auto_slave_in_bits_data(accumulator_auto_slave_in_bits_data),
    .auto_slave_in_bits_last(accumulator_auto_slave_in_bits_last)
  );
  AXI4DspQueueBlock dspQueue ( // @[AccChain.scala 29:27]
    .clock(dspQueue_clock),
    .reset(dspQueue_reset),
    .auto_stream_in_ready(dspQueue_auto_stream_in_ready),
    .auto_stream_in_valid(dspQueue_auto_stream_in_valid),
    .auto_stream_in_bits_data(dspQueue_auto_stream_in_bits_data),
    .auto_stream_in_bits_last(dspQueue_auto_stream_in_bits_last),
    .auto_stream_out_ready(dspQueue_auto_stream_out_ready),
    .auto_stream_out_valid(dspQueue_auto_stream_out_valid),
    .auto_stream_out_bits_data(dspQueue_auto_stream_out_bits_data),
    .auto_stream_out_bits_last(dspQueue_auto_stream_out_bits_last),
    .auto_in_aw_ready(dspQueue_auto_in_aw_ready),
    .auto_in_aw_valid(dspQueue_auto_in_aw_valid),
    .auto_in_aw_bits_id(dspQueue_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(dspQueue_auto_in_aw_bits_addr),
    .auto_in_w_ready(dspQueue_auto_in_w_ready),
    .auto_in_w_valid(dspQueue_auto_in_w_valid),
    .auto_in_w_bits_data(dspQueue_auto_in_w_bits_data),
    .auto_in_w_bits_strb(dspQueue_auto_in_w_bits_strb),
    .auto_in_b_ready(dspQueue_auto_in_b_ready),
    .auto_in_b_valid(dspQueue_auto_in_b_valid),
    .auto_in_b_bits_id(dspQueue_auto_in_b_bits_id),
    .auto_in_ar_ready(dspQueue_auto_in_ar_ready),
    .auto_in_ar_valid(dspQueue_auto_in_ar_valid),
    .auto_in_ar_bits_id(dspQueue_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(dspQueue_auto_in_ar_bits_addr),
    .auto_in_ar_bits_size(dspQueue_auto_in_ar_bits_size),
    .auto_in_r_ready(dspQueue_auto_in_r_ready),
    .auto_in_r_valid(dspQueue_auto_in_r_valid),
    .auto_in_r_bits_id(dspQueue_auto_in_r_bits_id),
    .auto_in_r_bits_data(dspQueue_auto_in_r_bits_data)
  );
  AXI4Xbar_1 bus ( // @[AccChain.scala 44:23]
    .clock(bus_clock),
    .reset(bus_reset),
    .auto_in_aw_ready(bus_auto_in_aw_ready),
    .auto_in_aw_valid(bus_auto_in_aw_valid),
    .auto_in_aw_bits_id(bus_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(bus_auto_in_aw_bits_addr),
    .auto_in_aw_bits_size(bus_auto_in_aw_bits_size),
    .auto_in_w_ready(bus_auto_in_w_ready),
    .auto_in_w_valid(bus_auto_in_w_valid),
    .auto_in_w_bits_data(bus_auto_in_w_bits_data),
    .auto_in_w_bits_strb(bus_auto_in_w_bits_strb),
    .auto_in_w_bits_last(bus_auto_in_w_bits_last),
    .auto_in_b_ready(bus_auto_in_b_ready),
    .auto_in_b_valid(bus_auto_in_b_valid),
    .auto_in_b_bits_resp(bus_auto_in_b_bits_resp),
    .auto_in_ar_ready(bus_auto_in_ar_ready),
    .auto_in_ar_valid(bus_auto_in_ar_valid),
    .auto_in_ar_bits_id(bus_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(bus_auto_in_ar_bits_addr),
    .auto_in_ar_bits_size(bus_auto_in_ar_bits_size),
    .auto_in_r_ready(bus_auto_in_r_ready),
    .auto_in_r_valid(bus_auto_in_r_valid),
    .auto_in_r_bits_data(bus_auto_in_r_bits_data),
    .auto_in_r_bits_resp(bus_auto_in_r_bits_resp),
    .auto_in_r_bits_last(bus_auto_in_r_bits_last),
    .auto_out_1_aw_ready(bus_auto_out_1_aw_ready),
    .auto_out_1_aw_valid(bus_auto_out_1_aw_valid),
    .auto_out_1_aw_bits_id(bus_auto_out_1_aw_bits_id),
    .auto_out_1_aw_bits_addr(bus_auto_out_1_aw_bits_addr),
    .auto_out_1_aw_bits_size(bus_auto_out_1_aw_bits_size),
    .auto_out_1_w_ready(bus_auto_out_1_w_ready),
    .auto_out_1_w_valid(bus_auto_out_1_w_valid),
    .auto_out_1_w_bits_data(bus_auto_out_1_w_bits_data),
    .auto_out_1_w_bits_strb(bus_auto_out_1_w_bits_strb),
    .auto_out_1_w_bits_last(bus_auto_out_1_w_bits_last),
    .auto_out_1_b_ready(bus_auto_out_1_b_ready),
    .auto_out_1_b_valid(bus_auto_out_1_b_valid),
    .auto_out_1_b_bits_id(bus_auto_out_1_b_bits_id),
    .auto_out_1_b_bits_resp(bus_auto_out_1_b_bits_resp),
    .auto_out_1_ar_ready(bus_auto_out_1_ar_ready),
    .auto_out_1_ar_valid(bus_auto_out_1_ar_valid),
    .auto_out_1_ar_bits_id(bus_auto_out_1_ar_bits_id),
    .auto_out_1_ar_bits_addr(bus_auto_out_1_ar_bits_addr),
    .auto_out_1_ar_bits_size(bus_auto_out_1_ar_bits_size),
    .auto_out_1_r_ready(bus_auto_out_1_r_ready),
    .auto_out_1_r_valid(bus_auto_out_1_r_valid),
    .auto_out_1_r_bits_id(bus_auto_out_1_r_bits_id),
    .auto_out_1_r_bits_data(bus_auto_out_1_r_bits_data),
    .auto_out_1_r_bits_resp(bus_auto_out_1_r_bits_resp),
    .auto_out_1_r_bits_last(bus_auto_out_1_r_bits_last),
    .auto_out_0_aw_ready(bus_auto_out_0_aw_ready),
    .auto_out_0_aw_valid(bus_auto_out_0_aw_valid),
    .auto_out_0_aw_bits_id(bus_auto_out_0_aw_bits_id),
    .auto_out_0_aw_bits_addr(bus_auto_out_0_aw_bits_addr),
    .auto_out_0_aw_bits_size(bus_auto_out_0_aw_bits_size),
    .auto_out_0_w_ready(bus_auto_out_0_w_ready),
    .auto_out_0_w_valid(bus_auto_out_0_w_valid),
    .auto_out_0_w_bits_data(bus_auto_out_0_w_bits_data),
    .auto_out_0_w_bits_strb(bus_auto_out_0_w_bits_strb),
    .auto_out_0_w_bits_last(bus_auto_out_0_w_bits_last),
    .auto_out_0_b_ready(bus_auto_out_0_b_ready),
    .auto_out_0_b_valid(bus_auto_out_0_b_valid),
    .auto_out_0_b_bits_id(bus_auto_out_0_b_bits_id),
    .auto_out_0_b_bits_resp(bus_auto_out_0_b_bits_resp),
    .auto_out_0_ar_ready(bus_auto_out_0_ar_ready),
    .auto_out_0_ar_valid(bus_auto_out_0_ar_valid),
    .auto_out_0_ar_bits_id(bus_auto_out_0_ar_bits_id),
    .auto_out_0_ar_bits_addr(bus_auto_out_0_ar_bits_addr),
    .auto_out_0_ar_bits_size(bus_auto_out_0_ar_bits_size),
    .auto_out_0_r_ready(bus_auto_out_0_r_ready),
    .auto_out_0_r_valid(bus_auto_out_0_r_valid),
    .auto_out_0_r_bits_id(bus_auto_out_0_r_bits_id),
    .auto_out_0_r_bits_data(bus_auto_out_0_r_bits_data),
    .auto_out_0_r_bits_resp(bus_auto_out_0_r_bits_resp),
    .auto_out_0_r_bits_last(bus_auto_out_0_r_bits_last)
  );
  AXI4Buffer axi4buf ( // @[Buffer.scala 58:29]
    .clock(axi4buf_clock),
    .reset(axi4buf_reset),
    .auto_in_aw_ready(axi4buf_auto_in_aw_ready),
    .auto_in_aw_valid(axi4buf_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4buf_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4buf_auto_in_aw_bits_addr),
    .auto_in_aw_bits_size(axi4buf_auto_in_aw_bits_size),
    .auto_in_w_ready(axi4buf_auto_in_w_ready),
    .auto_in_w_valid(axi4buf_auto_in_w_valid),
    .auto_in_w_bits_data(axi4buf_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi4buf_auto_in_w_bits_strb),
    .auto_in_w_bits_last(axi4buf_auto_in_w_bits_last),
    .auto_in_b_ready(axi4buf_auto_in_b_ready),
    .auto_in_b_valid(axi4buf_auto_in_b_valid),
    .auto_in_b_bits_id(axi4buf_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi4buf_auto_in_b_bits_resp),
    .auto_in_ar_ready(axi4buf_auto_in_ar_ready),
    .auto_in_ar_valid(axi4buf_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4buf_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4buf_auto_in_ar_bits_addr),
    .auto_in_ar_bits_size(axi4buf_auto_in_ar_bits_size),
    .auto_in_r_ready(axi4buf_auto_in_r_ready),
    .auto_in_r_valid(axi4buf_auto_in_r_valid),
    .auto_in_r_bits_id(axi4buf_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4buf_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4buf_auto_in_r_bits_resp),
    .auto_in_r_bits_last(axi4buf_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4buf_auto_out_aw_ready),
    .auto_out_aw_valid(axi4buf_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4buf_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4buf_auto_out_aw_bits_addr),
    .auto_out_w_ready(axi4buf_auto_out_w_ready),
    .auto_out_w_valid(axi4buf_auto_out_w_valid),
    .auto_out_w_bits_data(axi4buf_auto_out_w_bits_data),
    .auto_out_w_bits_strb(axi4buf_auto_out_w_bits_strb),
    .auto_out_w_bits_last(axi4buf_auto_out_w_bits_last),
    .auto_out_b_ready(axi4buf_auto_out_b_ready),
    .auto_out_b_valid(axi4buf_auto_out_b_valid),
    .auto_out_b_bits_id(axi4buf_auto_out_b_bits_id),
    .auto_out_b_bits_resp(axi4buf_auto_out_b_bits_resp),
    .auto_out_ar_ready(axi4buf_auto_out_ar_ready),
    .auto_out_ar_valid(axi4buf_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4buf_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4buf_auto_out_ar_bits_addr),
    .auto_out_ar_bits_size(axi4buf_auto_out_ar_bits_size),
    .auto_out_r_ready(axi4buf_auto_out_r_ready),
    .auto_out_r_valid(axi4buf_auto_out_r_valid),
    .auto_out_r_bits_id(axi4buf_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4buf_auto_out_r_bits_data),
    .auto_out_r_bits_resp(axi4buf_auto_out_r_bits_resp),
    .auto_out_r_bits_last(axi4buf_auto_out_r_bits_last)
  );
  AXI4Buffer axi4buf_1 ( // @[Buffer.scala 58:29]
    .clock(axi4buf_1_clock),
    .reset(axi4buf_1_reset),
    .auto_in_aw_ready(axi4buf_1_auto_in_aw_ready),
    .auto_in_aw_valid(axi4buf_1_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4buf_1_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4buf_1_auto_in_aw_bits_addr),
    .auto_in_aw_bits_size(axi4buf_1_auto_in_aw_bits_size),
    .auto_in_w_ready(axi4buf_1_auto_in_w_ready),
    .auto_in_w_valid(axi4buf_1_auto_in_w_valid),
    .auto_in_w_bits_data(axi4buf_1_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi4buf_1_auto_in_w_bits_strb),
    .auto_in_w_bits_last(axi4buf_1_auto_in_w_bits_last),
    .auto_in_b_ready(axi4buf_1_auto_in_b_ready),
    .auto_in_b_valid(axi4buf_1_auto_in_b_valid),
    .auto_in_b_bits_id(axi4buf_1_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi4buf_1_auto_in_b_bits_resp),
    .auto_in_ar_ready(axi4buf_1_auto_in_ar_ready),
    .auto_in_ar_valid(axi4buf_1_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4buf_1_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4buf_1_auto_in_ar_bits_addr),
    .auto_in_ar_bits_size(axi4buf_1_auto_in_ar_bits_size),
    .auto_in_r_ready(axi4buf_1_auto_in_r_ready),
    .auto_in_r_valid(axi4buf_1_auto_in_r_valid),
    .auto_in_r_bits_id(axi4buf_1_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4buf_1_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4buf_1_auto_in_r_bits_resp),
    .auto_in_r_bits_last(axi4buf_1_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4buf_1_auto_out_aw_ready),
    .auto_out_aw_valid(axi4buf_1_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4buf_1_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4buf_1_auto_out_aw_bits_addr),
    .auto_out_w_ready(axi4buf_1_auto_out_w_ready),
    .auto_out_w_valid(axi4buf_1_auto_out_w_valid),
    .auto_out_w_bits_data(axi4buf_1_auto_out_w_bits_data),
    .auto_out_w_bits_strb(axi4buf_1_auto_out_w_bits_strb),
    .auto_out_w_bits_last(axi4buf_1_auto_out_w_bits_last),
    .auto_out_b_ready(axi4buf_1_auto_out_b_ready),
    .auto_out_b_valid(axi4buf_1_auto_out_b_valid),
    .auto_out_b_bits_id(axi4buf_1_auto_out_b_bits_id),
    .auto_out_b_bits_resp(axi4buf_1_auto_out_b_bits_resp),
    .auto_out_ar_ready(axi4buf_1_auto_out_ar_ready),
    .auto_out_ar_valid(axi4buf_1_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4buf_1_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4buf_1_auto_out_ar_bits_addr),
    .auto_out_ar_bits_size(axi4buf_1_auto_out_ar_bits_size),
    .auto_out_r_ready(axi4buf_1_auto_out_r_ready),
    .auto_out_r_valid(axi4buf_1_auto_out_r_valid),
    .auto_out_r_bits_id(axi4buf_1_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4buf_1_auto_out_r_bits_data),
    .auto_out_r_bits_resp(axi4buf_1_auto_out_r_bits_resp),
    .auto_out_r_bits_last(axi4buf_1_auto_out_r_bits_last)
  );
  assign auto_bus_in_aw_ready = bus_auto_in_aw_ready; // @[LazyModule.scala 173:31]
  assign auto_bus_in_w_ready = bus_auto_in_w_ready; // @[LazyModule.scala 173:31]
  assign auto_bus_in_b_valid = bus_auto_in_b_valid; // @[LazyModule.scala 173:31]
  assign auto_bus_in_b_bits_resp = bus_auto_in_b_bits_resp; // @[LazyModule.scala 173:31]
  assign auto_bus_in_ar_ready = bus_auto_in_ar_ready; // @[LazyModule.scala 173:31]
  assign auto_bus_in_r_valid = bus_auto_in_r_valid; // @[LazyModule.scala 173:31]
  assign auto_bus_in_r_bits_data = bus_auto_in_r_bits_data; // @[LazyModule.scala 173:31]
  assign auto_bus_in_r_bits_resp = bus_auto_in_r_bits_resp; // @[LazyModule.scala 173:31]
  assign auto_bus_in_r_bits_last = bus_auto_in_r_bits_last; // @[LazyModule.scala 173:31]
  assign auto_dspQueue_stream_out_valid = dspQueue_auto_stream_out_valid; // @[LazyModule.scala 173:49]
  assign auto_dspQueue_stream_out_bits_data = dspQueue_auto_stream_out_bits_data; // @[LazyModule.scala 173:49]
  assign auto_dspQueue_stream_out_bits_last = dspQueue_auto_stream_out_bits_last; // @[LazyModule.scala 173:49]
  assign auto_accumulator_slave_in_ready = accumulator_auto_slave_in_ready; // @[LazyModule.scala 173:31]
  assign accumulator_clock = clock;
  assign accumulator_reset = reset;
  assign accumulator_auto_mem_in_aw_valid = axi4buf_1_auto_out_aw_valid; // @[LazyModule.scala 167:31]
  assign accumulator_auto_mem_in_aw_bits_id = axi4buf_1_auto_out_aw_bits_id; // @[LazyModule.scala 167:31]
  assign accumulator_auto_mem_in_aw_bits_addr = axi4buf_1_auto_out_aw_bits_addr; // @[LazyModule.scala 167:31]
  assign accumulator_auto_mem_in_w_valid = axi4buf_1_auto_out_w_valid; // @[LazyModule.scala 167:31]
  assign accumulator_auto_mem_in_w_bits_data = axi4buf_1_auto_out_w_bits_data; // @[LazyModule.scala 167:31]
  assign accumulator_auto_mem_in_w_bits_strb = axi4buf_1_auto_out_w_bits_strb; // @[LazyModule.scala 167:31]
  assign accumulator_auto_mem_in_b_ready = axi4buf_1_auto_out_b_ready; // @[LazyModule.scala 167:31]
  assign accumulator_auto_mem_in_ar_valid = axi4buf_1_auto_out_ar_valid; // @[LazyModule.scala 167:31]
  assign accumulator_auto_mem_in_ar_bits_id = axi4buf_1_auto_out_ar_bits_id; // @[LazyModule.scala 167:31]
  assign accumulator_auto_mem_in_ar_bits_addr = axi4buf_1_auto_out_ar_bits_addr; // @[LazyModule.scala 167:31]
  assign accumulator_auto_mem_in_ar_bits_size = axi4buf_1_auto_out_ar_bits_size; // @[LazyModule.scala 167:31]
  assign accumulator_auto_mem_in_r_ready = axi4buf_1_auto_out_r_ready; // @[LazyModule.scala 167:31]
  assign accumulator_auto_master_out_ready = dspQueue_auto_stream_in_ready; // @[LazyModule.scala 167:57]
  assign accumulator_auto_slave_in_valid = auto_accumulator_slave_in_valid; // @[LazyModule.scala 173:31]
  assign accumulator_auto_slave_in_bits_data = auto_accumulator_slave_in_bits_data; // @[LazyModule.scala 173:31]
  assign accumulator_auto_slave_in_bits_last = auto_accumulator_slave_in_bits_last; // @[LazyModule.scala 173:31]
  assign dspQueue_clock = clock;
  assign dspQueue_reset = reset;
  assign dspQueue_auto_stream_in_valid = accumulator_auto_master_out_valid; // @[LazyModule.scala 167:57]
  assign dspQueue_auto_stream_in_bits_data = accumulator_auto_master_out_bits_data; // @[LazyModule.scala 167:57]
  assign dspQueue_auto_stream_in_bits_last = accumulator_auto_master_out_bits_last; // @[LazyModule.scala 167:57]
  assign dspQueue_auto_stream_out_ready = auto_dspQueue_stream_out_ready; // @[LazyModule.scala 173:49]
  assign dspQueue_auto_in_aw_valid = axi4buf_auto_out_aw_valid; // @[LazyModule.scala 167:31]
  assign dspQueue_auto_in_aw_bits_id = axi4buf_auto_out_aw_bits_id; // @[LazyModule.scala 167:31]
  assign dspQueue_auto_in_aw_bits_addr = axi4buf_auto_out_aw_bits_addr; // @[LazyModule.scala 167:31]
  assign dspQueue_auto_in_w_valid = axi4buf_auto_out_w_valid; // @[LazyModule.scala 167:31]
  assign dspQueue_auto_in_w_bits_data = axi4buf_auto_out_w_bits_data; // @[LazyModule.scala 167:31]
  assign dspQueue_auto_in_w_bits_strb = axi4buf_auto_out_w_bits_strb; // @[LazyModule.scala 167:31]
  assign dspQueue_auto_in_b_ready = axi4buf_auto_out_b_ready; // @[LazyModule.scala 167:31]
  assign dspQueue_auto_in_ar_valid = axi4buf_auto_out_ar_valid; // @[LazyModule.scala 167:31]
  assign dspQueue_auto_in_ar_bits_id = axi4buf_auto_out_ar_bits_id; // @[LazyModule.scala 167:31]
  assign dspQueue_auto_in_ar_bits_addr = axi4buf_auto_out_ar_bits_addr; // @[LazyModule.scala 167:31]
  assign dspQueue_auto_in_ar_bits_size = axi4buf_auto_out_ar_bits_size; // @[LazyModule.scala 167:31]
  assign dspQueue_auto_in_r_ready = axi4buf_auto_out_r_ready; // @[LazyModule.scala 167:31]
  assign bus_clock = clock;
  assign bus_reset = reset;
  assign bus_auto_in_aw_valid = auto_bus_in_aw_valid; // @[LazyModule.scala 173:31]
  assign bus_auto_in_aw_bits_id = auto_bus_in_aw_bits_id; // @[LazyModule.scala 173:31]
  assign bus_auto_in_aw_bits_addr = auto_bus_in_aw_bits_addr; // @[LazyModule.scala 173:31]
  assign bus_auto_in_aw_bits_size = auto_bus_in_aw_bits_size; // @[LazyModule.scala 173:31]
  assign bus_auto_in_w_valid = auto_bus_in_w_valid; // @[LazyModule.scala 173:31]
  assign bus_auto_in_w_bits_data = auto_bus_in_w_bits_data; // @[LazyModule.scala 173:31]
  assign bus_auto_in_w_bits_strb = auto_bus_in_w_bits_strb; // @[LazyModule.scala 173:31]
  assign bus_auto_in_w_bits_last = auto_bus_in_w_bits_last; // @[LazyModule.scala 173:31]
  assign bus_auto_in_b_ready = auto_bus_in_b_ready; // @[LazyModule.scala 173:31]
  assign bus_auto_in_ar_valid = auto_bus_in_ar_valid; // @[LazyModule.scala 173:31]
  assign bus_auto_in_ar_bits_id = auto_bus_in_ar_bits_id; // @[LazyModule.scala 173:31]
  assign bus_auto_in_ar_bits_addr = auto_bus_in_ar_bits_addr; // @[LazyModule.scala 173:31]
  assign bus_auto_in_ar_bits_size = auto_bus_in_ar_bits_size; // @[LazyModule.scala 173:31]
  assign bus_auto_in_r_ready = auto_bus_in_r_ready; // @[LazyModule.scala 173:31]
  assign bus_auto_out_1_aw_ready = axi4buf_1_auto_in_aw_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_1_w_ready = axi4buf_1_auto_in_w_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_1_b_valid = axi4buf_1_auto_in_b_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_1_b_bits_id = axi4buf_1_auto_in_b_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_1_b_bits_resp = axi4buf_1_auto_in_b_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_1_ar_ready = axi4buf_1_auto_in_ar_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_1_r_valid = axi4buf_1_auto_in_r_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_1_r_bits_id = axi4buf_1_auto_in_r_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_1_r_bits_data = axi4buf_1_auto_in_r_bits_data; // @[LazyModule.scala 167:57]
  assign bus_auto_out_1_r_bits_resp = axi4buf_1_auto_in_r_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_1_r_bits_last = axi4buf_1_auto_in_r_bits_last; // @[LazyModule.scala 167:57]
  assign bus_auto_out_0_aw_ready = axi4buf_auto_in_aw_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_0_w_ready = axi4buf_auto_in_w_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_0_b_valid = axi4buf_auto_in_b_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_0_b_bits_id = axi4buf_auto_in_b_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_0_b_bits_resp = axi4buf_auto_in_b_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_0_ar_ready = axi4buf_auto_in_ar_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_0_r_valid = axi4buf_auto_in_r_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_0_r_bits_id = axi4buf_auto_in_r_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_0_r_bits_data = axi4buf_auto_in_r_bits_data; // @[LazyModule.scala 167:57]
  assign bus_auto_out_0_r_bits_resp = axi4buf_auto_in_r_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_0_r_bits_last = axi4buf_auto_in_r_bits_last; // @[LazyModule.scala 167:57]
  assign axi4buf_clock = clock;
  assign axi4buf_reset = reset;
  assign axi4buf_auto_in_aw_valid = bus_auto_out_0_aw_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_auto_in_aw_bits_id = bus_auto_out_0_aw_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_auto_in_aw_bits_addr = bus_auto_out_0_aw_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_auto_in_aw_bits_size = bus_auto_out_0_aw_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_auto_in_w_valid = bus_auto_out_0_w_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_auto_in_w_bits_data = bus_auto_out_0_w_bits_data; // @[LazyModule.scala 167:57]
  assign axi4buf_auto_in_w_bits_strb = bus_auto_out_0_w_bits_strb; // @[LazyModule.scala 167:57]
  assign axi4buf_auto_in_w_bits_last = bus_auto_out_0_w_bits_last; // @[LazyModule.scala 167:57]
  assign axi4buf_auto_in_b_ready = bus_auto_out_0_b_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_auto_in_ar_valid = bus_auto_out_0_ar_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_auto_in_ar_bits_id = bus_auto_out_0_ar_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_auto_in_ar_bits_addr = bus_auto_out_0_ar_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_auto_in_ar_bits_size = bus_auto_out_0_ar_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_auto_in_r_ready = bus_auto_out_0_r_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_auto_out_aw_ready = dspQueue_auto_in_aw_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_auto_out_w_ready = dspQueue_auto_in_w_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_auto_out_b_valid = dspQueue_auto_in_b_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_auto_out_b_bits_id = dspQueue_auto_in_b_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_auto_out_b_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_auto_out_ar_ready = dspQueue_auto_in_ar_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_auto_out_r_valid = dspQueue_auto_in_r_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_auto_out_r_bits_id = dspQueue_auto_in_r_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_auto_out_r_bits_data = dspQueue_auto_in_r_bits_data; // @[LazyModule.scala 167:31]
  assign axi4buf_auto_out_r_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_auto_out_r_bits_last = 1'h1; // @[LazyModule.scala 167:31]
  assign axi4buf_1_clock = clock;
  assign axi4buf_1_reset = reset;
  assign axi4buf_1_auto_in_aw_valid = bus_auto_out_1_aw_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_1_auto_in_aw_bits_id = bus_auto_out_1_aw_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_1_auto_in_aw_bits_addr = bus_auto_out_1_aw_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_1_auto_in_aw_bits_size = bus_auto_out_1_aw_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_1_auto_in_w_valid = bus_auto_out_1_w_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_1_auto_in_w_bits_data = bus_auto_out_1_w_bits_data; // @[LazyModule.scala 167:57]
  assign axi4buf_1_auto_in_w_bits_strb = bus_auto_out_1_w_bits_strb; // @[LazyModule.scala 167:57]
  assign axi4buf_1_auto_in_w_bits_last = bus_auto_out_1_w_bits_last; // @[LazyModule.scala 167:57]
  assign axi4buf_1_auto_in_b_ready = bus_auto_out_1_b_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_1_auto_in_ar_valid = bus_auto_out_1_ar_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_1_auto_in_ar_bits_id = bus_auto_out_1_ar_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_1_auto_in_ar_bits_addr = bus_auto_out_1_ar_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_1_auto_in_ar_bits_size = bus_auto_out_1_ar_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_1_auto_in_r_ready = bus_auto_out_1_r_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_1_auto_out_aw_ready = accumulator_auto_mem_in_aw_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_1_auto_out_w_ready = accumulator_auto_mem_in_w_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_1_auto_out_b_valid = accumulator_auto_mem_in_b_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_1_auto_out_b_bits_id = accumulator_auto_mem_in_b_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_1_auto_out_b_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_1_auto_out_ar_ready = accumulator_auto_mem_in_ar_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_1_auto_out_r_valid = accumulator_auto_mem_in_r_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_1_auto_out_r_bits_id = accumulator_auto_mem_in_r_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_1_auto_out_r_bits_data = accumulator_auto_mem_in_r_bits_data; // @[LazyModule.scala 167:31]
  assign axi4buf_1_auto_out_r_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_1_auto_out_r_bits_last = 1'h1; // @[LazyModule.scala 167:31]
endmodule
module AXI4StreamWidthAdapater_2_to_1(
  input         clock,
  input         reset,
  output        auto_in_ready,
  input         auto_in_valid,
  input  [15:0] auto_in_bits_data,
  input         auto_in_bits_last,
  input         auto_out_ready,
  output        auto_out_valid,
  output [31:0] auto_out_bits_data,
  output        auto_out_bits_last
);
  reg [15:0] _T; // @[AXI4StreamWidthAdapter.scala 101:37]
  reg [31:0] _RAND_0;
  reg  _T_1; // @[AXI4StreamWidthAdapter.scala 102:22]
  reg [31:0] _RAND_1;
  wire  _T_2 = auto_in_valid & auto_out_ready; // @[AXI4StreamWidthAdapter.scala 103:14]
  wire [1:0] _T_4 = _T_1 + 1'h1; // @[AXI4StreamWidthAdapter.scala 103:60]
  wire [1:0] _T_5 = _T_1 ? 2'h0 : _T_4; // @[AXI4StreamWidthAdapter.scala 103:33]
  wire [1:0] _GEN_0 = _T_2 ? _T_5 : {{1'd0}, _T_1}; // @[AXI4StreamWidthAdapter.scala 103:21]
  wire  _T_7 = ~_T_1; // @[AXI4StreamWidthAdapter.scala 106:29]
  wire  _T_8 = _T_2 & _T_7; // @[AXI4StreamWidthAdapter.scala 106:22]
  wire  ov0 = _T_1 & auto_in_valid; // @[AXI4StreamWidthAdapter.scala 112:32]
  reg  _T_10; // @[AXI4StreamWidthAdapter.scala 101:37]
  reg [31:0] _RAND_2;
  reg  _T_11; // @[AXI4StreamWidthAdapter.scala 102:22]
  reg [31:0] _RAND_3;
  wire [1:0] _T_14 = _T_11 + 1'h1; // @[AXI4StreamWidthAdapter.scala 103:60]
  wire [1:0] _T_15 = _T_11 ? 2'h0 : _T_14; // @[AXI4StreamWidthAdapter.scala 103:33]
  wire [1:0] _GEN_2 = _T_2 ? _T_15 : {{1'd0}, _T_11}; // @[AXI4StreamWidthAdapter.scala 103:21]
  wire  _T_17 = ~_T_11; // @[AXI4StreamWidthAdapter.scala 106:29]
  wire  _T_18 = _T_2 & _T_17; // @[AXI4StreamWidthAdapter.scala 106:22]
  wire [1:0] _T_19 = {auto_in_bits_last,_T_10}; // @[Cat.scala 29:58]
  wire  ov1 = _T_11 & auto_in_valid; // @[AXI4StreamWidthAdapter.scala 112:32]
  reg  _T_22; // @[AXI4StreamWidthAdapter.scala 102:22]
  reg [31:0] _RAND_4;
  wire [1:0] _T_25 = _T_22 + 1'h1; // @[AXI4StreamWidthAdapter.scala 103:60]
  wire [1:0] _T_26 = _T_22 ? 2'h0 : _T_25; // @[AXI4StreamWidthAdapter.scala 103:33]
  wire [1:0] _GEN_4 = _T_2 ? _T_26 : {{1'd0}, _T_22}; // @[AXI4StreamWidthAdapter.scala 103:21]
  wire  ov2 = _T_22 & auto_in_valid; // @[AXI4StreamWidthAdapter.scala 112:32]
  reg  _T_32; // @[AXI4StreamWidthAdapter.scala 102:22]
  reg [31:0] _RAND_5;
  wire [1:0] _T_35 = _T_32 + 1'h1; // @[AXI4StreamWidthAdapter.scala 103:60]
  wire [1:0] _T_36 = _T_32 ? 2'h0 : _T_35; // @[AXI4StreamWidthAdapter.scala 103:33]
  wire [1:0] _GEN_6 = _T_2 ? _T_36 : {{1'd0}, _T_32}; // @[AXI4StreamWidthAdapter.scala 103:21]
  wire  ov3 = _T_32 & auto_in_valid; // @[AXI4StreamWidthAdapter.scala 112:32]
  reg  _T_42; // @[AXI4StreamWidthAdapter.scala 102:22]
  reg [31:0] _RAND_6;
  wire [1:0] _T_45 = _T_42 + 1'h1; // @[AXI4StreamWidthAdapter.scala 103:60]
  wire [1:0] _T_46 = _T_42 ? 2'h0 : _T_45; // @[AXI4StreamWidthAdapter.scala 103:33]
  wire [1:0] _GEN_8 = _T_2 ? _T_46 : {{1'd0}, _T_42}; // @[AXI4StreamWidthAdapter.scala 103:21]
  wire  ov4 = _T_42 & auto_in_valid; // @[AXI4StreamWidthAdapter.scala 112:32]
  wire  _T_51 = ov0 == ov1; // @[AXI4StreamWidthAdapter.scala 42:16]
  wire  _T_53 = _T_51 | reset; // @[AXI4StreamWidthAdapter.scala 42:11]
  wire  _T_54 = ~_T_53; // @[AXI4StreamWidthAdapter.scala 42:11]
  wire  _T_55 = ov0 == ov2; // @[AXI4StreamWidthAdapter.scala 43:16]
  wire  _T_57 = _T_55 | reset; // @[AXI4StreamWidthAdapter.scala 43:11]
  wire  _T_58 = ~_T_57; // @[AXI4StreamWidthAdapter.scala 43:11]
  wire  _T_59 = ov0 == ov3; // @[AXI4StreamWidthAdapter.scala 44:16]
  wire  _T_61 = _T_59 | reset; // @[AXI4StreamWidthAdapter.scala 44:11]
  wire  _T_62 = ~_T_61; // @[AXI4StreamWidthAdapter.scala 44:11]
  wire  _T_63 = ov0 == ov4; // @[AXI4StreamWidthAdapter.scala 45:16]
  wire  _T_65 = _T_63 | reset; // @[AXI4StreamWidthAdapter.scala 45:11]
  wire  _T_66 = ~_T_65; // @[AXI4StreamWidthAdapter.scala 45:11]
  assign auto_in_ready = auto_out_ready; // @[LazyModule.scala 173:31]
  assign auto_out_valid = _T_1 & auto_in_valid; // @[LazyModule.scala 173:49]
  assign auto_out_bits_data = {auto_in_bits_data,_T}; // @[LazyModule.scala 173:49]
  assign auto_out_bits_last = _T_19 != 2'h0; // @[LazyModule.scala 173:49]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_10 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_11 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_22 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_32 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_42 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (_T_8) begin
      _T <= auto_in_bits_data;
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else begin
      _T_1 <= _GEN_0[0];
    end
    if (_T_18) begin
      _T_10 <= auto_in_bits_last;
    end
    if (reset) begin
      _T_11 <= 1'h0;
    end else begin
      _T_11 <= _GEN_2[0];
    end
    if (reset) begin
      _T_22 <= 1'h0;
    end else begin
      _T_22 <= _GEN_4[0];
    end
    if (reset) begin
      _T_32 <= 1'h0;
    end else begin
      _T_32 <= _GEN_6[0];
    end
    if (reset) begin
      _T_42 <= 1'h0;
    end else begin
      _T_42 <= _GEN_8[0];
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_54) begin
          $fwrite(32'h80000002,"Assertion failed\n    at AXI4StreamWidthAdapter.scala:42 assert(ov0 === ov1)\n"); // @[AXI4StreamWidthAdapter.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_54) begin
          $fatal; // @[AXI4StreamWidthAdapter.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_58) begin
          $fwrite(32'h80000002,"Assertion failed\n    at AXI4StreamWidthAdapter.scala:43 assert(ov0 === ov2)\n"); // @[AXI4StreamWidthAdapter.scala 43:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_58) begin
          $fatal; // @[AXI4StreamWidthAdapter.scala 43:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_62) begin
          $fwrite(32'h80000002,"Assertion failed\n    at AXI4StreamWidthAdapter.scala:44 assert(ov0 === ov3)\n"); // @[AXI4StreamWidthAdapter.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_62) begin
          $fatal; // @[AXI4StreamWidthAdapter.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_66) begin
          $fwrite(32'h80000002,"Assertion failed\n    at AXI4StreamWidthAdapter.scala:45 assert(ov0 === ov4)\n"); // @[AXI4StreamWidthAdapter.scala 45:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_66) begin
          $fatal; // @[AXI4StreamWidthAdapter.scala 45:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module Queue_35(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [31:0] io_enq_bits_data,
  input         io_enq_bits_last,
  input         io_deq_ready,
  output        io_deq_valid,
  output [31:0] io_deq_bits_data,
  output        io_deq_bits_last
);
  reg [31:0] _T_data [0:0]; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_0;
  wire [31:0] _T_data__T_14_data; // @[Decoupled.scala 218:24]
  wire  _T_data__T_14_addr; // @[Decoupled.scala 218:24]
  wire [31:0] _T_data__T_10_data; // @[Decoupled.scala 218:24]
  wire  _T_data__T_10_addr; // @[Decoupled.scala 218:24]
  wire  _T_data__T_10_mask; // @[Decoupled.scala 218:24]
  wire  _T_data__T_10_en; // @[Decoupled.scala 218:24]
  reg  _T_last [0:0]; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_1;
  wire  _T_last__T_14_data; // @[Decoupled.scala 218:24]
  wire  _T_last__T_14_addr; // @[Decoupled.scala 218:24]
  wire  _T_last__T_10_data; // @[Decoupled.scala 218:24]
  wire  _T_last__T_10_addr; // @[Decoupled.scala 218:24]
  wire  _T_last__T_10_mask; // @[Decoupled.scala 218:24]
  wire  _T_last__T_10_en; // @[Decoupled.scala 218:24]
  reg  _T_1; // @[Decoupled.scala 221:35]
  reg [31:0] _RAND_2;
  wire  _T_3 = ~_T_1; // @[Decoupled.scala 224:36]
  wire  _T_6 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  _T_8 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_13 = io_deq_ready ? 1'h0 : _T_6; // @[Decoupled.scala 249:27]
  wire  _GEN_22 = _T_3 ? _GEN_13 : _T_6; // @[Decoupled.scala 246:18]
  wire  _GEN_21 = _T_3 ? 1'h0 : _T_8; // @[Decoupled.scala 246:18]
  wire  _T_11 = _GEN_22 != _GEN_21; // @[Decoupled.scala 236:16]
  wire  _T_12 = ~_T_3; // @[Decoupled.scala 240:19]
  assign _T_data__T_14_addr = 1'h0;
  assign _T_data__T_14_data = _T_data[_T_data__T_14_addr]; // @[Decoupled.scala 218:24]
  assign _T_data__T_10_data = io_enq_bits_data;
  assign _T_data__T_10_addr = 1'h0;
  assign _T_data__T_10_mask = 1'h1;
  assign _T_data__T_10_en = _T_3 ? _GEN_13 : _T_6;
  assign _T_last__T_14_addr = 1'h0;
  assign _T_last__T_14_data = _T_last[_T_last__T_14_addr]; // @[Decoupled.scala 218:24]
  assign _T_last__T_10_data = io_enq_bits_last;
  assign _T_last__T_10_addr = 1'h0;
  assign _T_last__T_10_mask = 1'h1;
  assign _T_last__T_10_en = _T_3 ? _GEN_13 : _T_6;
  assign io_enq_ready = io_deq_ready | _T_3; // @[Decoupled.scala 241:16 Decoupled.scala 254:40]
  assign io_deq_valid = io_enq_valid | _T_12; // @[Decoupled.scala 240:16 Decoupled.scala 245:40]
  assign io_deq_bits_data = _T_3 ? io_enq_bits_data : _T_data__T_14_data; // @[Decoupled.scala 242:15 Decoupled.scala 247:19]
  assign io_deq_bits_last = _T_3 ? io_enq_bits_last : _T_last__T_14_data; // @[Decoupled.scala 242:15 Decoupled.scala 247:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_data[initvar] = _RAND_0[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_last[initvar] = _RAND_1[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_1 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T_data__T_10_en & _T_data__T_10_mask) begin
      _T_data[_T_data__T_10_addr] <= _T_data__T_10_data; // @[Decoupled.scala 218:24]
    end
    if(_T_last__T_10_en & _T_last__T_10_mask) begin
      _T_last[_T_last__T_10_addr] <= _T_last__T_10_data; // @[Decoupled.scala 218:24]
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else if (_T_11) begin
      if (_T_3) begin
        if (io_deq_ready) begin
          _T_1 <= 1'h0;
        end else begin
          _T_1 <= _T_6;
        end
      end else begin
        _T_1 <= _T_6;
      end
    end
  end
endmodule
module StreamBuffer_1(
  input         clock,
  input         reset,
  input         auto_out_out_ready,
  output        auto_out_out_valid,
  output [31:0] auto_out_out_bits_data,
  output        auto_out_out_bits_last,
  output        auto_in_in_ready,
  input         auto_in_in_valid,
  input  [31:0] auto_in_in_bits_data,
  input         auto_in_in_bits_last
);
  wire  Queue_clock; // @[Decoupled.scala 296:21]
  wire  Queue_reset; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [31:0] Queue_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_bits_last; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [31:0] Queue_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_bits_last; // @[Decoupled.scala 296:21]
  Queue_35 Queue ( // @[Decoupled.scala 296:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_last(Queue_io_enq_bits_last),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_last(Queue_io_deq_bits_last)
  );
  assign auto_out_out_valid = Queue_io_deq_valid; // @[LazyModule.scala 173:49]
  assign auto_out_out_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_out_bits_last = Queue_io_deq_bits_last; // @[LazyModule.scala 173:49]
  assign auto_in_in_ready = Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_in_in_valid; // @[Decoupled.scala 297:22]
  assign Queue_io_enq_bits_data = auto_in_in_bits_data; // @[Decoupled.scala 298:21]
  assign Queue_io_enq_bits_last = auto_in_in_bits_last; // @[Decoupled.scala 298:21]
  assign Queue_io_deq_ready = auto_out_out_ready; // @[Decoupled.scala 320:15]
endmodule
module AXI4StreamMux_8(
  input         clock,
  input         reset,
  output        auto_register_in_aw_ready,
  input         auto_register_in_aw_valid,
  input         auto_register_in_aw_bits_id,
  input  [29:0] auto_register_in_aw_bits_addr,
  output        auto_register_in_w_ready,
  input         auto_register_in_w_valid,
  input  [31:0] auto_register_in_w_bits_data,
  input  [3:0]  auto_register_in_w_bits_strb,
  input         auto_register_in_b_ready,
  output        auto_register_in_b_valid,
  output        auto_register_in_b_bits_id,
  output        auto_register_in_ar_ready,
  input         auto_register_in_ar_valid,
  input         auto_register_in_ar_bits_id,
  input  [29:0] auto_register_in_ar_bits_addr,
  input  [2:0]  auto_register_in_ar_bits_size,
  input         auto_register_in_r_ready,
  output        auto_register_in_r_valid,
  output        auto_register_in_r_bits_id,
  output [31:0] auto_register_in_r_bits_data,
  output        auto_stream_in_6_ready,
  input         auto_stream_in_6_valid,
  input  [31:0] auto_stream_in_6_bits_data,
  input         auto_stream_in_6_bits_last,
  output        auto_stream_in_5_ready,
  input         auto_stream_in_5_valid,
  input  [31:0] auto_stream_in_5_bits_data,
  input         auto_stream_in_5_bits_last,
  output        auto_stream_in_4_ready,
  input         auto_stream_in_4_valid,
  input  [31:0] auto_stream_in_4_bits_data,
  input         auto_stream_in_4_bits_last,
  output        auto_stream_in_3_ready,
  input         auto_stream_in_3_valid,
  input  [31:0] auto_stream_in_3_bits_data,
  input         auto_stream_in_3_bits_last,
  output        auto_stream_in_2_ready,
  input         auto_stream_in_2_valid,
  input  [31:0] auto_stream_in_2_bits_data,
  input         auto_stream_in_2_bits_last,
  output        auto_stream_in_1_ready,
  input         auto_stream_in_1_valid,
  input  [31:0] auto_stream_in_1_bits_data,
  input         auto_stream_in_1_bits_last,
  output        auto_stream_in_0_ready,
  input         auto_stream_in_0_valid,
  input  [31:0] auto_stream_in_0_bits_data,
  input         auto_stream_in_0_bits_last,
  input         auto_stream_out_1_ready,
  output        auto_stream_out_1_valid,
  output [31:0] auto_stream_out_1_bits_data,
  output        auto_stream_out_1_bits_last,
  input         auto_stream_out_0_ready,
  output        auto_stream_out_0_valid,
  output [31:0] auto_stream_out_0_bits_data,
  output        auto_stream_out_0_bits_last
);
  wire  Queue_clock; // @[Decoupled.scala 296:21]
  wire  Queue_reset; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_bits_read; // @[Decoupled.scala 296:21]
  wire [31:0] Queue_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_bits_extra; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_bits_read; // @[Decoupled.scala 296:21]
  wire [31:0] Queue_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_bits_extra; // @[Decoupled.scala 296:21]
  reg [2:0] sels_0; // @[Mux.scala 32:23]
  reg [31:0] _RAND_0;
  reg [2:0] sels_1; // @[Mux.scala 32:23]
  reg [31:0] _RAND_1;
  reg [2:0] sels_2; // @[Mux.scala 32:23]
  reg [31:0] _RAND_2;
  wire  _T_3 = sels_0 == 3'h0; // @[Mux.scala 45:28]
  wire  _GEN_7 = _T_3 & auto_stream_in_0_valid; // @[Mux.scala 45:41]
  wire  _GEN_8 = _T_3 & auto_stream_out_0_ready; // @[Mux.scala 45:41]
  wire  _T_4 = sels_0 == 3'h1; // @[Mux.scala 45:28]
  wire  _GEN_12 = _T_4 ? auto_stream_in_1_bits_last : auto_stream_in_0_bits_last; // @[Mux.scala 45:41]
  wire [31:0] _GEN_15 = _T_4 ? auto_stream_in_1_bits_data : auto_stream_in_0_bits_data; // @[Mux.scala 45:41]
  wire  _GEN_16 = _T_4 ? auto_stream_in_1_valid : _GEN_7; // @[Mux.scala 45:41]
  wire  _GEN_17 = _T_4 & auto_stream_out_0_ready; // @[Mux.scala 45:41]
  wire  _T_5 = sels_0 == 3'h2; // @[Mux.scala 45:28]
  wire  _GEN_21 = _T_5 ? auto_stream_in_2_bits_last : _GEN_12; // @[Mux.scala 45:41]
  wire [31:0] _GEN_24 = _T_5 ? auto_stream_in_2_bits_data : _GEN_15; // @[Mux.scala 45:41]
  wire  _GEN_25 = _T_5 ? auto_stream_in_2_valid : _GEN_16; // @[Mux.scala 45:41]
  wire  _GEN_26 = _T_5 & auto_stream_out_0_ready; // @[Mux.scala 45:41]
  wire  _T_6 = sels_0 == 3'h3; // @[Mux.scala 45:28]
  wire  _GEN_30 = _T_6 ? auto_stream_in_3_bits_last : _GEN_21; // @[Mux.scala 45:41]
  wire [31:0] _GEN_33 = _T_6 ? auto_stream_in_3_bits_data : _GEN_24; // @[Mux.scala 45:41]
  wire  _GEN_34 = _T_6 ? auto_stream_in_3_valid : _GEN_25; // @[Mux.scala 45:41]
  wire  _GEN_35 = _T_6 & auto_stream_out_0_ready; // @[Mux.scala 45:41]
  wire  _T_7 = sels_0 == 3'h4; // @[Mux.scala 45:28]
  wire  _GEN_39 = _T_7 ? auto_stream_in_4_bits_last : _GEN_30; // @[Mux.scala 45:41]
  wire [31:0] _GEN_42 = _T_7 ? auto_stream_in_4_bits_data : _GEN_33; // @[Mux.scala 45:41]
  wire  _GEN_43 = _T_7 ? auto_stream_in_4_valid : _GEN_34; // @[Mux.scala 45:41]
  wire  _GEN_44 = _T_7 & auto_stream_out_0_ready; // @[Mux.scala 45:41]
  wire  _T_8 = sels_0 == 3'h5; // @[Mux.scala 45:28]
  wire  _GEN_48 = _T_8 ? auto_stream_in_5_bits_last : _GEN_39; // @[Mux.scala 45:41]
  wire [31:0] _GEN_51 = _T_8 ? auto_stream_in_5_bits_data : _GEN_42; // @[Mux.scala 45:41]
  wire  _GEN_52 = _T_8 ? auto_stream_in_5_valid : _GEN_43; // @[Mux.scala 45:41]
  wire  _GEN_53 = _T_8 & auto_stream_out_0_ready; // @[Mux.scala 45:41]
  wire  _T_9 = sels_0 == 3'h6; // @[Mux.scala 45:28]
  wire  _GEN_62 = _T_9 & auto_stream_out_0_ready; // @[Mux.scala 45:41]
  wire  _T_10 = sels_0 == sels_1; // @[Mux.scala 40:46]
  wire [2:0] _T_12 = _T_10 ? 3'h7 : sels_1; // @[Mux.scala 41:29]
  wire  _T_13 = _T_12 == 3'h0; // @[Mux.scala 45:28]
  wire  _GEN_70 = _T_13 & auto_stream_in_0_valid; // @[Mux.scala 45:41]
  wire  _GEN_71 = _T_13 ? auto_stream_out_1_ready : _GEN_8; // @[Mux.scala 45:41]
  wire  _T_14 = _T_12 == 3'h1; // @[Mux.scala 45:28]
  wire  _GEN_75 = _T_14 ? auto_stream_in_1_bits_last : auto_stream_in_0_bits_last; // @[Mux.scala 45:41]
  wire [31:0] _GEN_78 = _T_14 ? auto_stream_in_1_bits_data : auto_stream_in_0_bits_data; // @[Mux.scala 45:41]
  wire  _GEN_79 = _T_14 ? auto_stream_in_1_valid : _GEN_70; // @[Mux.scala 45:41]
  wire  _GEN_80 = _T_14 ? auto_stream_out_1_ready : _GEN_17; // @[Mux.scala 45:41]
  wire  _T_15 = _T_12 == 3'h2; // @[Mux.scala 45:28]
  wire  _GEN_84 = _T_15 ? auto_stream_in_2_bits_last : _GEN_75; // @[Mux.scala 45:41]
  wire [31:0] _GEN_87 = _T_15 ? auto_stream_in_2_bits_data : _GEN_78; // @[Mux.scala 45:41]
  wire  _GEN_88 = _T_15 ? auto_stream_in_2_valid : _GEN_79; // @[Mux.scala 45:41]
  wire  _GEN_89 = _T_15 ? auto_stream_out_1_ready : _GEN_26; // @[Mux.scala 45:41]
  wire  _T_16 = _T_12 == 3'h3; // @[Mux.scala 45:28]
  wire  _GEN_93 = _T_16 ? auto_stream_in_3_bits_last : _GEN_84; // @[Mux.scala 45:41]
  wire [31:0] _GEN_96 = _T_16 ? auto_stream_in_3_bits_data : _GEN_87; // @[Mux.scala 45:41]
  wire  _GEN_97 = _T_16 ? auto_stream_in_3_valid : _GEN_88; // @[Mux.scala 45:41]
  wire  _GEN_98 = _T_16 ? auto_stream_out_1_ready : _GEN_35; // @[Mux.scala 45:41]
  wire  _T_17 = _T_12 == 3'h4; // @[Mux.scala 45:28]
  wire  _GEN_102 = _T_17 ? auto_stream_in_4_bits_last : _GEN_93; // @[Mux.scala 45:41]
  wire [31:0] _GEN_105 = _T_17 ? auto_stream_in_4_bits_data : _GEN_96; // @[Mux.scala 45:41]
  wire  _GEN_106 = _T_17 ? auto_stream_in_4_valid : _GEN_97; // @[Mux.scala 45:41]
  wire  _GEN_107 = _T_17 ? auto_stream_out_1_ready : _GEN_44; // @[Mux.scala 45:41]
  wire  _T_18 = _T_12 == 3'h5; // @[Mux.scala 45:28]
  wire  _GEN_111 = _T_18 ? auto_stream_in_5_bits_last : _GEN_102; // @[Mux.scala 45:41]
  wire [31:0] _GEN_114 = _T_18 ? auto_stream_in_5_bits_data : _GEN_105; // @[Mux.scala 45:41]
  wire  _GEN_115 = _T_18 ? auto_stream_in_5_valid : _GEN_106; // @[Mux.scala 45:41]
  wire  _GEN_116 = _T_18 ? auto_stream_out_1_ready : _GEN_53; // @[Mux.scala 45:41]
  wire  _T_19 = _T_12 == 3'h6; // @[Mux.scala 45:28]
  wire  _GEN_125 = _T_19 ? auto_stream_out_1_ready : _GEN_62; // @[Mux.scala 45:41]
  wire  _T_20 = sels_0 == sels_2; // @[Mux.scala 40:46]
  wire  _T_21 = sels_1 == sels_2; // @[Mux.scala 40:46]
  wire  _T_23 = _T_20 | _T_21; // @[Mux.scala 40:75]
  wire [2:0] _T_24 = _T_23 ? 3'h7 : sels_2; // @[Mux.scala 41:29]
  wire  _T_25 = _T_24 == 3'h0; // @[Mux.scala 45:28]
  wire  _T_26 = _T_24 == 3'h1; // @[Mux.scala 45:28]
  wire  _T_27 = _T_24 == 3'h2; // @[Mux.scala 45:28]
  wire  _T_28 = _T_24 == 3'h3; // @[Mux.scala 45:28]
  wire  _T_29 = _T_24 == 3'h4; // @[Mux.scala 45:28]
  wire  _T_30 = _T_24 == 3'h5; // @[Mux.scala 45:28]
  wire  _T_31 = _T_24 == 3'h6; // @[Mux.scala 45:28]
  wire  _T_33 = auto_register_in_aw_valid & auto_register_in_w_valid; // @[RegisterRouter.scala 40:39]
  wire  _T_34 = auto_register_in_ar_valid | _T_33; // @[RegisterRouter.scala 40:26]
  wire  _T_35 = ~auto_register_in_ar_valid; // @[RegisterRouter.scala 42:29]
  wire  _T_78_ready = Queue_io_enq_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 299:17]
  wire [29:0] _T_42 = auto_register_in_ar_valid ? auto_register_in_ar_bits_addr : auto_register_in_aw_bits_addr; // @[RegisterRouter.scala 48:19]
  wire [1:0] _T_197 = {_T_42[3],_T_42[2]}; // @[Cat.scala 29:58]
  wire  _T_36 = _T_78_ready & _T_35; // @[RegisterRouter.scala 42:26]
  wire [1:0] _T_45 = 2'h1 << auto_register_in_ar_bits_size[0]; // @[OneHot.scala 65:12]
  wire [1:0] _T_47 = _T_45 | 2'h1; // @[Misc.scala 200:81]
  wire  _T_48 = auto_register_in_ar_bits_size >= 3'h2; // @[Misc.scala 204:21]
  wire  _T_51 = ~auto_register_in_ar_bits_addr[1]; // @[Misc.scala 209:20]
  wire  _T_53 = _T_47[1] & _T_51; // @[Misc.scala 213:38]
  wire  _T_54 = _T_48 | _T_53; // @[Misc.scala 213:29]
  wire  _T_56 = _T_47[1] & auto_register_in_ar_bits_addr[1]; // @[Misc.scala 213:38]
  wire  _T_57 = _T_48 | _T_56; // @[Misc.scala 213:29]
  wire  _T_60 = ~auto_register_in_ar_bits_addr[0]; // @[Misc.scala 209:20]
  wire  _T_61 = _T_51 & _T_60; // @[Misc.scala 212:27]
  wire  _T_62 = _T_47[0] & _T_61; // @[Misc.scala 213:38]
  wire  _T_63 = _T_54 | _T_62; // @[Misc.scala 213:29]
  wire  _T_64 = _T_51 & auto_register_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  wire  _T_65 = _T_47[0] & _T_64; // @[Misc.scala 213:38]
  wire  _T_66 = _T_54 | _T_65; // @[Misc.scala 213:29]
  wire  _T_67 = auto_register_in_ar_bits_addr[1] & _T_60; // @[Misc.scala 212:27]
  wire  _T_68 = _T_47[0] & _T_67; // @[Misc.scala 213:38]
  wire  _T_69 = _T_57 | _T_68; // @[Misc.scala 213:29]
  wire  _T_70 = auto_register_in_ar_bits_addr[1] & auto_register_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  wire  _T_71 = _T_47[0] & _T_70; // @[Misc.scala 213:38]
  wire  _T_72 = _T_57 | _T_71; // @[Misc.scala 213:29]
  wire [3:0] _T_75 = {_T_72,_T_69,_T_66,_T_63}; // @[Cat.scala 29:58]
  wire [3:0] _T_77 = auto_register_in_ar_valid ? _T_75 : auto_register_in_w_bits_strb; // @[RegisterRouter.scala 54:25]
  wire [7:0] _T_98 = _T_77[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_100 = _T_77[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_102 = _T_77[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_104 = _T_77[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_107 = {_T_104,_T_102,_T_100,_T_98}; // @[Cat.scala 29:58]
  wire  _T_126 = _T_107[2:0] == 3'h7; // @[RegisterRouter.scala 59:16]
  wire  _T_208 = _T_34 & _T_78_ready; // @[RegisterRouter.scala 59:16]
  wire [3:0] _T_198 = 4'h1 << _T_197; // @[OneHot.scala 58:35]
  wire  _T_235 = _T_208 & _T_35; // @[RegisterRouter.scala 59:16]
  wire  _T_247 = _T_235 & _T_198[2]; // @[RegisterRouter.scala 59:16]
  wire  _T_133 = _T_247 & _T_126; // @[RegisterRouter.scala 59:16]
  wire  _T_242 = _T_235 & _T_198[1]; // @[RegisterRouter.scala 59:16]
  wire  _T_156 = _T_242 & _T_126; // @[RegisterRouter.scala 59:16]
  wire  _T_237 = _T_235 & _T_198[0]; // @[RegisterRouter.scala 59:16]
  wire  _T_179 = _T_237 & _T_126; // @[RegisterRouter.scala 59:16]
  wire [2:0] _GEN_213 = 2'h1 == _T_197 ? sels_1 : sels_0; // @[MuxLiteral.scala 48:10]
  wire [2:0] _GEN_214 = 2'h2 == _T_197 ? sels_2 : _GEN_213; // @[MuxLiteral.scala 48:10]
  wire [2:0] _GEN_215 = 2'h3 == _T_197 ? 3'h0 : _GEN_214; // @[MuxLiteral.scala 48:10]
  wire  _T_323_bits_read = Queue_io_deq_bits_read; // @[Decoupled.scala 317:19 Decoupled.scala 318:14]
  wire  _T_323_valid = Queue_io_deq_valid; // @[Decoupled.scala 317:19 Decoupled.scala 319:15]
  wire  _T_326 = ~_T_323_bits_read; // @[RegisterRouter.scala 65:29]
  Queue Queue ( // @[Decoupled.scala 296:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_read(Queue_io_enq_bits_read),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_extra(Queue_io_enq_bits_extra),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_read(Queue_io_deq_bits_read),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_extra(Queue_io_deq_bits_extra)
  );
  assign auto_register_in_aw_ready = _T_36 & auto_register_in_w_valid; // @[LazyModule.scala 173:31]
  assign auto_register_in_w_ready = _T_36 & auto_register_in_aw_valid; // @[LazyModule.scala 173:31]
  assign auto_register_in_b_valid = _T_323_valid & _T_326; // @[LazyModule.scala 173:31]
  assign auto_register_in_b_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_register_in_ar_ready = Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_register_in_r_valid = _T_323_valid & _T_323_bits_read; // @[LazyModule.scala 173:31]
  assign auto_register_in_r_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_register_in_r_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 173:31]
  assign auto_stream_in_6_ready = _T_31 | _GEN_125; // @[LazyModule.scala 173:31]
  assign auto_stream_in_5_ready = _T_30 | _GEN_116; // @[LazyModule.scala 173:31]
  assign auto_stream_in_4_ready = _T_29 | _GEN_107; // @[LazyModule.scala 173:31]
  assign auto_stream_in_3_ready = _T_28 | _GEN_98; // @[LazyModule.scala 173:31]
  assign auto_stream_in_2_ready = _T_27 | _GEN_89; // @[LazyModule.scala 173:31]
  assign auto_stream_in_1_ready = _T_26 | _GEN_80; // @[LazyModule.scala 173:31]
  assign auto_stream_in_0_ready = _T_25 | _GEN_71; // @[LazyModule.scala 173:31]
  assign auto_stream_out_1_valid = _T_19 ? auto_stream_in_6_valid : _GEN_115; // @[LazyModule.scala 173:49]
  assign auto_stream_out_1_bits_data = _T_19 ? auto_stream_in_6_bits_data : _GEN_114; // @[LazyModule.scala 173:49]
  assign auto_stream_out_1_bits_last = _T_19 ? auto_stream_in_6_bits_last : _GEN_111; // @[LazyModule.scala 173:49]
  assign auto_stream_out_0_valid = _T_9 ? auto_stream_in_6_valid : _GEN_52; // @[LazyModule.scala 173:49]
  assign auto_stream_out_0_bits_data = _T_9 ? auto_stream_in_6_bits_data : _GEN_51; // @[LazyModule.scala 173:49]
  assign auto_stream_out_0_bits_last = _T_9 ? auto_stream_in_6_bits_last : _GEN_48; // @[LazyModule.scala 173:49]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_register_in_ar_valid | _T_33; // @[Decoupled.scala 297:22]
  assign Queue_io_enq_bits_read = auto_register_in_ar_valid; // @[Decoupled.scala 298:21]
  assign Queue_io_enq_bits_data = {{29'd0}, _GEN_215}; // @[Decoupled.scala 298:21]
  assign Queue_io_enq_bits_extra = auto_register_in_ar_valid ? auto_register_in_ar_bits_id : auto_register_in_aw_bits_id; // @[Decoupled.scala 298:21]
  assign Queue_io_deq_ready = _T_323_bits_read ? auto_register_in_r_ready : auto_register_in_b_ready; // @[Decoupled.scala 320:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  sels_0 = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  sels_1 = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  sels_2 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      sels_0 <= 3'h7;
    end else if (_T_179) begin
      sels_0 <= auto_register_in_w_bits_data[2:0];
    end
    if (reset) begin
      sels_1 <= 3'h7;
    end else if (_T_156) begin
      sels_1 <= auto_register_in_w_bits_data[2:0];
    end
    if (reset) begin
      sels_2 <= 3'h7;
    end else if (_T_133) begin
      sels_2 <= auto_register_in_w_bits_data[2:0];
    end
  end
endmodule
module Queue_37(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [31:0] io_enq_bits_data,
  input         io_enq_bits_last,
  input         io_deq_ready,
  output        io_deq_valid,
  output [31:0] io_deq_bits_data,
  output        io_deq_bits_last
);
  reg [31:0] _T_data [0:0]; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_0;
  wire [31:0] _T_data__T_14_data; // @[Decoupled.scala 218:24]
  wire  _T_data__T_14_addr; // @[Decoupled.scala 218:24]
  wire [31:0] _T_data__T_10_data; // @[Decoupled.scala 218:24]
  wire  _T_data__T_10_addr; // @[Decoupled.scala 218:24]
  wire  _T_data__T_10_mask; // @[Decoupled.scala 218:24]
  wire  _T_data__T_10_en; // @[Decoupled.scala 218:24]
  reg  _T_last [0:0]; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_1;
  wire  _T_last__T_14_data; // @[Decoupled.scala 218:24]
  wire  _T_last__T_14_addr; // @[Decoupled.scala 218:24]
  wire  _T_last__T_10_data; // @[Decoupled.scala 218:24]
  wire  _T_last__T_10_addr; // @[Decoupled.scala 218:24]
  wire  _T_last__T_10_mask; // @[Decoupled.scala 218:24]
  wire  _T_last__T_10_en; // @[Decoupled.scala 218:24]
  reg  _T_1; // @[Decoupled.scala 221:35]
  reg [31:0] _RAND_2;
  wire  _T_3 = ~_T_1; // @[Decoupled.scala 224:36]
  wire  _T_6 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  _T_8 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_13 = io_deq_ready ? 1'h0 : _T_6; // @[Decoupled.scala 249:27]
  wire  _GEN_22 = _T_3 ? _GEN_13 : _T_6; // @[Decoupled.scala 246:18]
  wire  _GEN_21 = _T_3 ? 1'h0 : _T_8; // @[Decoupled.scala 246:18]
  wire  _T_11 = _GEN_22 != _GEN_21; // @[Decoupled.scala 236:16]
  wire  _T_12 = ~_T_3; // @[Decoupled.scala 240:19]
  assign _T_data__T_14_addr = 1'h0;
  assign _T_data__T_14_data = _T_data[_T_data__T_14_addr]; // @[Decoupled.scala 218:24]
  assign _T_data__T_10_data = io_enq_bits_data;
  assign _T_data__T_10_addr = 1'h0;
  assign _T_data__T_10_mask = 1'h1;
  assign _T_data__T_10_en = _T_3 ? _GEN_13 : _T_6;
  assign _T_last__T_14_addr = 1'h0;
  assign _T_last__T_14_data = _T_last[_T_last__T_14_addr]; // @[Decoupled.scala 218:24]
  assign _T_last__T_10_data = io_enq_bits_last;
  assign _T_last__T_10_addr = 1'h0;
  assign _T_last__T_10_mask = 1'h1;
  assign _T_last__T_10_en = _T_3 ? _GEN_13 : _T_6;
  assign io_enq_ready = io_deq_ready | _T_3; // @[Decoupled.scala 241:16 Decoupled.scala 254:40]
  assign io_deq_valid = io_enq_valid | _T_12; // @[Decoupled.scala 240:16 Decoupled.scala 245:40]
  assign io_deq_bits_data = _T_3 ? io_enq_bits_data : _T_data__T_14_data; // @[Decoupled.scala 242:15 Decoupled.scala 247:19]
  assign io_deq_bits_last = _T_3 ? io_enq_bits_last : _T_last__T_14_data; // @[Decoupled.scala 242:15 Decoupled.scala 247:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_data[initvar] = _RAND_0[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_last[initvar] = _RAND_1[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_1 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T_data__T_10_en & _T_data__T_10_mask) begin
      _T_data[_T_data__T_10_addr] <= _T_data__T_10_data; // @[Decoupled.scala 218:24]
    end
    if(_T_last__T_10_en & _T_last__T_10_mask) begin
      _T_last[_T_last__T_10_addr] <= _T_last__T_10_data; // @[Decoupled.scala 218:24]
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else if (_T_11) begin
      if (_T_3) begin
        if (io_deq_ready) begin
          _T_1 <= 1'h0;
        end else begin
          _T_1 <= _T_6;
        end
      end else begin
        _T_1 <= _T_6;
      end
    end
  end
endmodule
module StreamBuffer_2(
  input         clock,
  input         reset,
  input         auto_out_out_ready,
  output        auto_out_out_valid,
  output [31:0] auto_out_out_bits_data,
  output        auto_out_out_bits_last,
  output        auto_in_in_ready,
  input         auto_in_in_valid,
  input  [31:0] auto_in_in_bits_data,
  input         auto_in_in_bits_last
);
  wire  Queue_clock; // @[Decoupled.scala 296:21]
  wire  Queue_reset; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [31:0] Queue_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_bits_last; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [31:0] Queue_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_bits_last; // @[Decoupled.scala 296:21]
  Queue_37 Queue ( // @[Decoupled.scala 296:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_last(Queue_io_enq_bits_last),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_last(Queue_io_deq_bits_last)
  );
  assign auto_out_out_valid = Queue_io_deq_valid; // @[LazyModule.scala 173:49]
  assign auto_out_out_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_out_bits_last = Queue_io_deq_bits_last; // @[LazyModule.scala 173:49]
  assign auto_in_in_ready = Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_in_in_valid; // @[Decoupled.scala 297:22]
  assign Queue_io_enq_bits_data = auto_in_in_bits_data; // @[Decoupled.scala 298:21]
  assign Queue_io_enq_bits_last = auto_in_in_bits_last; // @[Decoupled.scala 298:21]
  assign Queue_io_deq_ready = auto_out_out_ready; // @[Decoupled.scala 320:15]
endmodule
module AXI4StreamWidthAdapater_1_to_4(
  input         clock,
  input         reset,
  output        auto_in_ready,
  input         auto_in_valid,
  input  [31:0] auto_in_bits_data,
  input         auto_in_bits_last,
  input         auto_out_ready,
  output        auto_out_valid,
  output [7:0]  auto_out_bits_data,
  output        auto_out_bits_last
);
  reg [1:0] _T_5; // @[AXI4StreamWidthAdapter.scala 158:22]
  reg [31:0] _RAND_0;
  wire  _T_6 = auto_in_valid & auto_out_ready; // @[AXI4StreamWidthAdapter.scala 159:14]
  wire  _T_7 = _T_5 == 2'h3; // @[AXI4StreamWidthAdapter.scala 159:38]
  wire [2:0] _T_8 = _T_5 + 2'h1; // @[AXI4StreamWidthAdapter.scala 159:60]
  wire [2:0] _T_9 = _T_7 ? 3'h0 : _T_8; // @[AXI4StreamWidthAdapter.scala 159:33]
  wire [2:0] _GEN_0 = _T_6 ? _T_9 : {{1'd0}, _T_5}; // @[AXI4StreamWidthAdapter.scala 159:21]
  wire  ir0 = _T_7 & auto_out_ready; // @[AXI4StreamWidthAdapter.scala 163:34]
  reg [1:0] _T_11; // @[AXI4StreamWidthAdapter.scala 167:22]
  reg [31:0] _RAND_1;
  wire  _T_13 = _T_11 == 2'h3; // @[AXI4StreamWidthAdapter.scala 168:38]
  wire [2:0] _T_14 = _T_11 + 2'h1; // @[AXI4StreamWidthAdapter.scala 168:60]
  wire [2:0] _T_15 = _T_13 ? 3'h0 : _T_14; // @[AXI4StreamWidthAdapter.scala 168:33]
  wire [2:0] _GEN_1 = _T_6 ? _T_15 : {{1'd0}, _T_11}; // @[AXI4StreamWidthAdapter.scala 168:21]
  wire  ir1 = _T_13 & auto_out_ready; // @[AXI4StreamWidthAdapter.scala 170:60]
  reg [1:0] _T_20; // @[AXI4StreamWidthAdapter.scala 158:22]
  reg [31:0] _RAND_2;
  wire  _T_22 = _T_20 == 2'h3; // @[AXI4StreamWidthAdapter.scala 159:38]
  wire [2:0] _T_23 = _T_20 + 2'h1; // @[AXI4StreamWidthAdapter.scala 159:60]
  wire [2:0] _T_24 = _T_22 ? 3'h0 : _T_23; // @[AXI4StreamWidthAdapter.scala 159:33]
  wire [2:0] _GEN_2 = _T_6 ? _T_24 : {{1'd0}, _T_20}; // @[AXI4StreamWidthAdapter.scala 159:21]
  wire  ir2 = _T_22 & auto_out_ready; // @[AXI4StreamWidthAdapter.scala 163:34]
  reg [1:0] _T_27; // @[AXI4StreamWidthAdapter.scala 158:22]
  reg [31:0] _RAND_3;
  wire  _T_29 = _T_27 == 2'h3; // @[AXI4StreamWidthAdapter.scala 159:38]
  wire [2:0] _T_30 = _T_27 + 2'h1; // @[AXI4StreamWidthAdapter.scala 159:60]
  wire [2:0] _T_31 = _T_29 ? 3'h0 : _T_30; // @[AXI4StreamWidthAdapter.scala 159:33]
  wire [2:0] _GEN_3 = _T_6 ? _T_31 : {{1'd0}, _T_27}; // @[AXI4StreamWidthAdapter.scala 159:21]
  wire  ir3 = _T_29 & auto_out_ready; // @[AXI4StreamWidthAdapter.scala 163:34]
  reg [1:0] _T_34; // @[AXI4StreamWidthAdapter.scala 158:22]
  reg [31:0] _RAND_4;
  wire  _T_36 = _T_34 == 2'h3; // @[AXI4StreamWidthAdapter.scala 159:38]
  wire [2:0] _T_37 = _T_34 + 2'h1; // @[AXI4StreamWidthAdapter.scala 159:60]
  wire [2:0] _T_38 = _T_36 ? 3'h0 : _T_37; // @[AXI4StreamWidthAdapter.scala 159:33]
  wire [2:0] _GEN_4 = _T_6 ? _T_38 : {{1'd0}, _T_34}; // @[AXI4StreamWidthAdapter.scala 159:21]
  wire  ir4 = _T_36 & auto_out_ready; // @[AXI4StreamWidthAdapter.scala 163:34]
  wire  _T_56 = ir0 == ir1; // @[AXI4StreamWidthAdapter.scala 46:16]
  wire  _T_58 = _T_56 | reset; // @[AXI4StreamWidthAdapter.scala 46:11]
  wire  _T_59 = ~_T_58; // @[AXI4StreamWidthAdapter.scala 46:11]
  wire  _T_60 = ir0 == ir2; // @[AXI4StreamWidthAdapter.scala 47:16]
  wire  _T_62 = _T_60 | reset; // @[AXI4StreamWidthAdapter.scala 47:11]
  wire  _T_63 = ~_T_62; // @[AXI4StreamWidthAdapter.scala 47:11]
  wire  _T_64 = ir0 == ir3; // @[AXI4StreamWidthAdapter.scala 48:16]
  wire  _T_66 = _T_64 | reset; // @[AXI4StreamWidthAdapter.scala 48:11]
  wire  _T_67 = ~_T_66; // @[AXI4StreamWidthAdapter.scala 48:11]
  wire  _T_68 = ir0 == ir4; // @[AXI4StreamWidthAdapter.scala 49:16]
  wire  _T_70 = _T_68 | reset; // @[AXI4StreamWidthAdapter.scala 49:11]
  wire  _T_71 = ~_T_70; // @[AXI4StreamWidthAdapter.scala 49:11]
  wire [7:0] _GEN_6 = 2'h1 == _T_5 ? auto_in_bits_data[15:8] : auto_in_bits_data[7:0]; // @[AXI4StreamWidthAdapter.scala 54:19]
  wire [7:0] _GEN_7 = 2'h2 == _T_5 ? auto_in_bits_data[23:16] : _GEN_6; // @[AXI4StreamWidthAdapter.scala 54:19]
  assign auto_in_ready = _T_7 & auto_out_ready; // @[LazyModule.scala 173:31]
  assign auto_out_valid = auto_in_valid; // @[LazyModule.scala 173:49]
  assign auto_out_bits_data = 2'h3 == _T_5 ? auto_in_bits_data[31:24] : _GEN_7; // @[LazyModule.scala 173:49]
  assign auto_out_bits_last = auto_in_bits_last & _T_13; // @[LazyModule.scala 173:49]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_5 = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_11 = _RAND_1[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_20 = _RAND_2[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_27 = _RAND_3[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_34 = _RAND_4[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      _T_5 <= 2'h0;
    end else begin
      _T_5 <= _GEN_0[1:0];
    end
    if (reset) begin
      _T_11 <= 2'h0;
    end else begin
      _T_11 <= _GEN_1[1:0];
    end
    if (reset) begin
      _T_20 <= 2'h0;
    end else begin
      _T_20 <= _GEN_2[1:0];
    end
    if (reset) begin
      _T_27 <= 2'h0;
    end else begin
      _T_27 <= _GEN_3[1:0];
    end
    if (reset) begin
      _T_34 <= 2'h0;
    end else begin
      _T_34 <= _GEN_4[1:0];
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_59) begin
          $fwrite(32'h80000002,"Assertion failed\n    at AXI4StreamWidthAdapter.scala:46 assert(ir0 === ir1)\n"); // @[AXI4StreamWidthAdapter.scala 46:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_59) begin
          $fatal; // @[AXI4StreamWidthAdapter.scala 46:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_63) begin
          $fwrite(32'h80000002,"Assertion failed\n    at AXI4StreamWidthAdapter.scala:47 assert(ir0 === ir2)\n"); // @[AXI4StreamWidthAdapter.scala 47:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_63) begin
          $fatal; // @[AXI4StreamWidthAdapter.scala 47:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_67) begin
          $fwrite(32'h80000002,"Assertion failed\n    at AXI4StreamWidthAdapter.scala:48 assert(ir0 === ir3)\n"); // @[AXI4StreamWidthAdapter.scala 48:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_67) begin
          $fatal; // @[AXI4StreamWidthAdapter.scala 48:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_71) begin
          $fwrite(32'h80000002,"Assertion failed\n    at AXI4StreamWidthAdapter.scala:49 assert(ir0 === ir4)\n"); // @[AXI4StreamWidthAdapter.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_71) begin
          $fatal; // @[AXI4StreamWidthAdapter.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module Queue_38(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [31:0] io_enq_bits_data,
  input         io_enq_bits_last,
  input         io_deq_ready,
  output        io_deq_valid,
  output [31:0] io_deq_bits_data,
  output        io_deq_bits_last
);
  reg [31:0] _T_data [0:3]; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_0;
  wire [31:0] _T_data__T_18_data; // @[Decoupled.scala 218:24]
  wire [1:0] _T_data__T_18_addr; // @[Decoupled.scala 218:24]
  wire [31:0] _T_data__T_10_data; // @[Decoupled.scala 218:24]
  wire [1:0] _T_data__T_10_addr; // @[Decoupled.scala 218:24]
  wire  _T_data__T_10_mask; // @[Decoupled.scala 218:24]
  wire  _T_data__T_10_en; // @[Decoupled.scala 218:24]
  reg  _T_last [0:3]; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_1;
  wire  _T_last__T_18_data; // @[Decoupled.scala 218:24]
  wire [1:0] _T_last__T_18_addr; // @[Decoupled.scala 218:24]
  wire  _T_last__T_10_data; // @[Decoupled.scala 218:24]
  wire [1:0] _T_last__T_10_addr; // @[Decoupled.scala 218:24]
  wire  _T_last__T_10_mask; // @[Decoupled.scala 218:24]
  wire  _T_last__T_10_en; // @[Decoupled.scala 218:24]
  reg [1:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_2;
  reg [1:0] value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_3;
  reg  _T_1; // @[Decoupled.scala 221:35]
  reg [31:0] _RAND_4;
  wire  _T_2 = value == value_1; // @[Decoupled.scala 223:41]
  wire  _T_3 = ~_T_1; // @[Decoupled.scala 224:36]
  wire  _T_4 = _T_2 & _T_3; // @[Decoupled.scala 224:33]
  wire  _T_5 = _T_2 & _T_1; // @[Decoupled.scala 225:32]
  wire  _T_6 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  _T_8 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire [1:0] _T_12 = value + 2'h1; // @[Counter.scala 39:22]
  wire [1:0] _T_14 = value_1 + 2'h1; // @[Counter.scala 39:22]
  wire  _T_15 = _T_6 != _T_8; // @[Decoupled.scala 236:16]
  assign _T_data__T_18_addr = value_1;
  assign _T_data__T_18_data = _T_data[_T_data__T_18_addr]; // @[Decoupled.scala 218:24]
  assign _T_data__T_10_data = io_enq_bits_data;
  assign _T_data__T_10_addr = value;
  assign _T_data__T_10_mask = 1'h1;
  assign _T_data__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_last__T_18_addr = value_1;
  assign _T_last__T_18_data = _T_last[_T_last__T_18_addr]; // @[Decoupled.scala 218:24]
  assign _T_last__T_10_data = io_enq_bits_last;
  assign _T_last__T_10_addr = value;
  assign _T_last__T_10_mask = 1'h1;
  assign _T_last__T_10_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~_T_5; // @[Decoupled.scala 241:16]
  assign io_deq_valid = ~_T_4; // @[Decoupled.scala 240:16]
  assign io_deq_bits_data = _T_data__T_18_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_last = _T_last__T_18_data; // @[Decoupled.scala 242:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    _T_data[initvar] = _RAND_0[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    _T_last[initvar] = _RAND_1[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  value = _RAND_2[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  value_1 = _RAND_3[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T_data__T_10_en & _T_data__T_10_mask) begin
      _T_data[_T_data__T_10_addr] <= _T_data__T_10_data; // @[Decoupled.scala 218:24]
    end
    if(_T_last__T_10_en & _T_last__T_10_mask) begin
      _T_last[_T_last__T_10_addr] <= _T_last__T_10_data; // @[Decoupled.scala 218:24]
    end
    if (reset) begin
      value <= 2'h0;
    end else if (_T_6) begin
      value <= _T_12;
    end
    if (reset) begin
      value_1 <= 2'h0;
    end else if (_T_8) begin
      value_1 <= _T_14;
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else if (_T_15) begin
      _T_1 <= _T_6;
    end
  end
endmodule
module StreamBuffer_3(
  input         clock,
  input         reset,
  input         auto_out_out_ready,
  output        auto_out_out_valid,
  output [31:0] auto_out_out_bits_data,
  output        auto_out_out_bits_last,
  output        auto_in_in_ready,
  input         auto_in_in_valid,
  input  [31:0] auto_in_in_bits_data,
  input         auto_in_in_bits_last
);
  wire  Queue_clock; // @[Decoupled.scala 296:21]
  wire  Queue_reset; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [31:0] Queue_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_bits_last; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [31:0] Queue_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_bits_last; // @[Decoupled.scala 296:21]
  Queue_38 Queue ( // @[Decoupled.scala 296:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_last(Queue_io_enq_bits_last),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_last(Queue_io_deq_bits_last)
  );
  assign auto_out_out_valid = Queue_io_deq_valid; // @[LazyModule.scala 173:49]
  assign auto_out_out_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_out_bits_last = Queue_io_deq_bits_last; // @[LazyModule.scala 173:49]
  assign auto_in_in_ready = Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_in_in_valid; // @[Decoupled.scala 297:22]
  assign Queue_io_enq_bits_data = auto_in_in_bits_data; // @[Decoupled.scala 298:21]
  assign Queue_io_enq_bits_last = auto_in_in_bits_last; // @[Decoupled.scala 298:21]
  assign Queue_io_deq_ready = auto_out_out_ready; // @[Decoupled.scala 320:15]
endmodule
module IntToBundleBridge(
  input   auto_in_0,
  output  auto_out_0
);
  assign auto_out_0 = auto_in_0; // @[LazyModule.scala 173:49]
endmodule
module UARTTx(
  input         clock,
  input         reset,
  input         io_en,
  output        io_in_ready,
  input         io_in_valid,
  input  [7:0]  io_in_bits,
  output        io_out,
  input  [15:0] io_div,
  input         io_nstop
);
  wire [31:0] plusarg_reader_out; // @[PlusArg.scala 44:11]
  reg [15:0] prescaler; // @[UARTTx.scala 21:22]
  reg [31:0] _RAND_0;
  wire  pulse = prescaler == 16'h0; // @[UARTTx.scala 22:26]
  reg [3:0] counter; // @[UARTTx.scala 25:20]
  reg [31:0] _RAND_1;
  reg [8:0] shifter; // @[UARTTx.scala 26:20]
  reg [31:0] _RAND_2;
  reg  out; // @[UARTTx.scala 27:16]
  reg [31:0] _RAND_3;
  wire  plusarg_tx = plusarg_reader_out != 32'h0; // @[UARTTx.scala 30:90]
  wire  busy = counter != 4'h0; // @[UARTTx.scala 32:23]
  wire  _T = ~busy; // @[UARTTx.scala 33:27]
  wire  _T_2 = io_in_ready & io_in_valid; // @[Decoupled.scala 40:37]
  wire  _T_4 = ~reset; // @[UARTTx.scala 36:11]
  wire  _T_6 = _T_2 & plusarg_tx; // @[UARTTx.scala 38:22]
  wire [9:0] _T_9 = {1'h1,io_in_bits,1'h0}; // @[Cat.scala 29:58]
  wire  _T_10 = ~io_nstop; // @[UARTTx.scala 55:19]
  wire [3:0] _T_12 = _T_10 ? 4'ha : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_13 = io_nstop ? 4'hb : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_14 = _T_12 | _T_13; // @[Mux.scala 27:72]
  wire [3:0] _T_17 = _T_14 - 4'h0; // @[UARTTx.scala 55:53]
  wire [9:0] _GEN_0 = _T_6 ? _T_9 : {{1'd0}, shifter}; // @[UARTTx.scala 38:37]
  wire [15:0] _T_20 = prescaler - 16'h1; // @[UARTTx.scala 59:78]
  wire  _T_22 = pulse & busy; // @[UARTTx.scala 61:15]
  wire [3:0] _T_24 = counter - 4'h1; // @[UARTTx.scala 62:24]
  wire [8:0] _T_26 = {1'h1,shifter[8:1]}; // @[Cat.scala 29:58]
  wire [9:0] _GEN_4 = _T_22 ? {{1'd0}, _T_26} : _GEN_0; // @[UARTTx.scala 61:24]
  wire  _GEN_5 = _T_22 ? shifter[0] : out; // @[UARTTx.scala 61:24]
  plusarg_reader #(.FORMAT("uart_tx=%d"), .DEFAULT(1), .WIDTH(32)) plusarg_reader ( // @[PlusArg.scala 44:11]
    .out(plusarg_reader_out)
  );
  assign io_in_ready = io_en & _T; // @[UARTTx.scala 33:15]
  assign io_out = out; // @[UARTTx.scala 28:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  prescaler = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  counter = _RAND_1[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  shifter = _RAND_2[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      prescaler <= 16'h0;
    end else if (busy) begin
      if (pulse) begin
        prescaler <= io_div;
      end else begin
        prescaler <= _T_20;
      end
    end
    if (reset) begin
      counter <= 4'h0;
    end else if (_T_22) begin
      counter <= _T_24;
    end else if (_T_6) begin
      counter <= _T_17;
    end
    shifter <= _GEN_4[8:0];
    out <= reset | _GEN_5;
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & _T_4) begin
          $fwrite(32'h80000002,"UART TX (%x): %c\n",io_in_bits,io_in_bits); // @[UARTTx.scala 36:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module QueueCompatibility_6(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input  [7:0] io_enq_bits,
  input        io_deq_ready,
  output       io_deq_valid,
  output [7:0] io_deq_bits,
  output [4:0] io_count
);
  reg [7:0] _T [0:15]; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_0;
  wire [7:0] _T__T_18_data; // @[Decoupled.scala 218:24]
  wire [3:0] _T__T_18_addr; // @[Decoupled.scala 218:24]
  wire [7:0] _T__T_10_data; // @[Decoupled.scala 218:24]
  wire [3:0] _T__T_10_addr; // @[Decoupled.scala 218:24]
  wire  _T__T_10_mask; // @[Decoupled.scala 218:24]
  wire  _T__T_10_en; // @[Decoupled.scala 218:24]
  reg [3:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_1;
  reg [3:0] value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_2;
  reg  _T_1; // @[Decoupled.scala 221:35]
  reg [31:0] _RAND_3;
  wire  _T_2 = value == value_1; // @[Decoupled.scala 223:41]
  wire  _T_3 = ~_T_1; // @[Decoupled.scala 224:36]
  wire  _T_4 = _T_2 & _T_3; // @[Decoupled.scala 224:33]
  wire  _T_5 = _T_2 & _T_1; // @[Decoupled.scala 225:32]
  wire  _T_6 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  _T_8 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire [3:0] _T_12 = value + 4'h1; // @[Counter.scala 39:22]
  wire [3:0] _T_14 = value_1 + 4'h1; // @[Counter.scala 39:22]
  wire  _T_15 = _T_6 != _T_8; // @[Decoupled.scala 236:16]
  wire [3:0] _T_20 = value - value_1; // @[Decoupled.scala 257:40]
  wire  _T_21 = _T_1 & _T_2; // @[Decoupled.scala 259:32]
  wire [4:0] _T_22 = _T_21 ? 5'h10 : 5'h0; // @[Decoupled.scala 259:20]
  wire [4:0] _GEN_8 = {{1'd0}, _T_20}; // @[Decoupled.scala 259:62]
  assign _T__T_18_addr = value_1;
  assign _T__T_18_data = _T[_T__T_18_addr]; // @[Decoupled.scala 218:24]
  assign _T__T_10_data = io_enq_bits;
  assign _T__T_10_addr = value;
  assign _T__T_10_mask = 1'h1;
  assign _T__T_10_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~_T_5; // @[Decoupled.scala 241:16]
  assign io_deq_valid = ~_T_4; // @[Decoupled.scala 240:16]
  assign io_deq_bits = _T__T_18_data; // @[Decoupled.scala 242:15]
  assign io_count = _T_22 | _GEN_8; // @[Decoupled.scala 259:14]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    _T[initvar] = _RAND_0[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  value = _RAND_1[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  value_1 = _RAND_2[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_1 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T__T_10_en & _T__T_10_mask) begin
      _T[_T__T_10_addr] <= _T__T_10_data; // @[Decoupled.scala 218:24]
    end
    if (reset) begin
      value <= 4'h0;
    end else if (_T_6) begin
      value <= _T_12;
    end
    if (reset) begin
      value_1 <= 4'h0;
    end else if (_T_8) begin
      value_1 <= _T_14;
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else if (_T_15) begin
      _T_1 <= _T_6;
    end
  end
endmodule
module UARTRx(
  input         clock,
  input         reset,
  input         io_en,
  input         io_in,
  output        io_out_valid,
  output [7:0]  io_out_bits,
  input  [15:0] io_div
);
  reg [1:0] debounce; // @[UARTRx.scala 22:21]
  reg [31:0] _RAND_0;
  wire  debounce_max = debounce == 2'h3; // @[UARTRx.scala 23:32]
  wire  debounce_min = debounce == 2'h0; // @[UARTRx.scala 24:32]
  reg [12:0] prescaler; // @[UARTRx.scala 26:22]
  reg [31:0] _RAND_1;
  wire  pulse = prescaler == 13'h0; // @[UARTRx.scala 28:26]
  reg [3:0] data_count; // @[UARTRx.scala 32:23]
  reg [31:0] _RAND_2;
  wire  data_last = data_count == 4'h0; // @[UARTRx.scala 33:31]
  reg [3:0] sample_count; // @[UARTRx.scala 35:25]
  reg [31:0] _RAND_3;
  wire  sample_mid = sample_count == 4'h7; // @[UARTRx.scala 36:34]
  wire [7:0] _T_1 = {data_count,sample_count}; // @[Cat.scala 29:58]
  wire [7:0] countdown = _T_1 - 8'h1; // @[UARTRx.scala 38:49]
  wire [3:0] remainder = io_div[3:0]; // @[UARTRx.scala 43:25]
  wire  extend = sample_count < remainder; // @[UARTRx.scala 44:30]
  reg  state; // @[UARTRx.scala 59:18]
  reg [31:0] _RAND_4;
  wire  _T_14 = ~state; // @[Conditional.scala 37:30]
  wire  _T_21 = ~io_in; // @[UARTRx.scala 66:13]
  wire  _GEN_8 = _T_21 & debounce_max; // @[UARTRx.scala 66:21]
  wire  start = _T_14 & _GEN_8; // @[Conditional.scala 40:58]
  wire  restore = start | pulse; // @[UARTRx.scala 45:23]
  wire [12:0] prescaler_in = restore ? {{1'd0}, io_div[15:4]} : prescaler; // @[UARTRx.scala 46:25]
  wire  _T_4 = restore & extend; // @[UARTRx.scala 47:51]
  wire  _T_5 = _T_4 ? 1'h0 : 1'h1; // @[UARTRx.scala 47:42]
  wire [12:0] _GEN_41 = {{12'd0}, _T_5}; // @[UARTRx.scala 47:37]
  wire [12:0] prescaler_next = prescaler_in - _GEN_41; // @[UARTRx.scala 47:37]
  reg [2:0] sample; // @[UARTRx.scala 49:19]
  reg [31:0] _RAND_5;
  wire  _T_10 = sample[0] & sample[1]; // @[Misc.scala 165:48]
  wire  _T_11 = sample[0] & sample[2]; // @[Misc.scala 165:48]
  wire  _T_12 = _T_10 | _T_11; // @[Misc.scala 166:22]
  wire  _T_13 = sample[1] & sample[2]; // @[Misc.scala 165:48]
  wire  voter = _T_12 | _T_13; // @[Misc.scala 166:22]
  reg [7:0] shifter; // @[UARTRx.scala 51:20]
  reg [31:0] _RAND_6;
  reg  valid; // @[UARTRx.scala 53:18]
  reg [31:0] _RAND_7;
  wire  _T_16 = ~_T_21; // @[UARTRx.scala 63:13]
  wire  _T_17 = ~debounce_min; // @[UARTRx.scala 63:26]
  wire  _T_18 = _T_16 & _T_17; // @[UARTRx.scala 63:23]
  wire [1:0] _T_20 = debounce - 2'h1; // @[UARTRx.scala 64:30]
  wire [1:0] _T_23 = debounce + 2'h1; // @[UARTRx.scala 67:30]
  wire [3:0] _T_27 = 4'h9 - 4'h0; // @[UARTRx.scala 72:94]
  wire  _GEN_1 = debounce_max | state; // @[UARTRx.scala 68:29]
  wire [3:0] _T_29 = {sample,io_in}; // @[Cat.scala 29:58]
  wire [7:0] _T_33 = {voter,shifter[7:1]}; // @[Cat.scala 29:58]
  wire  _GEN_16 = sample_mid & data_last; // @[UARTRx.scala 85:27]
  wire [3:0] _GEN_18 = pulse ? _T_29 : {{1'd0}, sample}; // @[UARTRx.scala 80:20]
  wire  _GEN_22 = pulse & _GEN_16; // @[UARTRx.scala 80:20]
  wire [3:0] _GEN_25 = state ? _GEN_18 : {{1'd0}, sample}; // @[Conditional.scala 39:67]
  wire  _GEN_29 = state & _GEN_22; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_37 = _T_14 ? {{1'd0}, sample} : _GEN_25; // @[Conditional.scala 40:58]
  wire  _T_34 = ~io_en; // @[UARTRx.scala 112:9]
  assign io_out_valid = valid; // @[UARTRx.scala 55:16]
  assign io_out_bits = shifter; // @[UARTRx.scala 56:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  debounce = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  prescaler = _RAND_1[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  data_count = _RAND_2[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  sample_count = _RAND_3[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  state = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  sample = _RAND_5[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  shifter = _RAND_6[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  valid = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      debounce <= 2'h0;
    end else if (_T_34) begin
      debounce <= 2'h0;
    end else if (_T_14) begin
      if (_T_21) begin
        debounce <= _T_23;
      end else if (_T_18) begin
        debounce <= _T_20;
      end
    end
    if (_T_14) begin
      if (_T_21) begin
        if (debounce_max) begin
          prescaler <= prescaler_next;
        end
      end
    end else if (state) begin
      prescaler <= prescaler_next;
    end
    if (_T_14) begin
      if (_T_21) begin
        if (debounce_max) begin
          data_count <= _T_27;
        end
      end
    end else if (state) begin
      if (pulse) begin
        data_count <= countdown[7:4];
      end
    end
    if (_T_14) begin
      if (_T_21) begin
        if (debounce_max) begin
          sample_count <= 4'hf;
        end
      end
    end else if (state) begin
      if (pulse) begin
        sample_count <= countdown[3:0];
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else if (_T_14) begin
      if (_T_21) begin
        state <= _GEN_1;
      end
    end else if (state) begin
      if (pulse) begin
        if (sample_mid) begin
          if (data_last) begin
            state <= 1'h0;
          end
        end
      end
    end
    sample <= _GEN_37[2:0];
    if (!(_T_14)) begin
      if (state) begin
        if (pulse) begin
          if (sample_mid) begin
            if (!(data_last)) begin
              shifter <= _T_33;
            end
          end
        end
      end
    end
    if (reset) begin
      valid <= 1'h0;
    end else if (_T_14) begin
      valid <= 1'h0;
    end else begin
      valid <= _GEN_29;
    end
  end
endmodule
module AXI4UARTBlock(
  input         clock,
  input         reset,
  output        auto_mem_in_aw_ready,
  input         auto_mem_in_aw_valid,
  input         auto_mem_in_aw_bits_id,
  input  [29:0] auto_mem_in_aw_bits_addr,
  output        auto_mem_in_w_ready,
  input         auto_mem_in_w_valid,
  input  [31:0] auto_mem_in_w_bits_data,
  input  [3:0]  auto_mem_in_w_bits_strb,
  input         auto_mem_in_b_ready,
  output        auto_mem_in_b_valid,
  output        auto_mem_in_b_bits_id,
  output        auto_mem_in_ar_ready,
  input         auto_mem_in_ar_valid,
  input         auto_mem_in_ar_bits_id,
  input  [29:0] auto_mem_in_ar_bits_addr,
  input  [2:0]  auto_mem_in_ar_bits_size,
  input         auto_mem_in_r_ready,
  output        auto_mem_in_r_valid,
  output        auto_mem_in_r_bits_id,
  output [31:0] auto_mem_in_r_bits_data,
  output        auto_in_in_ready,
  input         auto_in_in_valid,
  input  [7:0]  auto_in_in_bits_data,
  input         auto_out_out_ready,
  output        auto_out_out_valid,
  output [7:0]  auto_out_out_bits_data,
  output        int_0,
  output        io_txd,
  input         io_rxd
);
  wire  converter_auto_in_0; // @[Nodes.scala 31:31]
  wire  converter_auto_out_0; // @[Nodes.scala 31:31]
  wire  txm_clock; // @[DSPBlockUART.scala 101:21]
  wire  txm_reset; // @[DSPBlockUART.scala 101:21]
  wire  txm_io_en; // @[DSPBlockUART.scala 101:21]
  wire  txm_io_in_ready; // @[DSPBlockUART.scala 101:21]
  wire  txm_io_in_valid; // @[DSPBlockUART.scala 101:21]
  wire [7:0] txm_io_in_bits; // @[DSPBlockUART.scala 101:21]
  wire  txm_io_out; // @[DSPBlockUART.scala 101:21]
  wire [15:0] txm_io_div; // @[DSPBlockUART.scala 101:21]
  wire  txm_io_nstop; // @[DSPBlockUART.scala 101:21]
  wire  txq_clock; // @[DSPBlockUART.scala 102:21]
  wire  txq_reset; // @[DSPBlockUART.scala 102:21]
  wire  txq_io_enq_ready; // @[DSPBlockUART.scala 102:21]
  wire  txq_io_enq_valid; // @[DSPBlockUART.scala 102:21]
  wire [7:0] txq_io_enq_bits; // @[DSPBlockUART.scala 102:21]
  wire  txq_io_deq_ready; // @[DSPBlockUART.scala 102:21]
  wire  txq_io_deq_valid; // @[DSPBlockUART.scala 102:21]
  wire [7:0] txq_io_deq_bits; // @[DSPBlockUART.scala 102:21]
  wire [4:0] txq_io_count; // @[DSPBlockUART.scala 102:21]
  wire  rxm_clock; // @[DSPBlockUART.scala 104:21]
  wire  rxm_reset; // @[DSPBlockUART.scala 104:21]
  wire  rxm_io_en; // @[DSPBlockUART.scala 104:21]
  wire  rxm_io_in; // @[DSPBlockUART.scala 104:21]
  wire  rxm_io_out_valid; // @[DSPBlockUART.scala 104:21]
  wire [7:0] rxm_io_out_bits; // @[DSPBlockUART.scala 104:21]
  wire [15:0] rxm_io_div; // @[DSPBlockUART.scala 104:21]
  wire  rxq_clock; // @[DSPBlockUART.scala 105:21]
  wire  rxq_reset; // @[DSPBlockUART.scala 105:21]
  wire  rxq_io_enq_ready; // @[DSPBlockUART.scala 105:21]
  wire  rxq_io_enq_valid; // @[DSPBlockUART.scala 105:21]
  wire [7:0] rxq_io_enq_bits; // @[DSPBlockUART.scala 105:21]
  wire  rxq_io_deq_ready; // @[DSPBlockUART.scala 105:21]
  wire  rxq_io_deq_valid; // @[DSPBlockUART.scala 105:21]
  wire [7:0] rxq_io_deq_bits; // @[DSPBlockUART.scala 105:21]
  wire [4:0] rxq_io_count; // @[DSPBlockUART.scala 105:21]
  wire  Queue_clock; // @[Decoupled.scala 296:21]
  wire  Queue_reset; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_bits_read; // @[Decoupled.scala 296:21]
  wire [31:0] Queue_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_bits_extra; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_bits_read; // @[Decoupled.scala 296:21]
  wire [31:0] Queue_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_bits_extra; // @[Decoupled.scala 296:21]
  reg [15:0] div; // @[DSPBlockUART.scala 107:18]
  reg [31:0] _RAND_0;
  reg  txen; // @[DSPBlockUART.scala 113:19]
  reg [31:0] _RAND_1;
  reg  rxen; // @[DSPBlockUART.scala 114:19]
  reg [31:0] _RAND_2;
  reg [4:0] txwm; // @[DSPBlockUART.scala 121:19]
  reg [31:0] _RAND_3;
  reg [4:0] rxwm; // @[DSPBlockUART.scala 122:19]
  reg [31:0] _RAND_4;
  reg  nstop; // @[DSPBlockUART.scala 123:20]
  reg [31:0] _RAND_5;
  reg  ie_rxwm; // @[DSPBlockUART.scala 166:17]
  reg [31:0] _RAND_6;
  reg  ie_txwm; // @[DSPBlockUART.scala 166:17]
  reg [31:0] _RAND_7;
  wire  ip_txwm = txq_io_count < txwm; // @[DSPBlockUART.scala 169:30]
  wire  ip_rxwm = rxq_io_count > rxwm; // @[DSPBlockUART.scala 170:30]
  wire  _T_8 = ip_txwm & ie_txwm; // @[DSPBlockUART.scala 171:31]
  wire  _T_9 = ip_rxwm & ie_rxwm; // @[DSPBlockUART.scala 171:55]
  reg [31:0] _T_11; // @[DSPBlockUART.scala 175:53]
  reg [31:0] _RAND_8;
  reg [31:0] _T_12; // @[DSPBlockUART.scala 177:53]
  reg [31:0] _RAND_9;
  wire  _T_14 = auto_mem_in_aw_valid & auto_mem_in_w_valid; // @[RegisterRouter.scala 40:39]
  wire  _T_15 = auto_mem_in_ar_valid | _T_14; // @[RegisterRouter.scala 40:26]
  wire  _T_16 = ~auto_mem_in_ar_valid; // @[RegisterRouter.scala 42:29]
  wire  _T_59_ready = Queue_io_enq_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 299:17]
  wire [29:0] _T_23 = auto_mem_in_ar_valid ? auto_mem_in_ar_bits_addr : auto_mem_in_aw_bits_addr; // @[RegisterRouter.scala 48:19]
  wire [2:0] _T_413 = {_T_23[4],_T_23[3],_T_23[2]}; // @[Cat.scala 29:58]
  wire [5:0] _T_63 = _T_23[7:2] & 6'h38; // @[RegisterRouter.scala 59:16]
  wire  _T_71 = _T_63 == 6'h0; // @[RegisterRouter.scala 59:16]
  wire  _T_17 = _T_59_ready & _T_16; // @[RegisterRouter.scala 42:26]
  wire [1:0] _T_26 = 2'h1 << auto_mem_in_ar_bits_size[0]; // @[OneHot.scala 65:12]
  wire [1:0] _T_28 = _T_26 | 2'h1; // @[Misc.scala 200:81]
  wire  _T_29 = auto_mem_in_ar_bits_size >= 3'h2; // @[Misc.scala 204:21]
  wire  _T_32 = ~auto_mem_in_ar_bits_addr[1]; // @[Misc.scala 209:20]
  wire  _T_34 = _T_28[1] & _T_32; // @[Misc.scala 213:38]
  wire  _T_35 = _T_29 | _T_34; // @[Misc.scala 213:29]
  wire  _T_37 = _T_28[1] & auto_mem_in_ar_bits_addr[1]; // @[Misc.scala 213:38]
  wire  _T_38 = _T_29 | _T_37; // @[Misc.scala 213:29]
  wire  _T_41 = ~auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 209:20]
  wire  _T_42 = _T_32 & _T_41; // @[Misc.scala 212:27]
  wire  _T_43 = _T_28[0] & _T_42; // @[Misc.scala 213:38]
  wire  _T_44 = _T_35 | _T_43; // @[Misc.scala 213:29]
  wire  _T_45 = _T_32 & auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  wire  _T_46 = _T_28[0] & _T_45; // @[Misc.scala 213:38]
  wire  _T_47 = _T_35 | _T_46; // @[Misc.scala 213:29]
  wire  _T_48 = auto_mem_in_ar_bits_addr[1] & _T_41; // @[Misc.scala 212:27]
  wire  _T_49 = _T_28[0] & _T_48; // @[Misc.scala 213:38]
  wire  _T_50 = _T_38 | _T_49; // @[Misc.scala 213:29]
  wire  _T_51 = auto_mem_in_ar_bits_addr[1] & auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  wire  _T_52 = _T_28[0] & _T_51; // @[Misc.scala 213:38]
  wire  _T_53 = _T_38 | _T_52; // @[Misc.scala 213:29]
  wire [3:0] _T_56 = {_T_53,_T_50,_T_47,_T_44}; // @[Cat.scala 29:58]
  wire [3:0] _T_58 = auto_mem_in_ar_valid ? _T_56 : auto_mem_in_w_bits_strb; // @[RegisterRouter.scala 54:25]
  wire [7:0] _T_87 = _T_58[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_89 = _T_58[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_91 = _T_58[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_93 = _T_58[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_96 = {_T_93,_T_91,_T_89,_T_87}; // @[Cat.scala 29:58]
  wire  _T_115 = _T_96 == 32'hffffffff; // @[RegisterRouter.scala 59:16]
  wire  _T_432 = _T_15 & _T_59_ready; // @[RegisterRouter.scala 59:16]
  wire [7:0] _T_414 = 8'h1 << _T_413; // @[OneHot.scala 58:35]
  wire  _T_479 = _T_432 & _T_16; // @[RegisterRouter.scala 59:16]
  wire  _T_481 = _T_479 & _T_414[0]; // @[RegisterRouter.scala 59:16]
  wire  _T_482 = _T_481 & _T_71; // @[RegisterRouter.scala 59:16]
  wire  _T_122 = _T_482 & _T_115; // @[RegisterRouter.scala 59:16]
  wire [1:0] _T_180 = {ip_rxwm,ip_txwm}; // @[Cat.scala 29:58]
  wire  _T_486 = _T_479 & _T_414[1]; // @[RegisterRouter.scala 59:16]
  wire  _T_487 = _T_486 & _T_71; // @[RegisterRouter.scala 59:16]
  wire  _T_193 = _T_487 & _T_115; // @[RegisterRouter.scala 59:16]
  wire  _T_209 = _T_96[15:0] == 16'hffff; // @[RegisterRouter.scala 59:16]
  wire  _T_511 = _T_479 & _T_414[6]; // @[RegisterRouter.scala 59:16]
  wire  _T_512 = _T_511 & _T_71; // @[RegisterRouter.scala 59:16]
  wire  _T_216 = _T_512 & _T_209; // @[RegisterRouter.scala 59:16]
  wire  _T_491 = _T_479 & _T_414[2]; // @[RegisterRouter.scala 59:16]
  wire  _T_492 = _T_491 & _T_71; // @[RegisterRouter.scala 59:16]
  wire  _T_239 = _T_492 & _T_96[0]; // @[RegisterRouter.scala 59:16]
  wire  _T_262 = _T_492 & _T_96[1]; // @[RegisterRouter.scala 59:16]
  wire [1:0] _T_274 = {nstop,txen}; // @[Cat.scala 29:58]
  wire  _T_280 = _T_96[20:16] == 5'h1f; // @[RegisterRouter.scala 59:16]
  wire  _T_287 = _T_492 & _T_280; // @[RegisterRouter.scala 59:16]
  wire [15:0] _T_298 = {{14'd0}, _T_274}; // @[RegisterRouter.scala 59:16]
  wire [20:0] _T_299 = {txwm,_T_298}; // @[Cat.scala 29:58]
  wire  _T_496 = _T_479 & _T_414[3]; // @[RegisterRouter.scala 59:16]
  wire  _T_497 = _T_496 & _T_71; // @[RegisterRouter.scala 59:16]
  wire  _T_312 = _T_497 & _T_96[0]; // @[RegisterRouter.scala 59:16]
  wire  _T_335 = _T_497 & _T_280; // @[RegisterRouter.scala 59:16]
  wire [15:0] _T_346 = {{15'd0}, rxen}; // @[RegisterRouter.scala 59:16]
  wire [20:0] _T_347 = {rxwm,_T_346}; // @[Cat.scala 29:58]
  wire  _T_501 = _T_479 & _T_414[4]; // @[RegisterRouter.scala 59:16]
  wire  _T_502 = _T_501 & _T_71; // @[RegisterRouter.scala 59:16]
  wire  _T_360 = _T_502 & _T_96[0]; // @[RegisterRouter.scala 59:16]
  wire  _T_383 = _T_502 & _T_96[1]; // @[RegisterRouter.scala 59:16]
  wire [1:0] _T_395 = {ie_rxwm,ie_txwm}; // @[Cat.scala 29:58]
  wire  _GEN_43 = 3'h1 == _T_413 ? _T_71 : _T_71; // @[MuxLiteral.scala 48:10]
  wire  _GEN_44 = 3'h2 == _T_413 ? _T_71 : _GEN_43; // @[MuxLiteral.scala 48:10]
  wire  _GEN_45 = 3'h3 == _T_413 ? _T_71 : _GEN_44; // @[MuxLiteral.scala 48:10]
  wire  _GEN_46 = 3'h4 == _T_413 ? _T_71 : _GEN_45; // @[MuxLiteral.scala 48:10]
  wire  _GEN_47 = 3'h5 == _T_413 ? _T_71 : _GEN_46; // @[MuxLiteral.scala 48:10]
  wire  _GEN_48 = 3'h6 == _T_413 ? _T_71 : _GEN_47; // @[MuxLiteral.scala 48:10]
  wire  _GEN_58 = 3'h7 == _T_413; // @[MuxLiteral.scala 48:10]
  wire  _GEN_49 = _GEN_58 | _GEN_48; // @[MuxLiteral.scala 48:10]
  wire [31:0] _GEN_51 = 3'h1 == _T_413 ? _T_12 : _T_11; // @[MuxLiteral.scala 48:10]
  wire [31:0] _T_624_2 = {{11'd0}, _T_299}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [31:0] _GEN_52 = 3'h2 == _T_413 ? _T_624_2 : _GEN_51; // @[MuxLiteral.scala 48:10]
  wire [31:0] _T_624_3 = {{11'd0}, _T_347}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [31:0] _GEN_53 = 3'h3 == _T_413 ? _T_624_3 : _GEN_52; // @[MuxLiteral.scala 48:10]
  wire [31:0] _T_624_4 = {{30'd0}, _T_395}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [31:0] _GEN_54 = 3'h4 == _T_413 ? _T_624_4 : _GEN_53; // @[MuxLiteral.scala 48:10]
  wire [31:0] _T_624_5 = {{30'd0}, _T_180}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [31:0] _GEN_55 = 3'h5 == _T_413 ? _T_624_5 : _GEN_54; // @[MuxLiteral.scala 48:10]
  wire [31:0] _T_624_6 = {{16'd0}, div}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [31:0] _GEN_56 = 3'h6 == _T_413 ? _T_624_6 : _GEN_55; // @[MuxLiteral.scala 48:10]
  wire [31:0] _GEN_57 = 3'h7 == _T_413 ? 32'h0 : _GEN_56; // @[MuxLiteral.scala 48:10]
  wire  _T_627_bits_read = Queue_io_deq_bits_read; // @[Decoupled.scala 317:19 Decoupled.scala 318:14]
  wire  _T_627_valid = Queue_io_deq_valid; // @[Decoupled.scala 317:19 Decoupled.scala 319:15]
  wire  _T_630 = ~_T_627_bits_read; // @[RegisterRouter.scala 65:29]
  IntToBundleBridge converter ( // @[Nodes.scala 31:31]
    .auto_in_0(converter_auto_in_0),
    .auto_out_0(converter_auto_out_0)
  );
  UARTTx txm ( // @[DSPBlockUART.scala 101:21]
    .clock(txm_clock),
    .reset(txm_reset),
    .io_en(txm_io_en),
    .io_in_ready(txm_io_in_ready),
    .io_in_valid(txm_io_in_valid),
    .io_in_bits(txm_io_in_bits),
    .io_out(txm_io_out),
    .io_div(txm_io_div),
    .io_nstop(txm_io_nstop)
  );
  QueueCompatibility_6 txq ( // @[DSPBlockUART.scala 102:21]
    .clock(txq_clock),
    .reset(txq_reset),
    .io_enq_ready(txq_io_enq_ready),
    .io_enq_valid(txq_io_enq_valid),
    .io_enq_bits(txq_io_enq_bits),
    .io_deq_ready(txq_io_deq_ready),
    .io_deq_valid(txq_io_deq_valid),
    .io_deq_bits(txq_io_deq_bits),
    .io_count(txq_io_count)
  );
  UARTRx rxm ( // @[DSPBlockUART.scala 104:21]
    .clock(rxm_clock),
    .reset(rxm_reset),
    .io_en(rxm_io_en),
    .io_in(rxm_io_in),
    .io_out_valid(rxm_io_out_valid),
    .io_out_bits(rxm_io_out_bits),
    .io_div(rxm_io_div)
  );
  QueueCompatibility_6 rxq ( // @[DSPBlockUART.scala 105:21]
    .clock(rxq_clock),
    .reset(rxq_reset),
    .io_enq_ready(rxq_io_enq_ready),
    .io_enq_valid(rxq_io_enq_valid),
    .io_enq_bits(rxq_io_enq_bits),
    .io_deq_ready(rxq_io_deq_ready),
    .io_deq_valid(rxq_io_deq_valid),
    .io_deq_bits(rxq_io_deq_bits),
    .io_count(rxq_io_count)
  );
  Queue Queue ( // @[Decoupled.scala 296:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_read(Queue_io_enq_bits_read),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_extra(Queue_io_enq_bits_extra),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_read(Queue_io_deq_bits_read),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_extra(Queue_io_deq_bits_extra)
  );
  assign auto_mem_in_aw_ready = _T_17 & auto_mem_in_w_valid; // @[LazyModule.scala 173:31]
  assign auto_mem_in_w_ready = _T_17 & auto_mem_in_aw_valid; // @[LazyModule.scala 173:31]
  assign auto_mem_in_b_valid = _T_627_valid & _T_630; // @[LazyModule.scala 173:31]
  assign auto_mem_in_b_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_mem_in_ar_ready = Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_valid = _T_627_valid & _T_627_bits_read; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 173:31]
  assign auto_in_in_ready = txq_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_out_out_valid = rxq_io_deq_valid; // @[LazyModule.scala 173:49]
  assign auto_out_out_bits_data = rxq_io_deq_bits; // @[LazyModule.scala 173:49]
  assign int_0 = converter_auto_out_0; // @[SpectrometerTest.scala 173:12]
  assign io_txd = txm_io_out; // @[DSPBlockUART.scala 135:12]
  assign converter_auto_in_0 = _T_8 | _T_9; // @[LazyModule.scala 167:57]
  assign txm_clock = clock;
  assign txm_reset = reset;
  assign txm_io_en = txen; // @[DSPBlockUART.scala 131:19]
  assign txm_io_in_valid = txq_io_deq_valid; // @[DSPBlockUART.scala 132:15]
  assign txm_io_in_bits = txq_io_deq_bits; // @[DSPBlockUART.scala 132:15]
  assign txm_io_div = div; // @[DSPBlockUART.scala 133:16]
  assign txm_io_nstop = nstop; // @[DSPBlockUART.scala 134:18]
  assign txq_clock = clock;
  assign txq_reset = reset;
  assign txq_io_enq_valid = auto_in_in_valid; // @[DSPBlockUART.scala 139:22]
  assign txq_io_enq_bits = auto_in_in_bits_data; // @[DSPBlockUART.scala 138:22]
  assign txq_io_deq_ready = txm_io_in_ready; // @[DSPBlockUART.scala 132:15]
  assign rxm_clock = clock;
  assign rxm_reset = reset;
  assign rxm_io_en = rxen; // @[DSPBlockUART.scala 151:15]
  assign rxm_io_in = io_rxd; // @[DSPBlockUART.scala 152:15]
  assign rxm_io_div = div; // @[DSPBlockUART.scala 154:16]
  assign rxq_clock = clock;
  assign rxq_reset = reset;
  assign rxq_io_enq_valid = rxm_io_out_valid; // @[DSPBlockUART.scala 153:16]
  assign rxq_io_enq_bits = rxm_io_out_bits; // @[DSPBlockUART.scala 153:16]
  assign rxq_io_deq_ready = auto_out_out_ready; // @[DSPBlockUART.scala 144:22]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_mem_in_ar_valid | _T_14; // @[Decoupled.scala 297:22]
  assign Queue_io_enq_bits_read = auto_mem_in_ar_valid; // @[Decoupled.scala 298:21]
  assign Queue_io_enq_bits_data = _GEN_49 ? _GEN_57 : 32'h0; // @[Decoupled.scala 298:21]
  assign Queue_io_enq_bits_extra = auto_mem_in_ar_valid ? auto_mem_in_ar_bits_id : auto_mem_in_aw_bits_id; // @[Decoupled.scala 298:21]
  assign Queue_io_deq_ready = _T_627_bits_read ? auto_mem_in_r_ready : auto_mem_in_b_ready; // @[Decoupled.scala 320:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  div = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  txen = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  rxen = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  txwm = _RAND_3[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  rxwm = _RAND_4[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  nstop = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  ie_rxwm = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  ie_txwm = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_11 = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_12 = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      div <= 16'had;
    end else if (_T_216) begin
      div <= auto_mem_in_w_bits_data[15:0];
    end
    if (reset) begin
      txen <= 1'h0;
    end else if (_T_239) begin
      txen <= auto_mem_in_w_bits_data[0];
    end
    if (reset) begin
      rxen <= 1'h0;
    end else if (_T_312) begin
      rxen <= auto_mem_in_w_bits_data[0];
    end
    if (reset) begin
      txwm <= 5'h0;
    end else if (_T_287) begin
      txwm <= auto_mem_in_w_bits_data[20:16];
    end
    if (reset) begin
      rxwm <= 5'h0;
    end else if (_T_335) begin
      rxwm <= auto_mem_in_w_bits_data[20:16];
    end
    if (reset) begin
      nstop <= 1'h0;
    end else if (_T_262) begin
      nstop <= auto_mem_in_w_bits_data[1];
    end
    if (reset) begin
      ie_rxwm <= 1'h0;
    end else if (_T_383) begin
      ie_rxwm <= auto_mem_in_w_bits_data[1];
    end
    if (reset) begin
      ie_txwm <= 1'h0;
    end else if (_T_360) begin
      ie_txwm <= auto_mem_in_w_bits_data[0];
    end
    if (reset) begin
      _T_11 <= 32'h0;
    end else if (_T_122) begin
      _T_11 <= auto_mem_in_w_bits_data;
    end
    if (reset) begin
      _T_12 <= 32'h0;
    end else if (_T_193) begin
      _T_12 <= auto_mem_in_w_bits_data;
    end
  end
endmodule
module QueueCompatibility_8(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [20:0] io_enq_bits,
  input         io_deq_ready,
  output        io_deq_valid,
  output [20:0] io_deq_bits
);
  reg [20:0] _T [0:1]; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_0;
  wire [20:0] _T__T_18_data; // @[Decoupled.scala 218:24]
  wire  _T__T_18_addr; // @[Decoupled.scala 218:24]
  wire [20:0] _T__T_10_data; // @[Decoupled.scala 218:24]
  wire  _T__T_10_addr; // @[Decoupled.scala 218:24]
  wire  _T__T_10_mask; // @[Decoupled.scala 218:24]
  wire  _T__T_10_en; // @[Decoupled.scala 218:24]
  reg  value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_1;
  reg  value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_2;
  reg  _T_1; // @[Decoupled.scala 221:35]
  reg [31:0] _RAND_3;
  wire  _T_2 = value == value_1; // @[Decoupled.scala 223:41]
  wire  _T_3 = ~_T_1; // @[Decoupled.scala 224:36]
  wire  _T_4 = _T_2 & _T_3; // @[Decoupled.scala 224:33]
  wire  _T_5 = _T_2 & _T_1; // @[Decoupled.scala 225:32]
  wire  _T_6 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  _T_8 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire  _T_12 = value + 1'h1; // @[Counter.scala 39:22]
  wire  _GEN_9 = io_deq_ready ? 1'h0 : _T_6; // @[Decoupled.scala 249:27]
  wire  _GEN_12 = _T_4 ? _GEN_9 : _T_6; // @[Decoupled.scala 246:18]
  wire  _T_14 = value_1 + 1'h1; // @[Counter.scala 39:22]
  wire  _GEN_11 = _T_4 ? 1'h0 : _T_8; // @[Decoupled.scala 246:18]
  wire  _T_15 = _GEN_12 != _GEN_11; // @[Decoupled.scala 236:16]
  wire  _T_16 = ~_T_4; // @[Decoupled.scala 240:19]
  assign _T__T_18_addr = value_1;
  assign _T__T_18_data = _T[_T__T_18_addr]; // @[Decoupled.scala 218:24]
  assign _T__T_10_data = io_enq_bits;
  assign _T__T_10_addr = value;
  assign _T__T_10_mask = 1'h1;
  assign _T__T_10_en = _T_4 ? _GEN_9 : _T_6;
  assign io_enq_ready = ~_T_5; // @[Decoupled.scala 241:16]
  assign io_deq_valid = io_enq_valid | _T_16; // @[Decoupled.scala 240:16 Decoupled.scala 245:40]
  assign io_deq_bits = _T_4 ? io_enq_bits : _T__T_18_data; // @[Decoupled.scala 242:15 Decoupled.scala 247:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T[initvar] = _RAND_0[20:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  value = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  value_1 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_1 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T__T_10_en & _T__T_10_mask) begin
      _T[_T__T_10_addr] <= _T__T_10_data; // @[Decoupled.scala 218:24]
    end
    if (reset) begin
      value <= 1'h0;
    end else if (_GEN_12) begin
      value <= _T_12;
    end
    if (reset) begin
      value_1 <= 1'h0;
    end else if (_GEN_11) begin
      value_1 <= _T_14;
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else if (_T_15) begin
      if (_T_4) begin
        if (io_deq_ready) begin
          _T_1 <= 1'h0;
        end else begin
          _T_1 <= _T_6;
        end
      end else begin
        _T_1 <= _T_6;
      end
    end
  end
endmodule
module AXI4Xbar_2(
  input         clock,
  input         reset,
  output        auto_in_aw_ready,
  input         auto_in_aw_valid,
  input         auto_in_aw_bits_id,
  input  [29:0] auto_in_aw_bits_addr,
  input  [2:0]  auto_in_aw_bits_size,
  output        auto_in_w_ready,
  input         auto_in_w_valid,
  input  [31:0] auto_in_w_bits_data,
  input  [3:0]  auto_in_w_bits_strb,
  input         auto_in_w_bits_last,
  input         auto_in_b_ready,
  output        auto_in_b_valid,
  output [1:0]  auto_in_b_bits_resp,
  output        auto_in_ar_ready,
  input         auto_in_ar_valid,
  input         auto_in_ar_bits_id,
  input  [29:0] auto_in_ar_bits_addr,
  input  [2:0]  auto_in_ar_bits_size,
  input         auto_in_r_ready,
  output        auto_in_r_valid,
  output [31:0] auto_in_r_bits_data,
  output [1:0]  auto_in_r_bits_resp,
  output        auto_in_r_bits_last,
  input         auto_out_20_aw_ready,
  output        auto_out_20_aw_valid,
  output        auto_out_20_aw_bits_id,
  output [29:0] auto_out_20_aw_bits_addr,
  output [2:0]  auto_out_20_aw_bits_size,
  input         auto_out_20_w_ready,
  output        auto_out_20_w_valid,
  output [31:0] auto_out_20_w_bits_data,
  output [3:0]  auto_out_20_w_bits_strb,
  output        auto_out_20_w_bits_last,
  output        auto_out_20_b_ready,
  input         auto_out_20_b_valid,
  input  [1:0]  auto_out_20_b_bits_resp,
  input         auto_out_20_ar_ready,
  output        auto_out_20_ar_valid,
  output        auto_out_20_ar_bits_id,
  output [29:0] auto_out_20_ar_bits_addr,
  output [2:0]  auto_out_20_ar_bits_size,
  output        auto_out_20_r_ready,
  input         auto_out_20_r_valid,
  input  [31:0] auto_out_20_r_bits_data,
  input  [1:0]  auto_out_20_r_bits_resp,
  input         auto_out_20_r_bits_last,
  input         auto_out_19_aw_ready,
  output        auto_out_19_aw_valid,
  output        auto_out_19_aw_bits_id,
  output [29:0] auto_out_19_aw_bits_addr,
  output [2:0]  auto_out_19_aw_bits_size,
  input         auto_out_19_w_ready,
  output        auto_out_19_w_valid,
  output [31:0] auto_out_19_w_bits_data,
  output [3:0]  auto_out_19_w_bits_strb,
  output        auto_out_19_w_bits_last,
  output        auto_out_19_b_ready,
  input         auto_out_19_b_valid,
  input         auto_out_19_b_bits_id,
  input  [1:0]  auto_out_19_b_bits_resp,
  input         auto_out_19_ar_ready,
  output        auto_out_19_ar_valid,
  output        auto_out_19_ar_bits_id,
  output [29:0] auto_out_19_ar_bits_addr,
  output [2:0]  auto_out_19_ar_bits_size,
  output        auto_out_19_r_ready,
  input         auto_out_19_r_valid,
  input         auto_out_19_r_bits_id,
  input  [31:0] auto_out_19_r_bits_data,
  input  [1:0]  auto_out_19_r_bits_resp,
  input         auto_out_19_r_bits_last,
  input         auto_out_18_aw_ready,
  output        auto_out_18_aw_valid,
  output        auto_out_18_aw_bits_id,
  output [29:0] auto_out_18_aw_bits_addr,
  output [2:0]  auto_out_18_aw_bits_size,
  input         auto_out_18_w_ready,
  output        auto_out_18_w_valid,
  output [31:0] auto_out_18_w_bits_data,
  output [3:0]  auto_out_18_w_bits_strb,
  output        auto_out_18_w_bits_last,
  output        auto_out_18_b_ready,
  input         auto_out_18_b_valid,
  input         auto_out_18_b_bits_id,
  input  [1:0]  auto_out_18_b_bits_resp,
  input         auto_out_18_ar_ready,
  output        auto_out_18_ar_valid,
  output        auto_out_18_ar_bits_id,
  output [29:0] auto_out_18_ar_bits_addr,
  output [2:0]  auto_out_18_ar_bits_size,
  output        auto_out_18_r_ready,
  input         auto_out_18_r_valid,
  input         auto_out_18_r_bits_id,
  input  [31:0] auto_out_18_r_bits_data,
  input  [1:0]  auto_out_18_r_bits_resp,
  input         auto_out_18_r_bits_last,
  input         auto_out_17_aw_ready,
  output        auto_out_17_aw_valid,
  output        auto_out_17_aw_bits_id,
  output [29:0] auto_out_17_aw_bits_addr,
  output [2:0]  auto_out_17_aw_bits_size,
  input         auto_out_17_w_ready,
  output        auto_out_17_w_valid,
  output [31:0] auto_out_17_w_bits_data,
  output [3:0]  auto_out_17_w_bits_strb,
  output        auto_out_17_w_bits_last,
  output        auto_out_17_b_ready,
  input         auto_out_17_b_valid,
  input         auto_out_17_b_bits_id,
  input  [1:0]  auto_out_17_b_bits_resp,
  input         auto_out_17_ar_ready,
  output        auto_out_17_ar_valid,
  output        auto_out_17_ar_bits_id,
  output [29:0] auto_out_17_ar_bits_addr,
  output [2:0]  auto_out_17_ar_bits_size,
  output        auto_out_17_r_ready,
  input         auto_out_17_r_valid,
  input         auto_out_17_r_bits_id,
  input  [31:0] auto_out_17_r_bits_data,
  input  [1:0]  auto_out_17_r_bits_resp,
  input         auto_out_17_r_bits_last,
  input         auto_out_16_aw_ready,
  output        auto_out_16_aw_valid,
  output        auto_out_16_aw_bits_id,
  output [29:0] auto_out_16_aw_bits_addr,
  output [2:0]  auto_out_16_aw_bits_size,
  input         auto_out_16_w_ready,
  output        auto_out_16_w_valid,
  output [31:0] auto_out_16_w_bits_data,
  output [3:0]  auto_out_16_w_bits_strb,
  output        auto_out_16_w_bits_last,
  output        auto_out_16_b_ready,
  input         auto_out_16_b_valid,
  input         auto_out_16_b_bits_id,
  input  [1:0]  auto_out_16_b_bits_resp,
  input         auto_out_16_ar_ready,
  output        auto_out_16_ar_valid,
  output        auto_out_16_ar_bits_id,
  output [29:0] auto_out_16_ar_bits_addr,
  output [2:0]  auto_out_16_ar_bits_size,
  output        auto_out_16_r_ready,
  input         auto_out_16_r_valid,
  input         auto_out_16_r_bits_id,
  input  [31:0] auto_out_16_r_bits_data,
  input  [1:0]  auto_out_16_r_bits_resp,
  input         auto_out_16_r_bits_last,
  input         auto_out_15_aw_ready,
  output        auto_out_15_aw_valid,
  output        auto_out_15_aw_bits_id,
  output [29:0] auto_out_15_aw_bits_addr,
  output [2:0]  auto_out_15_aw_bits_size,
  input         auto_out_15_w_ready,
  output        auto_out_15_w_valid,
  output [31:0] auto_out_15_w_bits_data,
  output [3:0]  auto_out_15_w_bits_strb,
  output        auto_out_15_w_bits_last,
  output        auto_out_15_b_ready,
  input         auto_out_15_b_valid,
  input         auto_out_15_b_bits_id,
  input  [1:0]  auto_out_15_b_bits_resp,
  input         auto_out_15_ar_ready,
  output        auto_out_15_ar_valid,
  output        auto_out_15_ar_bits_id,
  output [29:0] auto_out_15_ar_bits_addr,
  output [2:0]  auto_out_15_ar_bits_size,
  output        auto_out_15_r_ready,
  input         auto_out_15_r_valid,
  input         auto_out_15_r_bits_id,
  input  [31:0] auto_out_15_r_bits_data,
  input  [1:0]  auto_out_15_r_bits_resp,
  input         auto_out_15_r_bits_last,
  input         auto_out_14_aw_ready,
  output        auto_out_14_aw_valid,
  output        auto_out_14_aw_bits_id,
  output [29:0] auto_out_14_aw_bits_addr,
  output [2:0]  auto_out_14_aw_bits_size,
  input         auto_out_14_w_ready,
  output        auto_out_14_w_valid,
  output [31:0] auto_out_14_w_bits_data,
  output [3:0]  auto_out_14_w_bits_strb,
  output        auto_out_14_w_bits_last,
  output        auto_out_14_b_ready,
  input         auto_out_14_b_valid,
  input         auto_out_14_b_bits_id,
  input  [1:0]  auto_out_14_b_bits_resp,
  input         auto_out_14_ar_ready,
  output        auto_out_14_ar_valid,
  output        auto_out_14_ar_bits_id,
  output [29:0] auto_out_14_ar_bits_addr,
  output [2:0]  auto_out_14_ar_bits_size,
  output        auto_out_14_r_ready,
  input         auto_out_14_r_valid,
  input         auto_out_14_r_bits_id,
  input  [31:0] auto_out_14_r_bits_data,
  input  [1:0]  auto_out_14_r_bits_resp,
  input         auto_out_14_r_bits_last,
  input         auto_out_13_aw_ready,
  output        auto_out_13_aw_valid,
  output        auto_out_13_aw_bits_id,
  output [29:0] auto_out_13_aw_bits_addr,
  output [2:0]  auto_out_13_aw_bits_size,
  input         auto_out_13_w_ready,
  output        auto_out_13_w_valid,
  output [31:0] auto_out_13_w_bits_data,
  output [3:0]  auto_out_13_w_bits_strb,
  output        auto_out_13_w_bits_last,
  output        auto_out_13_b_ready,
  input         auto_out_13_b_valid,
  input         auto_out_13_b_bits_id,
  input  [1:0]  auto_out_13_b_bits_resp,
  input         auto_out_13_ar_ready,
  output        auto_out_13_ar_valid,
  output        auto_out_13_ar_bits_id,
  output [29:0] auto_out_13_ar_bits_addr,
  output [2:0]  auto_out_13_ar_bits_size,
  output        auto_out_13_r_ready,
  input         auto_out_13_r_valid,
  input         auto_out_13_r_bits_id,
  input  [31:0] auto_out_13_r_bits_data,
  input  [1:0]  auto_out_13_r_bits_resp,
  input         auto_out_13_r_bits_last,
  input         auto_out_12_aw_ready,
  output        auto_out_12_aw_valid,
  output        auto_out_12_aw_bits_id,
  output [29:0] auto_out_12_aw_bits_addr,
  output [2:0]  auto_out_12_aw_bits_size,
  input         auto_out_12_w_ready,
  output        auto_out_12_w_valid,
  output [31:0] auto_out_12_w_bits_data,
  output [3:0]  auto_out_12_w_bits_strb,
  output        auto_out_12_w_bits_last,
  output        auto_out_12_b_ready,
  input         auto_out_12_b_valid,
  input         auto_out_12_b_bits_id,
  input  [1:0]  auto_out_12_b_bits_resp,
  input         auto_out_12_ar_ready,
  output        auto_out_12_ar_valid,
  output        auto_out_12_ar_bits_id,
  output [29:0] auto_out_12_ar_bits_addr,
  output [2:0]  auto_out_12_ar_bits_size,
  output        auto_out_12_r_ready,
  input         auto_out_12_r_valid,
  input         auto_out_12_r_bits_id,
  input  [31:0] auto_out_12_r_bits_data,
  input  [1:0]  auto_out_12_r_bits_resp,
  input         auto_out_12_r_bits_last,
  input         auto_out_11_aw_ready,
  output        auto_out_11_aw_valid,
  output        auto_out_11_aw_bits_id,
  output [29:0] auto_out_11_aw_bits_addr,
  output [2:0]  auto_out_11_aw_bits_size,
  input         auto_out_11_w_ready,
  output        auto_out_11_w_valid,
  output [31:0] auto_out_11_w_bits_data,
  output [3:0]  auto_out_11_w_bits_strb,
  output        auto_out_11_w_bits_last,
  output        auto_out_11_b_ready,
  input         auto_out_11_b_valid,
  input         auto_out_11_b_bits_id,
  input  [1:0]  auto_out_11_b_bits_resp,
  input         auto_out_11_ar_ready,
  output        auto_out_11_ar_valid,
  output        auto_out_11_ar_bits_id,
  output [29:0] auto_out_11_ar_bits_addr,
  output [2:0]  auto_out_11_ar_bits_size,
  output        auto_out_11_r_ready,
  input         auto_out_11_r_valid,
  input         auto_out_11_r_bits_id,
  input  [31:0] auto_out_11_r_bits_data,
  input  [1:0]  auto_out_11_r_bits_resp,
  input         auto_out_11_r_bits_last,
  input         auto_out_10_aw_ready,
  output        auto_out_10_aw_valid,
  output        auto_out_10_aw_bits_id,
  output [29:0] auto_out_10_aw_bits_addr,
  output [2:0]  auto_out_10_aw_bits_size,
  input         auto_out_10_w_ready,
  output        auto_out_10_w_valid,
  output [31:0] auto_out_10_w_bits_data,
  output [3:0]  auto_out_10_w_bits_strb,
  output        auto_out_10_w_bits_last,
  output        auto_out_10_b_ready,
  input         auto_out_10_b_valid,
  input         auto_out_10_b_bits_id,
  input  [1:0]  auto_out_10_b_bits_resp,
  input         auto_out_10_ar_ready,
  output        auto_out_10_ar_valid,
  output        auto_out_10_ar_bits_id,
  output [29:0] auto_out_10_ar_bits_addr,
  output [2:0]  auto_out_10_ar_bits_size,
  output        auto_out_10_r_ready,
  input         auto_out_10_r_valid,
  input         auto_out_10_r_bits_id,
  input  [31:0] auto_out_10_r_bits_data,
  input  [1:0]  auto_out_10_r_bits_resp,
  input         auto_out_10_r_bits_last,
  input         auto_out_9_aw_ready,
  output        auto_out_9_aw_valid,
  output        auto_out_9_aw_bits_id,
  output [29:0] auto_out_9_aw_bits_addr,
  output [2:0]  auto_out_9_aw_bits_size,
  input         auto_out_9_w_ready,
  output        auto_out_9_w_valid,
  output [31:0] auto_out_9_w_bits_data,
  output [3:0]  auto_out_9_w_bits_strb,
  output        auto_out_9_w_bits_last,
  output        auto_out_9_b_ready,
  input         auto_out_9_b_valid,
  input         auto_out_9_b_bits_id,
  input  [1:0]  auto_out_9_b_bits_resp,
  input         auto_out_9_ar_ready,
  output        auto_out_9_ar_valid,
  output        auto_out_9_ar_bits_id,
  output [29:0] auto_out_9_ar_bits_addr,
  output [2:0]  auto_out_9_ar_bits_size,
  output        auto_out_9_r_ready,
  input         auto_out_9_r_valid,
  input         auto_out_9_r_bits_id,
  input  [31:0] auto_out_9_r_bits_data,
  input  [1:0]  auto_out_9_r_bits_resp,
  input         auto_out_9_r_bits_last,
  input         auto_out_8_aw_ready,
  output        auto_out_8_aw_valid,
  output        auto_out_8_aw_bits_id,
  output [29:0] auto_out_8_aw_bits_addr,
  output [2:0]  auto_out_8_aw_bits_size,
  input         auto_out_8_w_ready,
  output        auto_out_8_w_valid,
  output [31:0] auto_out_8_w_bits_data,
  output [3:0]  auto_out_8_w_bits_strb,
  output        auto_out_8_w_bits_last,
  output        auto_out_8_b_ready,
  input         auto_out_8_b_valid,
  input         auto_out_8_b_bits_id,
  input  [1:0]  auto_out_8_b_bits_resp,
  input         auto_out_8_ar_ready,
  output        auto_out_8_ar_valid,
  output        auto_out_8_ar_bits_id,
  output [29:0] auto_out_8_ar_bits_addr,
  output [2:0]  auto_out_8_ar_bits_size,
  output        auto_out_8_r_ready,
  input         auto_out_8_r_valid,
  input         auto_out_8_r_bits_id,
  input  [31:0] auto_out_8_r_bits_data,
  input  [1:0]  auto_out_8_r_bits_resp,
  input         auto_out_8_r_bits_last,
  input         auto_out_7_aw_ready,
  output        auto_out_7_aw_valid,
  output        auto_out_7_aw_bits_id,
  output [29:0] auto_out_7_aw_bits_addr,
  output [2:0]  auto_out_7_aw_bits_size,
  input         auto_out_7_w_ready,
  output        auto_out_7_w_valid,
  output [31:0] auto_out_7_w_bits_data,
  output [3:0]  auto_out_7_w_bits_strb,
  output        auto_out_7_w_bits_last,
  output        auto_out_7_b_ready,
  input         auto_out_7_b_valid,
  input         auto_out_7_b_bits_id,
  input  [1:0]  auto_out_7_b_bits_resp,
  input         auto_out_7_ar_ready,
  output        auto_out_7_ar_valid,
  output        auto_out_7_ar_bits_id,
  output [29:0] auto_out_7_ar_bits_addr,
  output [2:0]  auto_out_7_ar_bits_size,
  output        auto_out_7_r_ready,
  input         auto_out_7_r_valid,
  input         auto_out_7_r_bits_id,
  input  [31:0] auto_out_7_r_bits_data,
  input  [1:0]  auto_out_7_r_bits_resp,
  input         auto_out_7_r_bits_last,
  input         auto_out_6_aw_ready,
  output        auto_out_6_aw_valid,
  output        auto_out_6_aw_bits_id,
  output [29:0] auto_out_6_aw_bits_addr,
  output [2:0]  auto_out_6_aw_bits_size,
  input         auto_out_6_w_ready,
  output        auto_out_6_w_valid,
  output [31:0] auto_out_6_w_bits_data,
  output [3:0]  auto_out_6_w_bits_strb,
  output        auto_out_6_w_bits_last,
  output        auto_out_6_b_ready,
  input         auto_out_6_b_valid,
  input         auto_out_6_b_bits_id,
  input  [1:0]  auto_out_6_b_bits_resp,
  input         auto_out_6_ar_ready,
  output        auto_out_6_ar_valid,
  output        auto_out_6_ar_bits_id,
  output [29:0] auto_out_6_ar_bits_addr,
  output [2:0]  auto_out_6_ar_bits_size,
  output        auto_out_6_r_ready,
  input         auto_out_6_r_valid,
  input         auto_out_6_r_bits_id,
  input  [31:0] auto_out_6_r_bits_data,
  input  [1:0]  auto_out_6_r_bits_resp,
  input         auto_out_6_r_bits_last,
  input         auto_out_5_aw_ready,
  output        auto_out_5_aw_valid,
  output        auto_out_5_aw_bits_id,
  output [29:0] auto_out_5_aw_bits_addr,
  output [2:0]  auto_out_5_aw_bits_size,
  input         auto_out_5_w_ready,
  output        auto_out_5_w_valid,
  output [31:0] auto_out_5_w_bits_data,
  output [3:0]  auto_out_5_w_bits_strb,
  output        auto_out_5_w_bits_last,
  output        auto_out_5_b_ready,
  input         auto_out_5_b_valid,
  input         auto_out_5_b_bits_id,
  input  [1:0]  auto_out_5_b_bits_resp,
  input         auto_out_5_ar_ready,
  output        auto_out_5_ar_valid,
  output        auto_out_5_ar_bits_id,
  output [29:0] auto_out_5_ar_bits_addr,
  output [2:0]  auto_out_5_ar_bits_size,
  output        auto_out_5_r_ready,
  input         auto_out_5_r_valid,
  input         auto_out_5_r_bits_id,
  input  [31:0] auto_out_5_r_bits_data,
  input  [1:0]  auto_out_5_r_bits_resp,
  input         auto_out_5_r_bits_last,
  input         auto_out_4_aw_ready,
  output        auto_out_4_aw_valid,
  output        auto_out_4_aw_bits_id,
  output [29:0] auto_out_4_aw_bits_addr,
  output [2:0]  auto_out_4_aw_bits_size,
  input         auto_out_4_w_ready,
  output        auto_out_4_w_valid,
  output [31:0] auto_out_4_w_bits_data,
  output [3:0]  auto_out_4_w_bits_strb,
  output        auto_out_4_w_bits_last,
  output        auto_out_4_b_ready,
  input         auto_out_4_b_valid,
  input         auto_out_4_b_bits_id,
  input  [1:0]  auto_out_4_b_bits_resp,
  input         auto_out_4_ar_ready,
  output        auto_out_4_ar_valid,
  output        auto_out_4_ar_bits_id,
  output [29:0] auto_out_4_ar_bits_addr,
  output [2:0]  auto_out_4_ar_bits_size,
  output        auto_out_4_r_ready,
  input         auto_out_4_r_valid,
  input         auto_out_4_r_bits_id,
  input  [31:0] auto_out_4_r_bits_data,
  input  [1:0]  auto_out_4_r_bits_resp,
  input         auto_out_4_r_bits_last,
  input         auto_out_3_aw_ready,
  output        auto_out_3_aw_valid,
  output        auto_out_3_aw_bits_id,
  output [29:0] auto_out_3_aw_bits_addr,
  output [2:0]  auto_out_3_aw_bits_size,
  input         auto_out_3_w_ready,
  output        auto_out_3_w_valid,
  output [31:0] auto_out_3_w_bits_data,
  output [3:0]  auto_out_3_w_bits_strb,
  output        auto_out_3_w_bits_last,
  output        auto_out_3_b_ready,
  input         auto_out_3_b_valid,
  input         auto_out_3_b_bits_id,
  input  [1:0]  auto_out_3_b_bits_resp,
  input         auto_out_3_ar_ready,
  output        auto_out_3_ar_valid,
  output        auto_out_3_ar_bits_id,
  output [29:0] auto_out_3_ar_bits_addr,
  output [2:0]  auto_out_3_ar_bits_size,
  output        auto_out_3_r_ready,
  input         auto_out_3_r_valid,
  input         auto_out_3_r_bits_id,
  input  [31:0] auto_out_3_r_bits_data,
  input  [1:0]  auto_out_3_r_bits_resp,
  input         auto_out_3_r_bits_last,
  input         auto_out_2_aw_ready,
  output        auto_out_2_aw_valid,
  output        auto_out_2_aw_bits_id,
  output [29:0] auto_out_2_aw_bits_addr,
  output [2:0]  auto_out_2_aw_bits_size,
  input         auto_out_2_w_ready,
  output        auto_out_2_w_valid,
  output [31:0] auto_out_2_w_bits_data,
  output [3:0]  auto_out_2_w_bits_strb,
  output        auto_out_2_w_bits_last,
  output        auto_out_2_b_ready,
  input         auto_out_2_b_valid,
  input         auto_out_2_b_bits_id,
  input  [1:0]  auto_out_2_b_bits_resp,
  input         auto_out_2_ar_ready,
  output        auto_out_2_ar_valid,
  output        auto_out_2_ar_bits_id,
  output [29:0] auto_out_2_ar_bits_addr,
  output [2:0]  auto_out_2_ar_bits_size,
  output        auto_out_2_r_ready,
  input         auto_out_2_r_valid,
  input         auto_out_2_r_bits_id,
  input  [31:0] auto_out_2_r_bits_data,
  input  [1:0]  auto_out_2_r_bits_resp,
  input         auto_out_2_r_bits_last,
  input         auto_out_1_aw_ready,
  output        auto_out_1_aw_valid,
  output        auto_out_1_aw_bits_id,
  output [29:0] auto_out_1_aw_bits_addr,
  output [2:0]  auto_out_1_aw_bits_size,
  input         auto_out_1_w_ready,
  output        auto_out_1_w_valid,
  output [31:0] auto_out_1_w_bits_data,
  output [3:0]  auto_out_1_w_bits_strb,
  output        auto_out_1_w_bits_last,
  output        auto_out_1_b_ready,
  input         auto_out_1_b_valid,
  input         auto_out_1_b_bits_id,
  input  [1:0]  auto_out_1_b_bits_resp,
  input         auto_out_1_ar_ready,
  output        auto_out_1_ar_valid,
  output        auto_out_1_ar_bits_id,
  output [29:0] auto_out_1_ar_bits_addr,
  output [2:0]  auto_out_1_ar_bits_size,
  output        auto_out_1_r_ready,
  input         auto_out_1_r_valid,
  input         auto_out_1_r_bits_id,
  input  [31:0] auto_out_1_r_bits_data,
  input  [1:0]  auto_out_1_r_bits_resp,
  input         auto_out_1_r_bits_last,
  input         auto_out_0_aw_ready,
  output        auto_out_0_aw_valid,
  output        auto_out_0_aw_bits_id,
  output [29:0] auto_out_0_aw_bits_addr,
  output [2:0]  auto_out_0_aw_bits_size,
  input         auto_out_0_w_ready,
  output        auto_out_0_w_valid,
  output [31:0] auto_out_0_w_bits_data,
  output [3:0]  auto_out_0_w_bits_strb,
  output        auto_out_0_w_bits_last,
  output        auto_out_0_b_ready,
  input         auto_out_0_b_valid,
  input         auto_out_0_b_bits_id,
  input  [1:0]  auto_out_0_b_bits_resp,
  input         auto_out_0_ar_ready,
  output        auto_out_0_ar_valid,
  output        auto_out_0_ar_bits_id,
  output [29:0] auto_out_0_ar_bits_addr,
  output [2:0]  auto_out_0_ar_bits_size,
  output        auto_out_0_r_ready,
  input         auto_out_0_r_valid,
  input         auto_out_0_r_bits_id,
  input  [31:0] auto_out_0_r_bits_data,
  input  [1:0]  auto_out_0_r_bits_resp,
  input         auto_out_0_r_bits_last
);
  wire  awIn_0_clock; // @[Xbar.scala 55:47]
  wire  awIn_0_reset; // @[Xbar.scala 55:47]
  wire  awIn_0_io_enq_ready; // @[Xbar.scala 55:47]
  wire  awIn_0_io_enq_valid; // @[Xbar.scala 55:47]
  wire [20:0] awIn_0_io_enq_bits; // @[Xbar.scala 55:47]
  wire  awIn_0_io_deq_ready; // @[Xbar.scala 55:47]
  wire  awIn_0_io_deq_valid; // @[Xbar.scala 55:47]
  wire [20:0] awIn_0_io_deq_bits; // @[Xbar.scala 55:47]
  wire [30:0] _T_1 = {1'b0,$signed(auto_in_ar_bits_addr)}; // @[Parameters.scala 137:49]
  wire [30:0] _T_3 = $signed(_T_1) & 31'shf130; // @[Parameters.scala 137:52]
  wire  requestARIO_0_0 = $signed(_T_3) == 31'sh0; // @[Parameters.scala 137:67]
  wire [29:0] _T_5 = auto_in_ar_bits_addr ^ 30'h1000; // @[Parameters.scala 137:31]
  wire [30:0] _T_6 = {1'b0,$signed(_T_5)}; // @[Parameters.scala 137:49]
  wire [30:0] _T_8 = $signed(_T_6) & 31'shf000; // @[Parameters.scala 137:52]
  wire  _T_9 = $signed(_T_8) == 31'sh0; // @[Parameters.scala 137:67]
  wire [29:0] _T_10 = auto_in_ar_bits_addr ^ 30'h2100; // @[Parameters.scala 137:31]
  wire [30:0] _T_11 = {1'b0,$signed(_T_10)}; // @[Parameters.scala 137:49]
  wire [30:0] _T_13 = $signed(_T_11) & 31'shf100; // @[Parameters.scala 137:52]
  wire  _T_14 = $signed(_T_13) == 31'sh0; // @[Parameters.scala 137:67]
  wire  requestARIO_0_1 = _T_9 | _T_14; // @[Xbar.scala 52:97]
  wire [29:0] _T_16 = auto_in_ar_bits_addr ^ 30'h2000; // @[Parameters.scala 137:31]
  wire [30:0] _T_17 = {1'b0,$signed(_T_16)}; // @[Parameters.scala 137:49]
  wire [30:0] _T_19 = $signed(_T_17) & 31'shf130; // @[Parameters.scala 137:52]
  wire  requestARIO_0_2 = $signed(_T_19) == 31'sh0; // @[Parameters.scala 137:67]
  wire [29:0] _T_21 = auto_in_ar_bits_addr ^ 30'h2010; // @[Parameters.scala 137:31]
  wire [30:0] _T_22 = {1'b0,$signed(_T_21)}; // @[Parameters.scala 137:49]
  wire [30:0] _T_24 = $signed(_T_22) & 31'shf130; // @[Parameters.scala 137:52]
  wire  requestARIO_0_3 = $signed(_T_24) == 31'sh0; // @[Parameters.scala 137:67]
  wire [29:0] _T_26 = auto_in_ar_bits_addr ^ 30'h2020; // @[Parameters.scala 137:31]
  wire [30:0] _T_27 = {1'b0,$signed(_T_26)}; // @[Parameters.scala 137:49]
  wire [30:0] _T_29 = $signed(_T_27) & 31'shf130; // @[Parameters.scala 137:52]
  wire  requestARIO_0_4 = $signed(_T_29) == 31'sh0; // @[Parameters.scala 137:67]
  wire [29:0] _T_31 = auto_in_ar_bits_addr ^ 30'h3000; // @[Parameters.scala 137:31]
  wire [30:0] _T_32 = {1'b0,$signed(_T_31)}; // @[Parameters.scala 137:49]
  wire [30:0] _T_34 = $signed(_T_32) & 31'shf130; // @[Parameters.scala 137:52]
  wire  requestARIO_0_5 = $signed(_T_34) == 31'sh0; // @[Parameters.scala 137:67]
  wire [29:0] _T_36 = auto_in_ar_bits_addr ^ 30'h3100; // @[Parameters.scala 137:31]
  wire [30:0] _T_37 = {1'b0,$signed(_T_36)}; // @[Parameters.scala 137:49]
  wire [30:0] _T_39 = $signed(_T_37) & 31'shf130; // @[Parameters.scala 137:52]
  wire  requestARIO_0_6 = $signed(_T_39) == 31'sh0; // @[Parameters.scala 137:67]
  wire [29:0] _T_41 = auto_in_ar_bits_addr ^ 30'h3110; // @[Parameters.scala 137:31]
  wire [30:0] _T_42 = {1'b0,$signed(_T_41)}; // @[Parameters.scala 137:49]
  wire [30:0] _T_44 = $signed(_T_42) & 31'shf130; // @[Parameters.scala 137:52]
  wire  requestARIO_0_7 = $signed(_T_44) == 31'sh0; // @[Parameters.scala 137:67]
  wire [29:0] _T_46 = auto_in_ar_bits_addr ^ 30'h3120; // @[Parameters.scala 137:31]
  wire [30:0] _T_47 = {1'b0,$signed(_T_46)}; // @[Parameters.scala 137:49]
  wire [30:0] _T_49 = $signed(_T_47) & 31'shf130; // @[Parameters.scala 137:52]
  wire  requestARIO_0_8 = $signed(_T_49) == 31'sh0; // @[Parameters.scala 137:67]
  wire [29:0] _T_51 = auto_in_ar_bits_addr ^ 30'h4000; // @[Parameters.scala 137:31]
  wire [30:0] _T_52 = {1'b0,$signed(_T_51)}; // @[Parameters.scala 137:49]
  wire [30:0] _T_54 = $signed(_T_52) & 31'shf100; // @[Parameters.scala 137:52]
  wire  requestARIO_0_9 = $signed(_T_54) == 31'sh0; // @[Parameters.scala 137:67]
  wire [29:0] _T_56 = auto_in_ar_bits_addr ^ 30'h4100; // @[Parameters.scala 137:31]
  wire [30:0] _T_57 = {1'b0,$signed(_T_56)}; // @[Parameters.scala 137:49]
  wire [30:0] _T_59 = $signed(_T_57) & 31'shf130; // @[Parameters.scala 137:52]
  wire  requestARIO_0_10 = $signed(_T_59) == 31'sh0; // @[Parameters.scala 137:67]
  wire [29:0] _T_61 = auto_in_ar_bits_addr ^ 30'h4110; // @[Parameters.scala 137:31]
  wire [30:0] _T_62 = {1'b0,$signed(_T_61)}; // @[Parameters.scala 137:49]
  wire [30:0] _T_64 = $signed(_T_62) & 31'shf130; // @[Parameters.scala 137:52]
  wire  requestARIO_0_11 = $signed(_T_64) == 31'sh0; // @[Parameters.scala 137:67]
  wire [29:0] _T_66 = auto_in_ar_bits_addr ^ 30'h4120; // @[Parameters.scala 137:31]
  wire [30:0] _T_67 = {1'b0,$signed(_T_66)}; // @[Parameters.scala 137:49]
  wire [30:0] _T_69 = $signed(_T_67) & 31'shf130; // @[Parameters.scala 137:52]
  wire  requestARIO_0_12 = $signed(_T_69) == 31'sh0; // @[Parameters.scala 137:67]
  wire [29:0] _T_71 = auto_in_ar_bits_addr ^ 30'h5000; // @[Parameters.scala 137:31]
  wire [30:0] _T_72 = {1'b0,$signed(_T_71)}; // @[Parameters.scala 137:49]
  wire [30:0] _T_74 = $signed(_T_72) & 31'shf100; // @[Parameters.scala 137:52]
  wire  requestARIO_0_13 = $signed(_T_74) == 31'sh0; // @[Parameters.scala 137:67]
  wire [29:0] _T_76 = auto_in_ar_bits_addr ^ 30'h5100; // @[Parameters.scala 137:31]
  wire [30:0] _T_77 = {1'b0,$signed(_T_76)}; // @[Parameters.scala 137:49]
  wire [30:0] _T_79 = $signed(_T_77) & 31'shf130; // @[Parameters.scala 137:52]
  wire  requestARIO_0_14 = $signed(_T_79) == 31'sh0; // @[Parameters.scala 137:67]
  wire [29:0] _T_81 = auto_in_ar_bits_addr ^ 30'h5110; // @[Parameters.scala 137:31]
  wire [30:0] _T_82 = {1'b0,$signed(_T_81)}; // @[Parameters.scala 137:49]
  wire [30:0] _T_84 = $signed(_T_82) & 31'shf130; // @[Parameters.scala 137:52]
  wire  requestARIO_0_15 = $signed(_T_84) == 31'sh0; // @[Parameters.scala 137:67]
  wire [29:0] _T_86 = auto_in_ar_bits_addr ^ 30'h5120; // @[Parameters.scala 137:31]
  wire [30:0] _T_87 = {1'b0,$signed(_T_86)}; // @[Parameters.scala 137:49]
  wire [30:0] _T_89 = $signed(_T_87) & 31'shf130; // @[Parameters.scala 137:52]
  wire  requestARIO_0_16 = $signed(_T_89) == 31'sh0; // @[Parameters.scala 137:67]
  wire [29:0] _T_91 = auto_in_ar_bits_addr ^ 30'h8000; // @[Parameters.scala 137:31]
  wire [30:0] _T_92 = {1'b0,$signed(_T_91)}; // @[Parameters.scala 137:49]
  wire [30:0] _T_94 = $signed(_T_92) & 31'shf130; // @[Parameters.scala 137:52]
  wire  requestARIO_0_17 = $signed(_T_94) == 31'sh0; // @[Parameters.scala 137:67]
  wire [29:0] _T_96 = auto_in_ar_bits_addr ^ 30'h9000; // @[Parameters.scala 137:31]
  wire [30:0] _T_97 = {1'b0,$signed(_T_96)}; // @[Parameters.scala 137:49]
  wire [30:0] _T_99 = $signed(_T_97) & 31'shf100; // @[Parameters.scala 137:52]
  wire  requestARIO_0_18 = $signed(_T_99) == 31'sh0; // @[Parameters.scala 137:67]
  wire [29:0] _T_101 = auto_in_ar_bits_addr ^ 30'h9100; // @[Parameters.scala 137:31]
  wire [30:0] _T_102 = {1'b0,$signed(_T_101)}; // @[Parameters.scala 137:49]
  wire [30:0] _T_104 = $signed(_T_102) & 31'shf130; // @[Parameters.scala 137:52]
  wire  requestARIO_0_19 = $signed(_T_104) == 31'sh0; // @[Parameters.scala 137:67]
  wire [29:0] _T_106 = auto_in_ar_bits_addr ^ 30'h6000; // @[Parameters.scala 137:31]
  wire [30:0] _T_107 = {1'b0,$signed(_T_106)}; // @[Parameters.scala 137:49]
  wire [30:0] _T_109 = $signed(_T_107) & 31'shf000; // @[Parameters.scala 137:52]
  wire  _T_110 = $signed(_T_109) == 31'sh0; // @[Parameters.scala 137:67]
  wire [29:0] _T_111 = auto_in_ar_bits_addr ^ 30'h7000; // @[Parameters.scala 137:31]
  wire [30:0] _T_112 = {1'b0,$signed(_T_111)}; // @[Parameters.scala 137:49]
  wire [30:0] _T_114 = $signed(_T_112) & 31'shf130; // @[Parameters.scala 137:52]
  wire  _T_115 = $signed(_T_114) == 31'sh0; // @[Parameters.scala 137:67]
  wire  requestARIO_0_20 = _T_110 | _T_115; // @[Xbar.scala 52:97]
  wire [30:0] _T_118 = {1'b0,$signed(auto_in_aw_bits_addr)}; // @[Parameters.scala 137:49]
  wire [30:0] _T_120 = $signed(_T_118) & 31'shf130; // @[Parameters.scala 137:52]
  wire  requestAWIO_0_0 = $signed(_T_120) == 31'sh0; // @[Parameters.scala 137:67]
  wire [29:0] _T_122 = auto_in_aw_bits_addr ^ 30'h1000; // @[Parameters.scala 137:31]
  wire [30:0] _T_123 = {1'b0,$signed(_T_122)}; // @[Parameters.scala 137:49]
  wire [30:0] _T_125 = $signed(_T_123) & 31'shf000; // @[Parameters.scala 137:52]
  wire  _T_126 = $signed(_T_125) == 31'sh0; // @[Parameters.scala 137:67]
  wire [29:0] _T_127 = auto_in_aw_bits_addr ^ 30'h2100; // @[Parameters.scala 137:31]
  wire [30:0] _T_128 = {1'b0,$signed(_T_127)}; // @[Parameters.scala 137:49]
  wire [30:0] _T_130 = $signed(_T_128) & 31'shf100; // @[Parameters.scala 137:52]
  wire  _T_131 = $signed(_T_130) == 31'sh0; // @[Parameters.scala 137:67]
  wire  requestAWIO_0_1 = _T_126 | _T_131; // @[Xbar.scala 52:97]
  wire [29:0] _T_133 = auto_in_aw_bits_addr ^ 30'h2000; // @[Parameters.scala 137:31]
  wire [30:0] _T_134 = {1'b0,$signed(_T_133)}; // @[Parameters.scala 137:49]
  wire [30:0] _T_136 = $signed(_T_134) & 31'shf130; // @[Parameters.scala 137:52]
  wire  requestAWIO_0_2 = $signed(_T_136) == 31'sh0; // @[Parameters.scala 137:67]
  wire [29:0] _T_138 = auto_in_aw_bits_addr ^ 30'h2010; // @[Parameters.scala 137:31]
  wire [30:0] _T_139 = {1'b0,$signed(_T_138)}; // @[Parameters.scala 137:49]
  wire [30:0] _T_141 = $signed(_T_139) & 31'shf130; // @[Parameters.scala 137:52]
  wire  requestAWIO_0_3 = $signed(_T_141) == 31'sh0; // @[Parameters.scala 137:67]
  wire [29:0] _T_143 = auto_in_aw_bits_addr ^ 30'h2020; // @[Parameters.scala 137:31]
  wire [30:0] _T_144 = {1'b0,$signed(_T_143)}; // @[Parameters.scala 137:49]
  wire [30:0] _T_146 = $signed(_T_144) & 31'shf130; // @[Parameters.scala 137:52]
  wire  requestAWIO_0_4 = $signed(_T_146) == 31'sh0; // @[Parameters.scala 137:67]
  wire [29:0] _T_148 = auto_in_aw_bits_addr ^ 30'h3000; // @[Parameters.scala 137:31]
  wire [30:0] _T_149 = {1'b0,$signed(_T_148)}; // @[Parameters.scala 137:49]
  wire [30:0] _T_151 = $signed(_T_149) & 31'shf130; // @[Parameters.scala 137:52]
  wire  requestAWIO_0_5 = $signed(_T_151) == 31'sh0; // @[Parameters.scala 137:67]
  wire [29:0] _T_153 = auto_in_aw_bits_addr ^ 30'h3100; // @[Parameters.scala 137:31]
  wire [30:0] _T_154 = {1'b0,$signed(_T_153)}; // @[Parameters.scala 137:49]
  wire [30:0] _T_156 = $signed(_T_154) & 31'shf130; // @[Parameters.scala 137:52]
  wire  requestAWIO_0_6 = $signed(_T_156) == 31'sh0; // @[Parameters.scala 137:67]
  wire [29:0] _T_158 = auto_in_aw_bits_addr ^ 30'h3110; // @[Parameters.scala 137:31]
  wire [30:0] _T_159 = {1'b0,$signed(_T_158)}; // @[Parameters.scala 137:49]
  wire [30:0] _T_161 = $signed(_T_159) & 31'shf130; // @[Parameters.scala 137:52]
  wire  requestAWIO_0_7 = $signed(_T_161) == 31'sh0; // @[Parameters.scala 137:67]
  wire [29:0] _T_163 = auto_in_aw_bits_addr ^ 30'h3120; // @[Parameters.scala 137:31]
  wire [30:0] _T_164 = {1'b0,$signed(_T_163)}; // @[Parameters.scala 137:49]
  wire [30:0] _T_166 = $signed(_T_164) & 31'shf130; // @[Parameters.scala 137:52]
  wire  requestAWIO_0_8 = $signed(_T_166) == 31'sh0; // @[Parameters.scala 137:67]
  wire [29:0] _T_168 = auto_in_aw_bits_addr ^ 30'h4000; // @[Parameters.scala 137:31]
  wire [30:0] _T_169 = {1'b0,$signed(_T_168)}; // @[Parameters.scala 137:49]
  wire [30:0] _T_171 = $signed(_T_169) & 31'shf100; // @[Parameters.scala 137:52]
  wire  requestAWIO_0_9 = $signed(_T_171) == 31'sh0; // @[Parameters.scala 137:67]
  wire [29:0] _T_173 = auto_in_aw_bits_addr ^ 30'h4100; // @[Parameters.scala 137:31]
  wire [30:0] _T_174 = {1'b0,$signed(_T_173)}; // @[Parameters.scala 137:49]
  wire [30:0] _T_176 = $signed(_T_174) & 31'shf130; // @[Parameters.scala 137:52]
  wire  requestAWIO_0_10 = $signed(_T_176) == 31'sh0; // @[Parameters.scala 137:67]
  wire [29:0] _T_178 = auto_in_aw_bits_addr ^ 30'h4110; // @[Parameters.scala 137:31]
  wire [30:0] _T_179 = {1'b0,$signed(_T_178)}; // @[Parameters.scala 137:49]
  wire [30:0] _T_181 = $signed(_T_179) & 31'shf130; // @[Parameters.scala 137:52]
  wire  requestAWIO_0_11 = $signed(_T_181) == 31'sh0; // @[Parameters.scala 137:67]
  wire [29:0] _T_183 = auto_in_aw_bits_addr ^ 30'h4120; // @[Parameters.scala 137:31]
  wire [30:0] _T_184 = {1'b0,$signed(_T_183)}; // @[Parameters.scala 137:49]
  wire [30:0] _T_186 = $signed(_T_184) & 31'shf130; // @[Parameters.scala 137:52]
  wire  requestAWIO_0_12 = $signed(_T_186) == 31'sh0; // @[Parameters.scala 137:67]
  wire [29:0] _T_188 = auto_in_aw_bits_addr ^ 30'h5000; // @[Parameters.scala 137:31]
  wire [30:0] _T_189 = {1'b0,$signed(_T_188)}; // @[Parameters.scala 137:49]
  wire [30:0] _T_191 = $signed(_T_189) & 31'shf100; // @[Parameters.scala 137:52]
  wire  requestAWIO_0_13 = $signed(_T_191) == 31'sh0; // @[Parameters.scala 137:67]
  wire [29:0] _T_193 = auto_in_aw_bits_addr ^ 30'h5100; // @[Parameters.scala 137:31]
  wire [30:0] _T_194 = {1'b0,$signed(_T_193)}; // @[Parameters.scala 137:49]
  wire [30:0] _T_196 = $signed(_T_194) & 31'shf130; // @[Parameters.scala 137:52]
  wire  requestAWIO_0_14 = $signed(_T_196) == 31'sh0; // @[Parameters.scala 137:67]
  wire [29:0] _T_198 = auto_in_aw_bits_addr ^ 30'h5110; // @[Parameters.scala 137:31]
  wire [30:0] _T_199 = {1'b0,$signed(_T_198)}; // @[Parameters.scala 137:49]
  wire [30:0] _T_201 = $signed(_T_199) & 31'shf130; // @[Parameters.scala 137:52]
  wire  requestAWIO_0_15 = $signed(_T_201) == 31'sh0; // @[Parameters.scala 137:67]
  wire [29:0] _T_203 = auto_in_aw_bits_addr ^ 30'h5120; // @[Parameters.scala 137:31]
  wire [30:0] _T_204 = {1'b0,$signed(_T_203)}; // @[Parameters.scala 137:49]
  wire [30:0] _T_206 = $signed(_T_204) & 31'shf130; // @[Parameters.scala 137:52]
  wire  requestAWIO_0_16 = $signed(_T_206) == 31'sh0; // @[Parameters.scala 137:67]
  wire [29:0] _T_208 = auto_in_aw_bits_addr ^ 30'h8000; // @[Parameters.scala 137:31]
  wire [30:0] _T_209 = {1'b0,$signed(_T_208)}; // @[Parameters.scala 137:49]
  wire [30:0] _T_211 = $signed(_T_209) & 31'shf130; // @[Parameters.scala 137:52]
  wire  requestAWIO_0_17 = $signed(_T_211) == 31'sh0; // @[Parameters.scala 137:67]
  wire [29:0] _T_213 = auto_in_aw_bits_addr ^ 30'h9000; // @[Parameters.scala 137:31]
  wire [30:0] _T_214 = {1'b0,$signed(_T_213)}; // @[Parameters.scala 137:49]
  wire [30:0] _T_216 = $signed(_T_214) & 31'shf100; // @[Parameters.scala 137:52]
  wire  requestAWIO_0_18 = $signed(_T_216) == 31'sh0; // @[Parameters.scala 137:67]
  wire [29:0] _T_218 = auto_in_aw_bits_addr ^ 30'h9100; // @[Parameters.scala 137:31]
  wire [30:0] _T_219 = {1'b0,$signed(_T_218)}; // @[Parameters.scala 137:49]
  wire [30:0] _T_221 = $signed(_T_219) & 31'shf130; // @[Parameters.scala 137:52]
  wire  requestAWIO_0_19 = $signed(_T_221) == 31'sh0; // @[Parameters.scala 137:67]
  wire [29:0] _T_223 = auto_in_aw_bits_addr ^ 30'h6000; // @[Parameters.scala 137:31]
  wire [30:0] _T_224 = {1'b0,$signed(_T_223)}; // @[Parameters.scala 137:49]
  wire [30:0] _T_226 = $signed(_T_224) & 31'shf000; // @[Parameters.scala 137:52]
  wire  _T_227 = $signed(_T_226) == 31'sh0; // @[Parameters.scala 137:67]
  wire [29:0] _T_228 = auto_in_aw_bits_addr ^ 30'h7000; // @[Parameters.scala 137:31]
  wire [30:0] _T_229 = {1'b0,$signed(_T_228)}; // @[Parameters.scala 137:49]
  wire [30:0] _T_231 = $signed(_T_229) & 31'shf130; // @[Parameters.scala 137:52]
  wire  _T_232 = $signed(_T_231) == 31'sh0; // @[Parameters.scala 137:67]
  wire  requestAWIO_0_20 = _T_227 | _T_232; // @[Xbar.scala 52:97]
  wire  requestROI_0_0 = ~auto_out_0_r_bits_id; // @[Parameters.scala 47:9]
  wire  requestROI_1_0 = ~auto_out_1_r_bits_id; // @[Parameters.scala 47:9]
  wire  requestROI_2_0 = ~auto_out_2_r_bits_id; // @[Parameters.scala 47:9]
  wire  requestROI_3_0 = ~auto_out_3_r_bits_id; // @[Parameters.scala 47:9]
  wire  requestROI_4_0 = ~auto_out_4_r_bits_id; // @[Parameters.scala 47:9]
  wire  requestROI_5_0 = ~auto_out_5_r_bits_id; // @[Parameters.scala 47:9]
  wire  requestROI_6_0 = ~auto_out_6_r_bits_id; // @[Parameters.scala 47:9]
  wire  requestROI_7_0 = ~auto_out_7_r_bits_id; // @[Parameters.scala 47:9]
  wire  requestROI_8_0 = ~auto_out_8_r_bits_id; // @[Parameters.scala 47:9]
  wire  requestROI_9_0 = ~auto_out_9_r_bits_id; // @[Parameters.scala 47:9]
  wire  requestROI_10_0 = ~auto_out_10_r_bits_id; // @[Parameters.scala 47:9]
  wire  requestROI_11_0 = ~auto_out_11_r_bits_id; // @[Parameters.scala 47:9]
  wire  requestROI_12_0 = ~auto_out_12_r_bits_id; // @[Parameters.scala 47:9]
  wire  requestROI_13_0 = ~auto_out_13_r_bits_id; // @[Parameters.scala 47:9]
  wire  requestROI_14_0 = ~auto_out_14_r_bits_id; // @[Parameters.scala 47:9]
  wire  requestROI_15_0 = ~auto_out_15_r_bits_id; // @[Parameters.scala 47:9]
  wire  requestROI_16_0 = ~auto_out_16_r_bits_id; // @[Parameters.scala 47:9]
  wire  requestROI_17_0 = ~auto_out_17_r_bits_id; // @[Parameters.scala 47:9]
  wire  requestROI_18_0 = ~auto_out_18_r_bits_id; // @[Parameters.scala 47:9]
  wire  requestROI_19_0 = ~auto_out_19_r_bits_id; // @[Parameters.scala 47:9]
  wire  requestBOI_0_0 = ~auto_out_0_b_bits_id; // @[Parameters.scala 47:9]
  wire  requestBOI_1_0 = ~auto_out_1_b_bits_id; // @[Parameters.scala 47:9]
  wire  requestBOI_2_0 = ~auto_out_2_b_bits_id; // @[Parameters.scala 47:9]
  wire  requestBOI_3_0 = ~auto_out_3_b_bits_id; // @[Parameters.scala 47:9]
  wire  requestBOI_4_0 = ~auto_out_4_b_bits_id; // @[Parameters.scala 47:9]
  wire  requestBOI_5_0 = ~auto_out_5_b_bits_id; // @[Parameters.scala 47:9]
  wire  requestBOI_6_0 = ~auto_out_6_b_bits_id; // @[Parameters.scala 47:9]
  wire  requestBOI_7_0 = ~auto_out_7_b_bits_id; // @[Parameters.scala 47:9]
  wire  requestBOI_8_0 = ~auto_out_8_b_bits_id; // @[Parameters.scala 47:9]
  wire  requestBOI_9_0 = ~auto_out_9_b_bits_id; // @[Parameters.scala 47:9]
  wire  requestBOI_10_0 = ~auto_out_10_b_bits_id; // @[Parameters.scala 47:9]
  wire  requestBOI_11_0 = ~auto_out_11_b_bits_id; // @[Parameters.scala 47:9]
  wire  requestBOI_12_0 = ~auto_out_12_b_bits_id; // @[Parameters.scala 47:9]
  wire  requestBOI_13_0 = ~auto_out_13_b_bits_id; // @[Parameters.scala 47:9]
  wire  requestBOI_14_0 = ~auto_out_14_b_bits_id; // @[Parameters.scala 47:9]
  wire  requestBOI_15_0 = ~auto_out_15_b_bits_id; // @[Parameters.scala 47:9]
  wire  requestBOI_16_0 = ~auto_out_16_b_bits_id; // @[Parameters.scala 47:9]
  wire  requestBOI_17_0 = ~auto_out_17_b_bits_id; // @[Parameters.scala 47:9]
  wire  requestBOI_18_0 = ~auto_out_18_b_bits_id; // @[Parameters.scala 47:9]
  wire  requestBOI_19_0 = ~auto_out_19_b_bits_id; // @[Parameters.scala 47:9]
  wire [9:0] _T_242 = {requestAWIO_0_9,requestAWIO_0_8,requestAWIO_0_7,requestAWIO_0_6,requestAWIO_0_5,requestAWIO_0_4,requestAWIO_0_3,requestAWIO_0_2,requestAWIO_0_1,requestAWIO_0_0}; // @[Xbar.scala 64:75]
  wire [4:0] _T_246 = {requestAWIO_0_14,requestAWIO_0_13,requestAWIO_0_12,requestAWIO_0_11,requestAWIO_0_10}; // @[Xbar.scala 64:75]
  wire [10:0] _T_252 = {requestAWIO_0_20,requestAWIO_0_19,requestAWIO_0_18,requestAWIO_0_17,requestAWIO_0_16,requestAWIO_0_15,_T_246}; // @[Xbar.scala 64:75]
  wire [20:0] _T_253 = {requestAWIO_0_20,requestAWIO_0_19,requestAWIO_0_18,requestAWIO_0_17,requestAWIO_0_16,requestAWIO_0_15,_T_246,_T_242}; // @[Xbar.scala 64:75]
  wire  requestWIO_0_0 = awIn_0_io_deq_bits[0]; // @[Xbar.scala 65:73]
  wire  requestWIO_0_1 = awIn_0_io_deq_bits[1]; // @[Xbar.scala 65:73]
  wire  requestWIO_0_2 = awIn_0_io_deq_bits[2]; // @[Xbar.scala 65:73]
  wire  requestWIO_0_3 = awIn_0_io_deq_bits[3]; // @[Xbar.scala 65:73]
  wire  requestWIO_0_4 = awIn_0_io_deq_bits[4]; // @[Xbar.scala 65:73]
  wire  requestWIO_0_5 = awIn_0_io_deq_bits[5]; // @[Xbar.scala 65:73]
  wire  requestWIO_0_6 = awIn_0_io_deq_bits[6]; // @[Xbar.scala 65:73]
  wire  requestWIO_0_7 = awIn_0_io_deq_bits[7]; // @[Xbar.scala 65:73]
  wire  requestWIO_0_8 = awIn_0_io_deq_bits[8]; // @[Xbar.scala 65:73]
  wire  requestWIO_0_9 = awIn_0_io_deq_bits[9]; // @[Xbar.scala 65:73]
  wire  requestWIO_0_10 = awIn_0_io_deq_bits[10]; // @[Xbar.scala 65:73]
  wire  requestWIO_0_11 = awIn_0_io_deq_bits[11]; // @[Xbar.scala 65:73]
  wire  requestWIO_0_12 = awIn_0_io_deq_bits[12]; // @[Xbar.scala 65:73]
  wire  requestWIO_0_13 = awIn_0_io_deq_bits[13]; // @[Xbar.scala 65:73]
  wire  requestWIO_0_14 = awIn_0_io_deq_bits[14]; // @[Xbar.scala 65:73]
  wire  requestWIO_0_15 = awIn_0_io_deq_bits[15]; // @[Xbar.scala 65:73]
  wire  requestWIO_0_16 = awIn_0_io_deq_bits[16]; // @[Xbar.scala 65:73]
  wire  requestWIO_0_17 = awIn_0_io_deq_bits[17]; // @[Xbar.scala 65:73]
  wire  requestWIO_0_18 = awIn_0_io_deq_bits[18]; // @[Xbar.scala 65:73]
  wire  requestWIO_0_19 = awIn_0_io_deq_bits[19]; // @[Xbar.scala 65:73]
  wire  requestWIO_0_20 = awIn_0_io_deq_bits[20]; // @[Xbar.scala 65:73]
  wire [9:0] _T_268 = {requestARIO_0_9,requestARIO_0_8,requestARIO_0_7,requestARIO_0_6,requestARIO_0_5,requestARIO_0_4,requestARIO_0_3,requestARIO_0_2,requestARIO_0_1,requestARIO_0_0}; // @[Xbar.scala 93:45]
  wire [4:0] _T_272 = {requestARIO_0_14,requestARIO_0_13,requestARIO_0_12,requestARIO_0_11,requestARIO_0_10}; // @[Xbar.scala 93:45]
  wire [20:0] _T_279 = {requestARIO_0_20,requestARIO_0_19,requestARIO_0_18,requestARIO_0_17,requestARIO_0_16,requestARIO_0_15,_T_272,_T_268}; // @[Xbar.scala 93:45]
  wire  _T_282 = _T_279[20:16] != 5'h0; // @[OneHot.scala 32:14]
  wire [15:0] _GEN_94 = {{11'd0}, _T_279[20:16]}; // @[OneHot.scala 32:28]
  wire [15:0] _T_283 = _GEN_94 | _T_279[15:0]; // @[OneHot.scala 32:28]
  wire  _T_286 = _T_283[15:8] != 8'h0; // @[OneHot.scala 32:14]
  wire [7:0] _T_287 = _T_283[15:8] | _T_283[7:0]; // @[OneHot.scala 32:28]
  wire  _T_290 = _T_287[7:4] != 4'h0; // @[OneHot.scala 32:14]
  wire [3:0] _T_291 = _T_287[7:4] | _T_287[3:0]; // @[OneHot.scala 32:28]
  wire  _T_294 = _T_291[3:2] != 2'h0; // @[OneHot.scala 32:14]
  wire [1:0] _T_295 = _T_291[3:2] | _T_291[1:0]; // @[OneHot.scala 32:28]
  wire [4:0] _T_300 = {_T_282,_T_286,_T_290,_T_294,_T_295[1]}; // @[Cat.scala 29:58]
  wire  _T_323 = _T_253[20:16] != 5'h0; // @[OneHot.scala 32:14]
  wire [15:0] _GEN_95 = {{11'd0}, _T_253[20:16]}; // @[OneHot.scala 32:28]
  wire [15:0] _T_324 = _GEN_95 | _T_253[15:0]; // @[OneHot.scala 32:28]
  wire  _T_327 = _T_324[15:8] != 8'h0; // @[OneHot.scala 32:14]
  wire [7:0] _T_328 = _T_324[15:8] | _T_324[7:0]; // @[OneHot.scala 32:28]
  wire  _T_331 = _T_328[7:4] != 4'h0; // @[OneHot.scala 32:14]
  wire [3:0] _T_332 = _T_328[7:4] | _T_328[3:0]; // @[OneHot.scala 32:28]
  wire  _T_335 = _T_332[3:2] != 2'h0; // @[OneHot.scala 32:14]
  wire [1:0] _T_336 = _T_332[3:2] | _T_332[1:0]; // @[OneHot.scala 32:28]
  wire [4:0] _T_341 = {_T_323,_T_327,_T_331,_T_335,_T_336[1]}; // @[Cat.scala 29:58]
  wire  _T_438 = requestARIO_0_0 & auto_out_0_ar_ready; // @[Mux.scala 27:72]
  wire  _T_439 = requestARIO_0_1 & auto_out_1_ar_ready; // @[Mux.scala 27:72]
  wire  _T_459 = _T_438 | _T_439; // @[Mux.scala 27:72]
  wire  _T_440 = requestARIO_0_2 & auto_out_2_ar_ready; // @[Mux.scala 27:72]
  wire  _T_460 = _T_459 | _T_440; // @[Mux.scala 27:72]
  wire  _T_441 = requestARIO_0_3 & auto_out_3_ar_ready; // @[Mux.scala 27:72]
  wire  _T_461 = _T_460 | _T_441; // @[Mux.scala 27:72]
  wire  _T_442 = requestARIO_0_4 & auto_out_4_ar_ready; // @[Mux.scala 27:72]
  wire  _T_462 = _T_461 | _T_442; // @[Mux.scala 27:72]
  wire  _T_443 = requestARIO_0_5 & auto_out_5_ar_ready; // @[Mux.scala 27:72]
  wire  _T_463 = _T_462 | _T_443; // @[Mux.scala 27:72]
  wire  _T_444 = requestARIO_0_6 & auto_out_6_ar_ready; // @[Mux.scala 27:72]
  wire  _T_464 = _T_463 | _T_444; // @[Mux.scala 27:72]
  wire  _T_445 = requestARIO_0_7 & auto_out_7_ar_ready; // @[Mux.scala 27:72]
  wire  _T_465 = _T_464 | _T_445; // @[Mux.scala 27:72]
  wire  _T_446 = requestARIO_0_8 & auto_out_8_ar_ready; // @[Mux.scala 27:72]
  wire  _T_466 = _T_465 | _T_446; // @[Mux.scala 27:72]
  wire  _T_447 = requestARIO_0_9 & auto_out_9_ar_ready; // @[Mux.scala 27:72]
  wire  _T_467 = _T_466 | _T_447; // @[Mux.scala 27:72]
  wire  _T_448 = requestARIO_0_10 & auto_out_10_ar_ready; // @[Mux.scala 27:72]
  wire  _T_468 = _T_467 | _T_448; // @[Mux.scala 27:72]
  wire  _T_449 = requestARIO_0_11 & auto_out_11_ar_ready; // @[Mux.scala 27:72]
  wire  _T_469 = _T_468 | _T_449; // @[Mux.scala 27:72]
  wire  _T_450 = requestARIO_0_12 & auto_out_12_ar_ready; // @[Mux.scala 27:72]
  wire  _T_470 = _T_469 | _T_450; // @[Mux.scala 27:72]
  wire  _T_451 = requestARIO_0_13 & auto_out_13_ar_ready; // @[Mux.scala 27:72]
  wire  _T_471 = _T_470 | _T_451; // @[Mux.scala 27:72]
  wire  _T_452 = requestARIO_0_14 & auto_out_14_ar_ready; // @[Mux.scala 27:72]
  wire  _T_472 = _T_471 | _T_452; // @[Mux.scala 27:72]
  wire  _T_453 = requestARIO_0_15 & auto_out_15_ar_ready; // @[Mux.scala 27:72]
  wire  _T_473 = _T_472 | _T_453; // @[Mux.scala 27:72]
  wire  _T_454 = requestARIO_0_16 & auto_out_16_ar_ready; // @[Mux.scala 27:72]
  wire  _T_474 = _T_473 | _T_454; // @[Mux.scala 27:72]
  wire  _T_455 = requestARIO_0_17 & auto_out_17_ar_ready; // @[Mux.scala 27:72]
  wire  _T_475 = _T_474 | _T_455; // @[Mux.scala 27:72]
  wire  _T_456 = requestARIO_0_18 & auto_out_18_ar_ready; // @[Mux.scala 27:72]
  wire  _T_476 = _T_475 | _T_456; // @[Mux.scala 27:72]
  wire  _T_457 = requestARIO_0_19 & auto_out_19_ar_ready; // @[Mux.scala 27:72]
  wire  _T_477 = _T_476 | _T_457; // @[Mux.scala 27:72]
  wire  _T_458 = requestARIO_0_20 & auto_out_20_ar_ready; // @[Mux.scala 27:72]
  wire  in_0_ar_ready = _T_477 | _T_458; // @[Mux.scala 27:72]
  reg [2:0] _T_347; // @[Xbar.scala 104:34]
  reg [31:0] _RAND_0;
  wire  _T_366 = _T_347 == 3'h0; // @[Xbar.scala 112:22]
  reg [4:0] _T_348; // @[Xbar.scala 105:29]
  reg [31:0] _RAND_1;
  wire  _T_365 = _T_348 == _T_300; // @[Xbar.scala 111:75]
  wire  _T_367 = _T_366 | _T_365; // @[Xbar.scala 112:34]
  wire  _T_368 = _T_347 != 3'h7; // @[Xbar.scala 112:80]
  wire  _T_370 = _T_367 & _T_368; // @[Xbar.scala 112:48]
  wire  io_in_0_ar_ready = in_0_ar_ready & _T_370; // @[Xbar.scala 130:45]
  wire  _T_342 = io_in_0_ar_ready & auto_in_ar_valid; // @[Decoupled.scala 40:37]
  reg  _T_1616; // @[Xbar.scala 242:23]
  reg [31:0] _RAND_2;
  wire  _T_609 = auto_out_0_r_valid & requestROI_0_0; // @[Xbar.scala 222:40]
  wire  _T_611 = auto_out_1_r_valid & requestROI_1_0; // @[Xbar.scala 222:40]
  wire  _T_1617 = _T_609 | _T_611; // @[Xbar.scala 246:36]
  wire  _T_613 = auto_out_2_r_valid & requestROI_2_0; // @[Xbar.scala 222:40]
  wire  _T_1618 = _T_1617 | _T_613; // @[Xbar.scala 246:36]
  wire  _T_615 = auto_out_3_r_valid & requestROI_3_0; // @[Xbar.scala 222:40]
  wire  _T_1619 = _T_1618 | _T_615; // @[Xbar.scala 246:36]
  wire  _T_617 = auto_out_4_r_valid & requestROI_4_0; // @[Xbar.scala 222:40]
  wire  _T_1620 = _T_1619 | _T_617; // @[Xbar.scala 246:36]
  wire  _T_619 = auto_out_5_r_valid & requestROI_5_0; // @[Xbar.scala 222:40]
  wire  _T_1621 = _T_1620 | _T_619; // @[Xbar.scala 246:36]
  wire  _T_621 = auto_out_6_r_valid & requestROI_6_0; // @[Xbar.scala 222:40]
  wire  _T_1622 = _T_1621 | _T_621; // @[Xbar.scala 246:36]
  wire  _T_623 = auto_out_7_r_valid & requestROI_7_0; // @[Xbar.scala 222:40]
  wire  _T_1623 = _T_1622 | _T_623; // @[Xbar.scala 246:36]
  wire  _T_625 = auto_out_8_r_valid & requestROI_8_0; // @[Xbar.scala 222:40]
  wire  _T_1624 = _T_1623 | _T_625; // @[Xbar.scala 246:36]
  wire  _T_627 = auto_out_9_r_valid & requestROI_9_0; // @[Xbar.scala 222:40]
  wire  _T_1625 = _T_1624 | _T_627; // @[Xbar.scala 246:36]
  wire  _T_629 = auto_out_10_r_valid & requestROI_10_0; // @[Xbar.scala 222:40]
  wire  _T_1626 = _T_1625 | _T_629; // @[Xbar.scala 246:36]
  wire  _T_631 = auto_out_11_r_valid & requestROI_11_0; // @[Xbar.scala 222:40]
  wire  _T_1627 = _T_1626 | _T_631; // @[Xbar.scala 246:36]
  wire  _T_633 = auto_out_12_r_valid & requestROI_12_0; // @[Xbar.scala 222:40]
  wire  _T_1628 = _T_1627 | _T_633; // @[Xbar.scala 246:36]
  wire  _T_635 = auto_out_13_r_valid & requestROI_13_0; // @[Xbar.scala 222:40]
  wire  _T_1629 = _T_1628 | _T_635; // @[Xbar.scala 246:36]
  wire  _T_637 = auto_out_14_r_valid & requestROI_14_0; // @[Xbar.scala 222:40]
  wire  _T_1630 = _T_1629 | _T_637; // @[Xbar.scala 246:36]
  wire  _T_639 = auto_out_15_r_valid & requestROI_15_0; // @[Xbar.scala 222:40]
  wire  _T_1631 = _T_1630 | _T_639; // @[Xbar.scala 246:36]
  wire  _T_641 = auto_out_16_r_valid & requestROI_16_0; // @[Xbar.scala 222:40]
  wire  _T_1632 = _T_1631 | _T_641; // @[Xbar.scala 246:36]
  wire  _T_643 = auto_out_17_r_valid & requestROI_17_0; // @[Xbar.scala 222:40]
  wire  _T_1633 = _T_1632 | _T_643; // @[Xbar.scala 246:36]
  wire  _T_645 = auto_out_18_r_valid & requestROI_18_0; // @[Xbar.scala 222:40]
  wire  _T_1634 = _T_1633 | _T_645; // @[Xbar.scala 246:36]
  wire  _T_647 = auto_out_19_r_valid & requestROI_19_0; // @[Xbar.scala 222:40]
  wire  _T_1635 = _T_1634 | _T_647; // @[Xbar.scala 246:36]
  wire  _T_1636 = _T_1635 | auto_out_20_r_valid; // @[Xbar.scala 246:36]
  reg  _T_1882_0; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_3;
  wire  _T_1907 = _T_1882_0 & _T_609; // @[Mux.scala 27:72]
  reg  _T_1882_1; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_4;
  wire  _T_1908 = _T_1882_1 & _T_611; // @[Mux.scala 27:72]
  wire  _T_1928 = _T_1907 | _T_1908; // @[Mux.scala 27:72]
  reg  _T_1882_2; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_5;
  wire  _T_1909 = _T_1882_2 & _T_613; // @[Mux.scala 27:72]
  wire  _T_1929 = _T_1928 | _T_1909; // @[Mux.scala 27:72]
  reg  _T_1882_3; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_6;
  wire  _T_1910 = _T_1882_3 & _T_615; // @[Mux.scala 27:72]
  wire  _T_1930 = _T_1929 | _T_1910; // @[Mux.scala 27:72]
  reg  _T_1882_4; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_7;
  wire  _T_1911 = _T_1882_4 & _T_617; // @[Mux.scala 27:72]
  wire  _T_1931 = _T_1930 | _T_1911; // @[Mux.scala 27:72]
  reg  _T_1882_5; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_8;
  wire  _T_1912 = _T_1882_5 & _T_619; // @[Mux.scala 27:72]
  wire  _T_1932 = _T_1931 | _T_1912; // @[Mux.scala 27:72]
  reg  _T_1882_6; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_9;
  wire  _T_1913 = _T_1882_6 & _T_621; // @[Mux.scala 27:72]
  wire  _T_1933 = _T_1932 | _T_1913; // @[Mux.scala 27:72]
  reg  _T_1882_7; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_10;
  wire  _T_1914 = _T_1882_7 & _T_623; // @[Mux.scala 27:72]
  wire  _T_1934 = _T_1933 | _T_1914; // @[Mux.scala 27:72]
  reg  _T_1882_8; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_11;
  wire  _T_1915 = _T_1882_8 & _T_625; // @[Mux.scala 27:72]
  wire  _T_1935 = _T_1934 | _T_1915; // @[Mux.scala 27:72]
  reg  _T_1882_9; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_12;
  wire  _T_1916 = _T_1882_9 & _T_627; // @[Mux.scala 27:72]
  wire  _T_1936 = _T_1935 | _T_1916; // @[Mux.scala 27:72]
  reg  _T_1882_10; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_13;
  wire  _T_1917 = _T_1882_10 & _T_629; // @[Mux.scala 27:72]
  wire  _T_1937 = _T_1936 | _T_1917; // @[Mux.scala 27:72]
  reg  _T_1882_11; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_14;
  wire  _T_1918 = _T_1882_11 & _T_631; // @[Mux.scala 27:72]
  wire  _T_1938 = _T_1937 | _T_1918; // @[Mux.scala 27:72]
  reg  _T_1882_12; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_15;
  wire  _T_1919 = _T_1882_12 & _T_633; // @[Mux.scala 27:72]
  wire  _T_1939 = _T_1938 | _T_1919; // @[Mux.scala 27:72]
  reg  _T_1882_13; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_16;
  wire  _T_1920 = _T_1882_13 & _T_635; // @[Mux.scala 27:72]
  wire  _T_1940 = _T_1939 | _T_1920; // @[Mux.scala 27:72]
  reg  _T_1882_14; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_17;
  wire  _T_1921 = _T_1882_14 & _T_637; // @[Mux.scala 27:72]
  wire  _T_1941 = _T_1940 | _T_1921; // @[Mux.scala 27:72]
  reg  _T_1882_15; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_18;
  wire  _T_1922 = _T_1882_15 & _T_639; // @[Mux.scala 27:72]
  wire  _T_1942 = _T_1941 | _T_1922; // @[Mux.scala 27:72]
  reg  _T_1882_16; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_19;
  wire  _T_1923 = _T_1882_16 & _T_641; // @[Mux.scala 27:72]
  wire  _T_1943 = _T_1942 | _T_1923; // @[Mux.scala 27:72]
  reg  _T_1882_17; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_20;
  wire  _T_1924 = _T_1882_17 & _T_643; // @[Mux.scala 27:72]
  wire  _T_1944 = _T_1943 | _T_1924; // @[Mux.scala 27:72]
  reg  _T_1882_18; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_21;
  wire  _T_1925 = _T_1882_18 & _T_645; // @[Mux.scala 27:72]
  wire  _T_1945 = _T_1944 | _T_1925; // @[Mux.scala 27:72]
  reg  _T_1882_19; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_22;
  wire  _T_1926 = _T_1882_19 & _T_647; // @[Mux.scala 27:72]
  wire  _T_1946 = _T_1945 | _T_1926; // @[Mux.scala 27:72]
  reg  _T_1882_20; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_23;
  wire  _T_1927 = _T_1882_20 & auto_out_20_r_valid; // @[Mux.scala 27:72]
  wire  _T_1947 = _T_1946 | _T_1927; // @[Mux.scala 27:72]
  wire  in_0_r_valid = _T_1616 ? _T_1636 : _T_1947; // @[Xbar.scala 278:22]
  wire  _T_344 = auto_in_r_ready & in_0_r_valid; // @[Decoupled.scala 40:37]
  wire [4:0] _T_1649 = {_T_637,_T_635,_T_633,_T_631,_T_629}; // @[Cat.scala 29:58]
  wire [9:0] _T_1645 = {_T_627,_T_625,_T_623,_T_621,_T_619,_T_617,_T_615,_T_613,_T_611,_T_609}; // @[Cat.scala 29:58]
  wire [20:0] _T_1656 = {auto_out_20_r_valid,_T_647,_T_645,_T_643,_T_641,_T_639,_T_1649,_T_1645}; // @[Cat.scala 29:58]
  reg [20:0] _T_1663; // @[Arbiter.scala 20:23]
  reg [31:0] _RAND_24;
  wire [20:0] _T_1664 = ~_T_1663; // @[Arbiter.scala 21:30]
  wire [20:0] _T_1665 = _T_1656 & _T_1664; // @[Arbiter.scala 21:28]
  wire [41:0] _T_1666 = {_T_1665,auto_out_20_r_valid,_T_647,_T_645,_T_643,_T_641,_T_639,_T_1649,_T_1645}; // @[Cat.scala 29:58]
  wire [41:0] _GEN_96 = {{1'd0}, _T_1666[41:1]}; // @[package.scala 208:43]
  wire [41:0] _T_1668 = _T_1666 | _GEN_96; // @[package.scala 208:43]
  wire [41:0] _GEN_97 = {{2'd0}, _T_1668[41:2]}; // @[package.scala 208:43]
  wire [41:0] _T_1670 = _T_1668 | _GEN_97; // @[package.scala 208:43]
  wire [41:0] _GEN_98 = {{4'd0}, _T_1670[41:4]}; // @[package.scala 208:43]
  wire [41:0] _T_1672 = _T_1670 | _GEN_98; // @[package.scala 208:43]
  wire [41:0] _GEN_99 = {{8'd0}, _T_1672[41:8]}; // @[package.scala 208:43]
  wire [41:0] _T_1674 = _T_1672 | _GEN_99; // @[package.scala 208:43]
  wire [41:0] _GEN_100 = {{16'd0}, _T_1674[41:16]}; // @[package.scala 208:43]
  wire [41:0] _T_1676 = _T_1674 | _GEN_100; // @[package.scala 208:43]
  wire [41:0] _T_1679 = {_T_1663, 21'h0}; // @[Arbiter.scala 22:66]
  wire [41:0] _GEN_101 = {{1'd0}, _T_1676[41:1]}; // @[Arbiter.scala 22:58]
  wire [41:0] _T_1680 = _GEN_101 | _T_1679; // @[Arbiter.scala 22:58]
  wire [20:0] _T_1683 = _T_1680[41:21] & _T_1680[20:0]; // @[Arbiter.scala 23:39]
  wire [20:0] _T_1684 = ~_T_1683; // @[Arbiter.scala 23:18]
  wire  _T_1727 = _T_1684[0] & _T_609; // @[Xbar.scala 250:63]
  wire  _T_1883_0 = _T_1616 ? _T_1727 : _T_1882_0; // @[Xbar.scala 262:23]
  wire [35:0] _T_1952 = {auto_out_0_r_bits_id,auto_out_0_r_bits_data,auto_out_0_r_bits_resp,auto_out_0_r_bits_last}; // @[Mux.scala 27:72]
  wire [35:0] _T_1953 = _T_1883_0 ? _T_1952 : 36'h0; // @[Mux.scala 27:72]
  wire  _T_1728 = _T_1684[1] & _T_611; // @[Xbar.scala 250:63]
  wire  _T_1883_1 = _T_1616 ? _T_1728 : _T_1882_1; // @[Xbar.scala 262:23]
  wire [35:0] _T_1956 = {auto_out_1_r_bits_id,auto_out_1_r_bits_data,auto_out_1_r_bits_resp,auto_out_1_r_bits_last}; // @[Mux.scala 27:72]
  wire [35:0] _T_1957 = _T_1883_1 ? _T_1956 : 36'h0; // @[Mux.scala 27:72]
  wire [35:0] _T_2034 = _T_1953 | _T_1957; // @[Mux.scala 27:72]
  wire  _T_1729 = _T_1684[2] & _T_613; // @[Xbar.scala 250:63]
  wire  _T_1883_2 = _T_1616 ? _T_1729 : _T_1882_2; // @[Xbar.scala 262:23]
  wire [35:0] _T_1960 = {auto_out_2_r_bits_id,auto_out_2_r_bits_data,auto_out_2_r_bits_resp,auto_out_2_r_bits_last}; // @[Mux.scala 27:72]
  wire [35:0] _T_1961 = _T_1883_2 ? _T_1960 : 36'h0; // @[Mux.scala 27:72]
  wire [35:0] _T_2035 = _T_2034 | _T_1961; // @[Mux.scala 27:72]
  wire  _T_1730 = _T_1684[3] & _T_615; // @[Xbar.scala 250:63]
  wire  _T_1883_3 = _T_1616 ? _T_1730 : _T_1882_3; // @[Xbar.scala 262:23]
  wire [35:0] _T_1964 = {auto_out_3_r_bits_id,auto_out_3_r_bits_data,auto_out_3_r_bits_resp,auto_out_3_r_bits_last}; // @[Mux.scala 27:72]
  wire [35:0] _T_1965 = _T_1883_3 ? _T_1964 : 36'h0; // @[Mux.scala 27:72]
  wire [35:0] _T_2036 = _T_2035 | _T_1965; // @[Mux.scala 27:72]
  wire  _T_1731 = _T_1684[4] & _T_617; // @[Xbar.scala 250:63]
  wire  _T_1883_4 = _T_1616 ? _T_1731 : _T_1882_4; // @[Xbar.scala 262:23]
  wire [35:0] _T_1968 = {auto_out_4_r_bits_id,auto_out_4_r_bits_data,auto_out_4_r_bits_resp,auto_out_4_r_bits_last}; // @[Mux.scala 27:72]
  wire [35:0] _T_1969 = _T_1883_4 ? _T_1968 : 36'h0; // @[Mux.scala 27:72]
  wire [35:0] _T_2037 = _T_2036 | _T_1969; // @[Mux.scala 27:72]
  wire  _T_1732 = _T_1684[5] & _T_619; // @[Xbar.scala 250:63]
  wire  _T_1883_5 = _T_1616 ? _T_1732 : _T_1882_5; // @[Xbar.scala 262:23]
  wire [35:0] _T_1972 = {auto_out_5_r_bits_id,auto_out_5_r_bits_data,auto_out_5_r_bits_resp,auto_out_5_r_bits_last}; // @[Mux.scala 27:72]
  wire [35:0] _T_1973 = _T_1883_5 ? _T_1972 : 36'h0; // @[Mux.scala 27:72]
  wire [35:0] _T_2038 = _T_2037 | _T_1973; // @[Mux.scala 27:72]
  wire  _T_1733 = _T_1684[6] & _T_621; // @[Xbar.scala 250:63]
  wire  _T_1883_6 = _T_1616 ? _T_1733 : _T_1882_6; // @[Xbar.scala 262:23]
  wire [35:0] _T_1976 = {auto_out_6_r_bits_id,auto_out_6_r_bits_data,auto_out_6_r_bits_resp,auto_out_6_r_bits_last}; // @[Mux.scala 27:72]
  wire [35:0] _T_1977 = _T_1883_6 ? _T_1976 : 36'h0; // @[Mux.scala 27:72]
  wire [35:0] _T_2039 = _T_2038 | _T_1977; // @[Mux.scala 27:72]
  wire  _T_1734 = _T_1684[7] & _T_623; // @[Xbar.scala 250:63]
  wire  _T_1883_7 = _T_1616 ? _T_1734 : _T_1882_7; // @[Xbar.scala 262:23]
  wire [35:0] _T_1980 = {auto_out_7_r_bits_id,auto_out_7_r_bits_data,auto_out_7_r_bits_resp,auto_out_7_r_bits_last}; // @[Mux.scala 27:72]
  wire [35:0] _T_1981 = _T_1883_7 ? _T_1980 : 36'h0; // @[Mux.scala 27:72]
  wire [35:0] _T_2040 = _T_2039 | _T_1981; // @[Mux.scala 27:72]
  wire  _T_1735 = _T_1684[8] & _T_625; // @[Xbar.scala 250:63]
  wire  _T_1883_8 = _T_1616 ? _T_1735 : _T_1882_8; // @[Xbar.scala 262:23]
  wire [35:0] _T_1984 = {auto_out_8_r_bits_id,auto_out_8_r_bits_data,auto_out_8_r_bits_resp,auto_out_8_r_bits_last}; // @[Mux.scala 27:72]
  wire [35:0] _T_1985 = _T_1883_8 ? _T_1984 : 36'h0; // @[Mux.scala 27:72]
  wire [35:0] _T_2041 = _T_2040 | _T_1985; // @[Mux.scala 27:72]
  wire  _T_1736 = _T_1684[9] & _T_627; // @[Xbar.scala 250:63]
  wire  _T_1883_9 = _T_1616 ? _T_1736 : _T_1882_9; // @[Xbar.scala 262:23]
  wire [35:0] _T_1988 = {auto_out_9_r_bits_id,auto_out_9_r_bits_data,auto_out_9_r_bits_resp,auto_out_9_r_bits_last}; // @[Mux.scala 27:72]
  wire [35:0] _T_1989 = _T_1883_9 ? _T_1988 : 36'h0; // @[Mux.scala 27:72]
  wire [35:0] _T_2042 = _T_2041 | _T_1989; // @[Mux.scala 27:72]
  wire  _T_1737 = _T_1684[10] & _T_629; // @[Xbar.scala 250:63]
  wire  _T_1883_10 = _T_1616 ? _T_1737 : _T_1882_10; // @[Xbar.scala 262:23]
  wire [35:0] _T_1992 = {auto_out_10_r_bits_id,auto_out_10_r_bits_data,auto_out_10_r_bits_resp,auto_out_10_r_bits_last}; // @[Mux.scala 27:72]
  wire [35:0] _T_1993 = _T_1883_10 ? _T_1992 : 36'h0; // @[Mux.scala 27:72]
  wire [35:0] _T_2043 = _T_2042 | _T_1993; // @[Mux.scala 27:72]
  wire  _T_1738 = _T_1684[11] & _T_631; // @[Xbar.scala 250:63]
  wire  _T_1883_11 = _T_1616 ? _T_1738 : _T_1882_11; // @[Xbar.scala 262:23]
  wire [35:0] _T_1996 = {auto_out_11_r_bits_id,auto_out_11_r_bits_data,auto_out_11_r_bits_resp,auto_out_11_r_bits_last}; // @[Mux.scala 27:72]
  wire [35:0] _T_1997 = _T_1883_11 ? _T_1996 : 36'h0; // @[Mux.scala 27:72]
  wire [35:0] _T_2044 = _T_2043 | _T_1997; // @[Mux.scala 27:72]
  wire  _T_1739 = _T_1684[12] & _T_633; // @[Xbar.scala 250:63]
  wire  _T_1883_12 = _T_1616 ? _T_1739 : _T_1882_12; // @[Xbar.scala 262:23]
  wire [35:0] _T_2000 = {auto_out_12_r_bits_id,auto_out_12_r_bits_data,auto_out_12_r_bits_resp,auto_out_12_r_bits_last}; // @[Mux.scala 27:72]
  wire [35:0] _T_2001 = _T_1883_12 ? _T_2000 : 36'h0; // @[Mux.scala 27:72]
  wire [35:0] _T_2045 = _T_2044 | _T_2001; // @[Mux.scala 27:72]
  wire  _T_1740 = _T_1684[13] & _T_635; // @[Xbar.scala 250:63]
  wire  _T_1883_13 = _T_1616 ? _T_1740 : _T_1882_13; // @[Xbar.scala 262:23]
  wire [35:0] _T_2004 = {auto_out_13_r_bits_id,auto_out_13_r_bits_data,auto_out_13_r_bits_resp,auto_out_13_r_bits_last}; // @[Mux.scala 27:72]
  wire [35:0] _T_2005 = _T_1883_13 ? _T_2004 : 36'h0; // @[Mux.scala 27:72]
  wire [35:0] _T_2046 = _T_2045 | _T_2005; // @[Mux.scala 27:72]
  wire  _T_1741 = _T_1684[14] & _T_637; // @[Xbar.scala 250:63]
  wire  _T_1883_14 = _T_1616 ? _T_1741 : _T_1882_14; // @[Xbar.scala 262:23]
  wire [35:0] _T_2008 = {auto_out_14_r_bits_id,auto_out_14_r_bits_data,auto_out_14_r_bits_resp,auto_out_14_r_bits_last}; // @[Mux.scala 27:72]
  wire [35:0] _T_2009 = _T_1883_14 ? _T_2008 : 36'h0; // @[Mux.scala 27:72]
  wire [35:0] _T_2047 = _T_2046 | _T_2009; // @[Mux.scala 27:72]
  wire  _T_1742 = _T_1684[15] & _T_639; // @[Xbar.scala 250:63]
  wire  _T_1883_15 = _T_1616 ? _T_1742 : _T_1882_15; // @[Xbar.scala 262:23]
  wire [35:0] _T_2012 = {auto_out_15_r_bits_id,auto_out_15_r_bits_data,auto_out_15_r_bits_resp,auto_out_15_r_bits_last}; // @[Mux.scala 27:72]
  wire [35:0] _T_2013 = _T_1883_15 ? _T_2012 : 36'h0; // @[Mux.scala 27:72]
  wire [35:0] _T_2048 = _T_2047 | _T_2013; // @[Mux.scala 27:72]
  wire  _T_1743 = _T_1684[16] & _T_641; // @[Xbar.scala 250:63]
  wire  _T_1883_16 = _T_1616 ? _T_1743 : _T_1882_16; // @[Xbar.scala 262:23]
  wire [35:0] _T_2016 = {auto_out_16_r_bits_id,auto_out_16_r_bits_data,auto_out_16_r_bits_resp,auto_out_16_r_bits_last}; // @[Mux.scala 27:72]
  wire [35:0] _T_2017 = _T_1883_16 ? _T_2016 : 36'h0; // @[Mux.scala 27:72]
  wire [35:0] _T_2049 = _T_2048 | _T_2017; // @[Mux.scala 27:72]
  wire  _T_1744 = _T_1684[17] & _T_643; // @[Xbar.scala 250:63]
  wire  _T_1883_17 = _T_1616 ? _T_1744 : _T_1882_17; // @[Xbar.scala 262:23]
  wire [35:0] _T_2020 = {auto_out_17_r_bits_id,auto_out_17_r_bits_data,auto_out_17_r_bits_resp,auto_out_17_r_bits_last}; // @[Mux.scala 27:72]
  wire [35:0] _T_2021 = _T_1883_17 ? _T_2020 : 36'h0; // @[Mux.scala 27:72]
  wire [35:0] _T_2050 = _T_2049 | _T_2021; // @[Mux.scala 27:72]
  wire  _T_1745 = _T_1684[18] & _T_645; // @[Xbar.scala 250:63]
  wire  _T_1883_18 = _T_1616 ? _T_1745 : _T_1882_18; // @[Xbar.scala 262:23]
  wire [35:0] _T_2024 = {auto_out_18_r_bits_id,auto_out_18_r_bits_data,auto_out_18_r_bits_resp,auto_out_18_r_bits_last}; // @[Mux.scala 27:72]
  wire [35:0] _T_2025 = _T_1883_18 ? _T_2024 : 36'h0; // @[Mux.scala 27:72]
  wire [35:0] _T_2051 = _T_2050 | _T_2025; // @[Mux.scala 27:72]
  wire  _T_1746 = _T_1684[19] & _T_647; // @[Xbar.scala 250:63]
  wire  _T_1883_19 = _T_1616 ? _T_1746 : _T_1882_19; // @[Xbar.scala 262:23]
  wire [35:0] _T_2028 = {auto_out_19_r_bits_id,auto_out_19_r_bits_data,auto_out_19_r_bits_resp,auto_out_19_r_bits_last}; // @[Mux.scala 27:72]
  wire [35:0] _T_2029 = _T_1883_19 ? _T_2028 : 36'h0; // @[Mux.scala 27:72]
  wire [35:0] _T_2052 = _T_2051 | _T_2029; // @[Mux.scala 27:72]
  wire  _T_1747 = _T_1684[20] & auto_out_20_r_valid; // @[Xbar.scala 250:63]
  wire  _T_1883_20 = _T_1616 ? _T_1747 : _T_1882_20; // @[Xbar.scala 262:23]
  wire [35:0] _T_2032 = {1'h0,auto_out_20_r_bits_data,auto_out_20_r_bits_resp,auto_out_20_r_bits_last}; // @[Mux.scala 27:72]
  wire [35:0] _T_2033 = _T_1883_20 ? _T_2032 : 36'h0; // @[Mux.scala 27:72]
  wire [35:0] _T_2053 = _T_2052 | _T_2033; // @[Mux.scala 27:72]
  wire  in_0_r_bits_last = _T_2053[0]; // @[Mux.scala 27:72]
  wire  _T_346 = _T_344 & in_0_r_bits_last; // @[Xbar.scala 120:45]
  wire [2:0] _GEN_102 = {{2'd0}, _T_342}; // @[Xbar.scala 106:30]
  wire [2:0] _T_350 = _T_347 + _GEN_102; // @[Xbar.scala 106:30]
  wire [2:0] _GEN_103 = {{2'd0}, _T_346}; // @[Xbar.scala 106:48]
  wire [2:0] _T_352 = _T_350 - _GEN_103; // @[Xbar.scala 106:48]
  wire  _T_353 = ~_T_346; // @[Xbar.scala 107:23]
  wire  _T_354 = _T_347 != 3'h0; // @[Xbar.scala 107:43]
  wire  _T_355 = _T_353 | _T_354; // @[Xbar.scala 107:34]
  wire  _T_357 = _T_355 | reset; // @[Xbar.scala 107:22]
  wire  _T_358 = ~_T_357; // @[Xbar.scala 107:22]
  wire  _T_359 = ~_T_342; // @[Xbar.scala 108:23]
  wire  _T_361 = _T_359 | _T_368; // @[Xbar.scala 108:34]
  wire  _T_363 = _T_361 | reset; // @[Xbar.scala 108:22]
  wire  _T_364 = ~_T_363; // @[Xbar.scala 108:22]
  wire  _T_502 = requestAWIO_0_0 & auto_out_0_aw_ready; // @[Mux.scala 27:72]
  wire  _T_503 = requestAWIO_0_1 & auto_out_1_aw_ready; // @[Mux.scala 27:72]
  wire  _T_523 = _T_502 | _T_503; // @[Mux.scala 27:72]
  wire  _T_504 = requestAWIO_0_2 & auto_out_2_aw_ready; // @[Mux.scala 27:72]
  wire  _T_524 = _T_523 | _T_504; // @[Mux.scala 27:72]
  wire  _T_505 = requestAWIO_0_3 & auto_out_3_aw_ready; // @[Mux.scala 27:72]
  wire  _T_525 = _T_524 | _T_505; // @[Mux.scala 27:72]
  wire  _T_506 = requestAWIO_0_4 & auto_out_4_aw_ready; // @[Mux.scala 27:72]
  wire  _T_526 = _T_525 | _T_506; // @[Mux.scala 27:72]
  wire  _T_507 = requestAWIO_0_5 & auto_out_5_aw_ready; // @[Mux.scala 27:72]
  wire  _T_527 = _T_526 | _T_507; // @[Mux.scala 27:72]
  wire  _T_508 = requestAWIO_0_6 & auto_out_6_aw_ready; // @[Mux.scala 27:72]
  wire  _T_528 = _T_527 | _T_508; // @[Mux.scala 27:72]
  wire  _T_509 = requestAWIO_0_7 & auto_out_7_aw_ready; // @[Mux.scala 27:72]
  wire  _T_529 = _T_528 | _T_509; // @[Mux.scala 27:72]
  wire  _T_510 = requestAWIO_0_8 & auto_out_8_aw_ready; // @[Mux.scala 27:72]
  wire  _T_530 = _T_529 | _T_510; // @[Mux.scala 27:72]
  wire  _T_511 = requestAWIO_0_9 & auto_out_9_aw_ready; // @[Mux.scala 27:72]
  wire  _T_531 = _T_530 | _T_511; // @[Mux.scala 27:72]
  wire  _T_512 = requestAWIO_0_10 & auto_out_10_aw_ready; // @[Mux.scala 27:72]
  wire  _T_532 = _T_531 | _T_512; // @[Mux.scala 27:72]
  wire  _T_513 = requestAWIO_0_11 & auto_out_11_aw_ready; // @[Mux.scala 27:72]
  wire  _T_533 = _T_532 | _T_513; // @[Mux.scala 27:72]
  wire  _T_514 = requestAWIO_0_12 & auto_out_12_aw_ready; // @[Mux.scala 27:72]
  wire  _T_534 = _T_533 | _T_514; // @[Mux.scala 27:72]
  wire  _T_515 = requestAWIO_0_13 & auto_out_13_aw_ready; // @[Mux.scala 27:72]
  wire  _T_535 = _T_534 | _T_515; // @[Mux.scala 27:72]
  wire  _T_516 = requestAWIO_0_14 & auto_out_14_aw_ready; // @[Mux.scala 27:72]
  wire  _T_536 = _T_535 | _T_516; // @[Mux.scala 27:72]
  wire  _T_517 = requestAWIO_0_15 & auto_out_15_aw_ready; // @[Mux.scala 27:72]
  wire  _T_537 = _T_536 | _T_517; // @[Mux.scala 27:72]
  wire  _T_518 = requestAWIO_0_16 & auto_out_16_aw_ready; // @[Mux.scala 27:72]
  wire  _T_538 = _T_537 | _T_518; // @[Mux.scala 27:72]
  wire  _T_519 = requestAWIO_0_17 & auto_out_17_aw_ready; // @[Mux.scala 27:72]
  wire  _T_539 = _T_538 | _T_519; // @[Mux.scala 27:72]
  wire  _T_520 = requestAWIO_0_18 & auto_out_18_aw_ready; // @[Mux.scala 27:72]
  wire  _T_540 = _T_539 | _T_520; // @[Mux.scala 27:72]
  wire  _T_521 = requestAWIO_0_19 & auto_out_19_aw_ready; // @[Mux.scala 27:72]
  wire  _T_541 = _T_540 | _T_521; // @[Mux.scala 27:72]
  wire  _T_522 = requestAWIO_0_20 & auto_out_20_aw_ready; // @[Mux.scala 27:72]
  wire  in_0_aw_ready = _T_541 | _T_522; // @[Mux.scala 27:72]
  reg  _T_401; // @[Xbar.scala 137:30]
  reg [31:0] _RAND_25;
  wire  _T_405 = _T_401 | awIn_0_io_enq_ready; // @[Xbar.scala 139:57]
  wire  _T_406 = in_0_aw_ready & _T_405; // @[Xbar.scala 139:45]
  reg [2:0] _T_375; // @[Xbar.scala 104:34]
  reg [31:0] _RAND_26;
  wire  _T_394 = _T_375 == 3'h0; // @[Xbar.scala 112:22]
  reg [4:0] _T_376; // @[Xbar.scala 105:29]
  reg [31:0] _RAND_27;
  wire  _T_393 = _T_376 == _T_341; // @[Xbar.scala 111:75]
  wire  _T_395 = _T_394 | _T_393; // @[Xbar.scala 112:34]
  wire  _T_396 = _T_375 != 3'h7; // @[Xbar.scala 112:80]
  wire  _T_398 = _T_395 & _T_396; // @[Xbar.scala 112:48]
  wire  io_in_0_aw_ready = _T_406 & _T_398; // @[Xbar.scala 139:82]
  wire  _T_371 = io_in_0_aw_ready & auto_in_aw_valid; // @[Decoupled.scala 40:37]
  reg  _T_2060; // @[Xbar.scala 242:23]
  reg [31:0] _RAND_28;
  wire  _T_651 = auto_out_0_b_valid & requestBOI_0_0; // @[Xbar.scala 222:40]
  wire  _T_653 = auto_out_1_b_valid & requestBOI_1_0; // @[Xbar.scala 222:40]
  wire  _T_2061 = _T_651 | _T_653; // @[Xbar.scala 246:36]
  wire  _T_655 = auto_out_2_b_valid & requestBOI_2_0; // @[Xbar.scala 222:40]
  wire  _T_2062 = _T_2061 | _T_655; // @[Xbar.scala 246:36]
  wire  _T_657 = auto_out_3_b_valid & requestBOI_3_0; // @[Xbar.scala 222:40]
  wire  _T_2063 = _T_2062 | _T_657; // @[Xbar.scala 246:36]
  wire  _T_659 = auto_out_4_b_valid & requestBOI_4_0; // @[Xbar.scala 222:40]
  wire  _T_2064 = _T_2063 | _T_659; // @[Xbar.scala 246:36]
  wire  _T_661 = auto_out_5_b_valid & requestBOI_5_0; // @[Xbar.scala 222:40]
  wire  _T_2065 = _T_2064 | _T_661; // @[Xbar.scala 246:36]
  wire  _T_663 = auto_out_6_b_valid & requestBOI_6_0; // @[Xbar.scala 222:40]
  wire  _T_2066 = _T_2065 | _T_663; // @[Xbar.scala 246:36]
  wire  _T_665 = auto_out_7_b_valid & requestBOI_7_0; // @[Xbar.scala 222:40]
  wire  _T_2067 = _T_2066 | _T_665; // @[Xbar.scala 246:36]
  wire  _T_667 = auto_out_8_b_valid & requestBOI_8_0; // @[Xbar.scala 222:40]
  wire  _T_2068 = _T_2067 | _T_667; // @[Xbar.scala 246:36]
  wire  _T_669 = auto_out_9_b_valid & requestBOI_9_0; // @[Xbar.scala 222:40]
  wire  _T_2069 = _T_2068 | _T_669; // @[Xbar.scala 246:36]
  wire  _T_671 = auto_out_10_b_valid & requestBOI_10_0; // @[Xbar.scala 222:40]
  wire  _T_2070 = _T_2069 | _T_671; // @[Xbar.scala 246:36]
  wire  _T_673 = auto_out_11_b_valid & requestBOI_11_0; // @[Xbar.scala 222:40]
  wire  _T_2071 = _T_2070 | _T_673; // @[Xbar.scala 246:36]
  wire  _T_675 = auto_out_12_b_valid & requestBOI_12_0; // @[Xbar.scala 222:40]
  wire  _T_2072 = _T_2071 | _T_675; // @[Xbar.scala 246:36]
  wire  _T_677 = auto_out_13_b_valid & requestBOI_13_0; // @[Xbar.scala 222:40]
  wire  _T_2073 = _T_2072 | _T_677; // @[Xbar.scala 246:36]
  wire  _T_679 = auto_out_14_b_valid & requestBOI_14_0; // @[Xbar.scala 222:40]
  wire  _T_2074 = _T_2073 | _T_679; // @[Xbar.scala 246:36]
  wire  _T_681 = auto_out_15_b_valid & requestBOI_15_0; // @[Xbar.scala 222:40]
  wire  _T_2075 = _T_2074 | _T_681; // @[Xbar.scala 246:36]
  wire  _T_683 = auto_out_16_b_valid & requestBOI_16_0; // @[Xbar.scala 222:40]
  wire  _T_2076 = _T_2075 | _T_683; // @[Xbar.scala 246:36]
  wire  _T_685 = auto_out_17_b_valid & requestBOI_17_0; // @[Xbar.scala 222:40]
  wire  _T_2077 = _T_2076 | _T_685; // @[Xbar.scala 246:36]
  wire  _T_687 = auto_out_18_b_valid & requestBOI_18_0; // @[Xbar.scala 222:40]
  wire  _T_2078 = _T_2077 | _T_687; // @[Xbar.scala 246:36]
  wire  _T_689 = auto_out_19_b_valid & requestBOI_19_0; // @[Xbar.scala 222:40]
  wire  _T_2079 = _T_2078 | _T_689; // @[Xbar.scala 246:36]
  wire  _T_2080 = _T_2079 | auto_out_20_b_valid; // @[Xbar.scala 246:36]
  reg  _T_2326_0; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_29;
  wire  _T_2351 = _T_2326_0 & _T_651; // @[Mux.scala 27:72]
  reg  _T_2326_1; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_30;
  wire  _T_2352 = _T_2326_1 & _T_653; // @[Mux.scala 27:72]
  wire  _T_2372 = _T_2351 | _T_2352; // @[Mux.scala 27:72]
  reg  _T_2326_2; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_31;
  wire  _T_2353 = _T_2326_2 & _T_655; // @[Mux.scala 27:72]
  wire  _T_2373 = _T_2372 | _T_2353; // @[Mux.scala 27:72]
  reg  _T_2326_3; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_32;
  wire  _T_2354 = _T_2326_3 & _T_657; // @[Mux.scala 27:72]
  wire  _T_2374 = _T_2373 | _T_2354; // @[Mux.scala 27:72]
  reg  _T_2326_4; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_33;
  wire  _T_2355 = _T_2326_4 & _T_659; // @[Mux.scala 27:72]
  wire  _T_2375 = _T_2374 | _T_2355; // @[Mux.scala 27:72]
  reg  _T_2326_5; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_34;
  wire  _T_2356 = _T_2326_5 & _T_661; // @[Mux.scala 27:72]
  wire  _T_2376 = _T_2375 | _T_2356; // @[Mux.scala 27:72]
  reg  _T_2326_6; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_35;
  wire  _T_2357 = _T_2326_6 & _T_663; // @[Mux.scala 27:72]
  wire  _T_2377 = _T_2376 | _T_2357; // @[Mux.scala 27:72]
  reg  _T_2326_7; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_36;
  wire  _T_2358 = _T_2326_7 & _T_665; // @[Mux.scala 27:72]
  wire  _T_2378 = _T_2377 | _T_2358; // @[Mux.scala 27:72]
  reg  _T_2326_8; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_37;
  wire  _T_2359 = _T_2326_8 & _T_667; // @[Mux.scala 27:72]
  wire  _T_2379 = _T_2378 | _T_2359; // @[Mux.scala 27:72]
  reg  _T_2326_9; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_38;
  wire  _T_2360 = _T_2326_9 & _T_669; // @[Mux.scala 27:72]
  wire  _T_2380 = _T_2379 | _T_2360; // @[Mux.scala 27:72]
  reg  _T_2326_10; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_39;
  wire  _T_2361 = _T_2326_10 & _T_671; // @[Mux.scala 27:72]
  wire  _T_2381 = _T_2380 | _T_2361; // @[Mux.scala 27:72]
  reg  _T_2326_11; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_40;
  wire  _T_2362 = _T_2326_11 & _T_673; // @[Mux.scala 27:72]
  wire  _T_2382 = _T_2381 | _T_2362; // @[Mux.scala 27:72]
  reg  _T_2326_12; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_41;
  wire  _T_2363 = _T_2326_12 & _T_675; // @[Mux.scala 27:72]
  wire  _T_2383 = _T_2382 | _T_2363; // @[Mux.scala 27:72]
  reg  _T_2326_13; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_42;
  wire  _T_2364 = _T_2326_13 & _T_677; // @[Mux.scala 27:72]
  wire  _T_2384 = _T_2383 | _T_2364; // @[Mux.scala 27:72]
  reg  _T_2326_14; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_43;
  wire  _T_2365 = _T_2326_14 & _T_679; // @[Mux.scala 27:72]
  wire  _T_2385 = _T_2384 | _T_2365; // @[Mux.scala 27:72]
  reg  _T_2326_15; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_44;
  wire  _T_2366 = _T_2326_15 & _T_681; // @[Mux.scala 27:72]
  wire  _T_2386 = _T_2385 | _T_2366; // @[Mux.scala 27:72]
  reg  _T_2326_16; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_45;
  wire  _T_2367 = _T_2326_16 & _T_683; // @[Mux.scala 27:72]
  wire  _T_2387 = _T_2386 | _T_2367; // @[Mux.scala 27:72]
  reg  _T_2326_17; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_46;
  wire  _T_2368 = _T_2326_17 & _T_685; // @[Mux.scala 27:72]
  wire  _T_2388 = _T_2387 | _T_2368; // @[Mux.scala 27:72]
  reg  _T_2326_18; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_47;
  wire  _T_2369 = _T_2326_18 & _T_687; // @[Mux.scala 27:72]
  wire  _T_2389 = _T_2388 | _T_2369; // @[Mux.scala 27:72]
  reg  _T_2326_19; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_48;
  wire  _T_2370 = _T_2326_19 & _T_689; // @[Mux.scala 27:72]
  wire  _T_2390 = _T_2389 | _T_2370; // @[Mux.scala 27:72]
  reg  _T_2326_20; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_49;
  wire  _T_2371 = _T_2326_20 & auto_out_20_b_valid; // @[Mux.scala 27:72]
  wire  _T_2391 = _T_2390 | _T_2371; // @[Mux.scala 27:72]
  wire  in_0_b_valid = _T_2060 ? _T_2080 : _T_2391; // @[Xbar.scala 278:22]
  wire  _T_373 = auto_in_b_ready & in_0_b_valid; // @[Decoupled.scala 40:37]
  wire [2:0] _GEN_104 = {{2'd0}, _T_371}; // @[Xbar.scala 106:30]
  wire [2:0] _T_378 = _T_375 + _GEN_104; // @[Xbar.scala 106:30]
  wire [2:0] _GEN_105 = {{2'd0}, _T_373}; // @[Xbar.scala 106:48]
  wire [2:0] _T_380 = _T_378 - _GEN_105; // @[Xbar.scala 106:48]
  wire  _T_381 = ~_T_373; // @[Xbar.scala 107:23]
  wire  _T_382 = _T_375 != 3'h0; // @[Xbar.scala 107:43]
  wire  _T_383 = _T_381 | _T_382; // @[Xbar.scala 107:34]
  wire  _T_385 = _T_383 | reset; // @[Xbar.scala 107:22]
  wire  _T_386 = ~_T_385; // @[Xbar.scala 107:22]
  wire  _T_387 = ~_T_371; // @[Xbar.scala 108:23]
  wire  _T_389 = _T_387 | _T_396; // @[Xbar.scala 108:34]
  wire  _T_391 = _T_389 | reset; // @[Xbar.scala 108:22]
  wire  _T_392 = ~_T_391; // @[Xbar.scala 108:22]
  wire  in_0_ar_valid = auto_in_ar_valid & _T_370; // @[Xbar.scala 129:45]
  wire  _T_403 = auto_in_aw_valid & _T_405; // @[Xbar.scala 138:45]
  wire  in_0_aw_valid = _T_403 & _T_398; // @[Xbar.scala 138:82]
  wire  _T_408 = ~_T_401; // @[Xbar.scala 140:54]
  wire  _T_410 = awIn_0_io_enq_ready & awIn_0_io_enq_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_2 = _T_410 | _T_401; // @[Xbar.scala 141:38]
  wire  _T_411 = in_0_aw_ready & in_0_aw_valid; // @[Decoupled.scala 40:37]
  wire  in_0_w_valid = auto_in_w_valid & awIn_0_io_deq_valid; // @[Xbar.scala 145:43]
  wire  _T_566 = requestWIO_0_0 & auto_out_0_w_ready; // @[Mux.scala 27:72]
  wire  _T_567 = requestWIO_0_1 & auto_out_1_w_ready; // @[Mux.scala 27:72]
  wire  _T_587 = _T_566 | _T_567; // @[Mux.scala 27:72]
  wire  _T_568 = requestWIO_0_2 & auto_out_2_w_ready; // @[Mux.scala 27:72]
  wire  _T_588 = _T_587 | _T_568; // @[Mux.scala 27:72]
  wire  _T_569 = requestWIO_0_3 & auto_out_3_w_ready; // @[Mux.scala 27:72]
  wire  _T_589 = _T_588 | _T_569; // @[Mux.scala 27:72]
  wire  _T_570 = requestWIO_0_4 & auto_out_4_w_ready; // @[Mux.scala 27:72]
  wire  _T_590 = _T_589 | _T_570; // @[Mux.scala 27:72]
  wire  _T_571 = requestWIO_0_5 & auto_out_5_w_ready; // @[Mux.scala 27:72]
  wire  _T_591 = _T_590 | _T_571; // @[Mux.scala 27:72]
  wire  _T_572 = requestWIO_0_6 & auto_out_6_w_ready; // @[Mux.scala 27:72]
  wire  _T_592 = _T_591 | _T_572; // @[Mux.scala 27:72]
  wire  _T_573 = requestWIO_0_7 & auto_out_7_w_ready; // @[Mux.scala 27:72]
  wire  _T_593 = _T_592 | _T_573; // @[Mux.scala 27:72]
  wire  _T_574 = requestWIO_0_8 & auto_out_8_w_ready; // @[Mux.scala 27:72]
  wire  _T_594 = _T_593 | _T_574; // @[Mux.scala 27:72]
  wire  _T_575 = requestWIO_0_9 & auto_out_9_w_ready; // @[Mux.scala 27:72]
  wire  _T_595 = _T_594 | _T_575; // @[Mux.scala 27:72]
  wire  _T_576 = requestWIO_0_10 & auto_out_10_w_ready; // @[Mux.scala 27:72]
  wire  _T_596 = _T_595 | _T_576; // @[Mux.scala 27:72]
  wire  _T_577 = requestWIO_0_11 & auto_out_11_w_ready; // @[Mux.scala 27:72]
  wire  _T_597 = _T_596 | _T_577; // @[Mux.scala 27:72]
  wire  _T_578 = requestWIO_0_12 & auto_out_12_w_ready; // @[Mux.scala 27:72]
  wire  _T_598 = _T_597 | _T_578; // @[Mux.scala 27:72]
  wire  _T_579 = requestWIO_0_13 & auto_out_13_w_ready; // @[Mux.scala 27:72]
  wire  _T_599 = _T_598 | _T_579; // @[Mux.scala 27:72]
  wire  _T_580 = requestWIO_0_14 & auto_out_14_w_ready; // @[Mux.scala 27:72]
  wire  _T_600 = _T_599 | _T_580; // @[Mux.scala 27:72]
  wire  _T_581 = requestWIO_0_15 & auto_out_15_w_ready; // @[Mux.scala 27:72]
  wire  _T_601 = _T_600 | _T_581; // @[Mux.scala 27:72]
  wire  _T_582 = requestWIO_0_16 & auto_out_16_w_ready; // @[Mux.scala 27:72]
  wire  _T_602 = _T_601 | _T_582; // @[Mux.scala 27:72]
  wire  _T_583 = requestWIO_0_17 & auto_out_17_w_ready; // @[Mux.scala 27:72]
  wire  _T_603 = _T_602 | _T_583; // @[Mux.scala 27:72]
  wire  _T_584 = requestWIO_0_18 & auto_out_18_w_ready; // @[Mux.scala 27:72]
  wire  _T_604 = _T_603 | _T_584; // @[Mux.scala 27:72]
  wire  _T_585 = requestWIO_0_19 & auto_out_19_w_ready; // @[Mux.scala 27:72]
  wire  _T_605 = _T_604 | _T_585; // @[Mux.scala 27:72]
  wire  _T_586 = requestWIO_0_20 & auto_out_20_w_ready; // @[Mux.scala 27:72]
  wire  in_0_w_ready = _T_605 | _T_586; // @[Mux.scala 27:72]
  wire  _T_414 = auto_in_w_valid & auto_in_w_bits_last; // @[Xbar.scala 147:50]
  wire  out_0_ar_valid = in_0_ar_valid & requestARIO_0_0; // @[Xbar.scala 222:40]
  wire  out_1_ar_valid = in_0_ar_valid & requestARIO_0_1; // @[Xbar.scala 222:40]
  wire  out_2_ar_valid = in_0_ar_valid & requestARIO_0_2; // @[Xbar.scala 222:40]
  wire  out_3_ar_valid = in_0_ar_valid & requestARIO_0_3; // @[Xbar.scala 222:40]
  wire  out_4_ar_valid = in_0_ar_valid & requestARIO_0_4; // @[Xbar.scala 222:40]
  wire  out_5_ar_valid = in_0_ar_valid & requestARIO_0_5; // @[Xbar.scala 222:40]
  wire  out_6_ar_valid = in_0_ar_valid & requestARIO_0_6; // @[Xbar.scala 222:40]
  wire  out_7_ar_valid = in_0_ar_valid & requestARIO_0_7; // @[Xbar.scala 222:40]
  wire  out_8_ar_valid = in_0_ar_valid & requestARIO_0_8; // @[Xbar.scala 222:40]
  wire  out_9_ar_valid = in_0_ar_valid & requestARIO_0_9; // @[Xbar.scala 222:40]
  wire  out_10_ar_valid = in_0_ar_valid & requestARIO_0_10; // @[Xbar.scala 222:40]
  wire  out_11_ar_valid = in_0_ar_valid & requestARIO_0_11; // @[Xbar.scala 222:40]
  wire  out_12_ar_valid = in_0_ar_valid & requestARIO_0_12; // @[Xbar.scala 222:40]
  wire  out_13_ar_valid = in_0_ar_valid & requestARIO_0_13; // @[Xbar.scala 222:40]
  wire  out_14_ar_valid = in_0_ar_valid & requestARIO_0_14; // @[Xbar.scala 222:40]
  wire  out_15_ar_valid = in_0_ar_valid & requestARIO_0_15; // @[Xbar.scala 222:40]
  wire  out_16_ar_valid = in_0_ar_valid & requestARIO_0_16; // @[Xbar.scala 222:40]
  wire  out_17_ar_valid = in_0_ar_valid & requestARIO_0_17; // @[Xbar.scala 222:40]
  wire  out_18_ar_valid = in_0_ar_valid & requestARIO_0_18; // @[Xbar.scala 222:40]
  wire  out_19_ar_valid = in_0_ar_valid & requestARIO_0_19; // @[Xbar.scala 222:40]
  wire  out_20_ar_valid = in_0_ar_valid & requestARIO_0_20; // @[Xbar.scala 222:40]
  wire  out_0_aw_valid = in_0_aw_valid & requestAWIO_0_0; // @[Xbar.scala 222:40]
  wire  out_1_aw_valid = in_0_aw_valid & requestAWIO_0_1; // @[Xbar.scala 222:40]
  wire  out_2_aw_valid = in_0_aw_valid & requestAWIO_0_2; // @[Xbar.scala 222:40]
  wire  out_3_aw_valid = in_0_aw_valid & requestAWIO_0_3; // @[Xbar.scala 222:40]
  wire  out_4_aw_valid = in_0_aw_valid & requestAWIO_0_4; // @[Xbar.scala 222:40]
  wire  out_5_aw_valid = in_0_aw_valid & requestAWIO_0_5; // @[Xbar.scala 222:40]
  wire  out_6_aw_valid = in_0_aw_valid & requestAWIO_0_6; // @[Xbar.scala 222:40]
  wire  out_7_aw_valid = in_0_aw_valid & requestAWIO_0_7; // @[Xbar.scala 222:40]
  wire  out_8_aw_valid = in_0_aw_valid & requestAWIO_0_8; // @[Xbar.scala 222:40]
  wire  out_9_aw_valid = in_0_aw_valid & requestAWIO_0_9; // @[Xbar.scala 222:40]
  wire  out_10_aw_valid = in_0_aw_valid & requestAWIO_0_10; // @[Xbar.scala 222:40]
  wire  out_11_aw_valid = in_0_aw_valid & requestAWIO_0_11; // @[Xbar.scala 222:40]
  wire  out_12_aw_valid = in_0_aw_valid & requestAWIO_0_12; // @[Xbar.scala 222:40]
  wire  out_13_aw_valid = in_0_aw_valid & requestAWIO_0_13; // @[Xbar.scala 222:40]
  wire  out_14_aw_valid = in_0_aw_valid & requestAWIO_0_14; // @[Xbar.scala 222:40]
  wire  out_15_aw_valid = in_0_aw_valid & requestAWIO_0_15; // @[Xbar.scala 222:40]
  wire  out_16_aw_valid = in_0_aw_valid & requestAWIO_0_16; // @[Xbar.scala 222:40]
  wire  out_17_aw_valid = in_0_aw_valid & requestAWIO_0_17; // @[Xbar.scala 222:40]
  wire  out_18_aw_valid = in_0_aw_valid & requestAWIO_0_18; // @[Xbar.scala 222:40]
  wire  out_19_aw_valid = in_0_aw_valid & requestAWIO_0_19; // @[Xbar.scala 222:40]
  wire  out_20_aw_valid = in_0_aw_valid & requestAWIO_0_20; // @[Xbar.scala 222:40]
  wire  _T_698 = ~out_0_aw_valid; // @[Xbar.scala 256:60]
  wire  _T_704 = _T_698 | out_0_aw_valid; // @[Xbar.scala 258:23]
  wire  _T_706 = _T_704 | reset; // @[Xbar.scala 258:12]
  wire  _T_707 = ~_T_706; // @[Xbar.scala 258:12]
  wire  _T_719 = ~out_0_ar_valid; // @[Xbar.scala 256:60]
  wire  _T_725 = _T_719 | out_0_ar_valid; // @[Xbar.scala 258:23]
  wire  _T_727 = _T_725 | reset; // @[Xbar.scala 258:12]
  wire  _T_728 = ~_T_727; // @[Xbar.scala 258:12]
  wire  _T_742 = ~out_1_aw_valid; // @[Xbar.scala 256:60]
  wire  _T_748 = _T_742 | out_1_aw_valid; // @[Xbar.scala 258:23]
  wire  _T_750 = _T_748 | reset; // @[Xbar.scala 258:12]
  wire  _T_751 = ~_T_750; // @[Xbar.scala 258:12]
  wire  _T_763 = ~out_1_ar_valid; // @[Xbar.scala 256:60]
  wire  _T_769 = _T_763 | out_1_ar_valid; // @[Xbar.scala 258:23]
  wire  _T_771 = _T_769 | reset; // @[Xbar.scala 258:12]
  wire  _T_772 = ~_T_771; // @[Xbar.scala 258:12]
  wire  _T_786 = ~out_2_aw_valid; // @[Xbar.scala 256:60]
  wire  _T_792 = _T_786 | out_2_aw_valid; // @[Xbar.scala 258:23]
  wire  _T_794 = _T_792 | reset; // @[Xbar.scala 258:12]
  wire  _T_795 = ~_T_794; // @[Xbar.scala 258:12]
  wire  _T_807 = ~out_2_ar_valid; // @[Xbar.scala 256:60]
  wire  _T_813 = _T_807 | out_2_ar_valid; // @[Xbar.scala 258:23]
  wire  _T_815 = _T_813 | reset; // @[Xbar.scala 258:12]
  wire  _T_816 = ~_T_815; // @[Xbar.scala 258:12]
  wire  _T_830 = ~out_3_aw_valid; // @[Xbar.scala 256:60]
  wire  _T_836 = _T_830 | out_3_aw_valid; // @[Xbar.scala 258:23]
  wire  _T_838 = _T_836 | reset; // @[Xbar.scala 258:12]
  wire  _T_839 = ~_T_838; // @[Xbar.scala 258:12]
  wire  _T_851 = ~out_3_ar_valid; // @[Xbar.scala 256:60]
  wire  _T_857 = _T_851 | out_3_ar_valid; // @[Xbar.scala 258:23]
  wire  _T_859 = _T_857 | reset; // @[Xbar.scala 258:12]
  wire  _T_860 = ~_T_859; // @[Xbar.scala 258:12]
  wire  _T_874 = ~out_4_aw_valid; // @[Xbar.scala 256:60]
  wire  _T_880 = _T_874 | out_4_aw_valid; // @[Xbar.scala 258:23]
  wire  _T_882 = _T_880 | reset; // @[Xbar.scala 258:12]
  wire  _T_883 = ~_T_882; // @[Xbar.scala 258:12]
  wire  _T_895 = ~out_4_ar_valid; // @[Xbar.scala 256:60]
  wire  _T_901 = _T_895 | out_4_ar_valid; // @[Xbar.scala 258:23]
  wire  _T_903 = _T_901 | reset; // @[Xbar.scala 258:12]
  wire  _T_904 = ~_T_903; // @[Xbar.scala 258:12]
  wire  _T_918 = ~out_5_aw_valid; // @[Xbar.scala 256:60]
  wire  _T_924 = _T_918 | out_5_aw_valid; // @[Xbar.scala 258:23]
  wire  _T_926 = _T_924 | reset; // @[Xbar.scala 258:12]
  wire  _T_927 = ~_T_926; // @[Xbar.scala 258:12]
  wire  _T_939 = ~out_5_ar_valid; // @[Xbar.scala 256:60]
  wire  _T_945 = _T_939 | out_5_ar_valid; // @[Xbar.scala 258:23]
  wire  _T_947 = _T_945 | reset; // @[Xbar.scala 258:12]
  wire  _T_948 = ~_T_947; // @[Xbar.scala 258:12]
  wire  _T_962 = ~out_6_aw_valid; // @[Xbar.scala 256:60]
  wire  _T_968 = _T_962 | out_6_aw_valid; // @[Xbar.scala 258:23]
  wire  _T_970 = _T_968 | reset; // @[Xbar.scala 258:12]
  wire  _T_971 = ~_T_970; // @[Xbar.scala 258:12]
  wire  _T_983 = ~out_6_ar_valid; // @[Xbar.scala 256:60]
  wire  _T_989 = _T_983 | out_6_ar_valid; // @[Xbar.scala 258:23]
  wire  _T_991 = _T_989 | reset; // @[Xbar.scala 258:12]
  wire  _T_992 = ~_T_991; // @[Xbar.scala 258:12]
  wire  _T_1006 = ~out_7_aw_valid; // @[Xbar.scala 256:60]
  wire  _T_1012 = _T_1006 | out_7_aw_valid; // @[Xbar.scala 258:23]
  wire  _T_1014 = _T_1012 | reset; // @[Xbar.scala 258:12]
  wire  _T_1015 = ~_T_1014; // @[Xbar.scala 258:12]
  wire  _T_1027 = ~out_7_ar_valid; // @[Xbar.scala 256:60]
  wire  _T_1033 = _T_1027 | out_7_ar_valid; // @[Xbar.scala 258:23]
  wire  _T_1035 = _T_1033 | reset; // @[Xbar.scala 258:12]
  wire  _T_1036 = ~_T_1035; // @[Xbar.scala 258:12]
  wire  _T_1050 = ~out_8_aw_valid; // @[Xbar.scala 256:60]
  wire  _T_1056 = _T_1050 | out_8_aw_valid; // @[Xbar.scala 258:23]
  wire  _T_1058 = _T_1056 | reset; // @[Xbar.scala 258:12]
  wire  _T_1059 = ~_T_1058; // @[Xbar.scala 258:12]
  wire  _T_1071 = ~out_8_ar_valid; // @[Xbar.scala 256:60]
  wire  _T_1077 = _T_1071 | out_8_ar_valid; // @[Xbar.scala 258:23]
  wire  _T_1079 = _T_1077 | reset; // @[Xbar.scala 258:12]
  wire  _T_1080 = ~_T_1079; // @[Xbar.scala 258:12]
  wire  _T_1094 = ~out_9_aw_valid; // @[Xbar.scala 256:60]
  wire  _T_1100 = _T_1094 | out_9_aw_valid; // @[Xbar.scala 258:23]
  wire  _T_1102 = _T_1100 | reset; // @[Xbar.scala 258:12]
  wire  _T_1103 = ~_T_1102; // @[Xbar.scala 258:12]
  wire  _T_1115 = ~out_9_ar_valid; // @[Xbar.scala 256:60]
  wire  _T_1121 = _T_1115 | out_9_ar_valid; // @[Xbar.scala 258:23]
  wire  _T_1123 = _T_1121 | reset; // @[Xbar.scala 258:12]
  wire  _T_1124 = ~_T_1123; // @[Xbar.scala 258:12]
  wire  _T_1138 = ~out_10_aw_valid; // @[Xbar.scala 256:60]
  wire  _T_1144 = _T_1138 | out_10_aw_valid; // @[Xbar.scala 258:23]
  wire  _T_1146 = _T_1144 | reset; // @[Xbar.scala 258:12]
  wire  _T_1147 = ~_T_1146; // @[Xbar.scala 258:12]
  wire  _T_1159 = ~out_10_ar_valid; // @[Xbar.scala 256:60]
  wire  _T_1165 = _T_1159 | out_10_ar_valid; // @[Xbar.scala 258:23]
  wire  _T_1167 = _T_1165 | reset; // @[Xbar.scala 258:12]
  wire  _T_1168 = ~_T_1167; // @[Xbar.scala 258:12]
  wire  _T_1182 = ~out_11_aw_valid; // @[Xbar.scala 256:60]
  wire  _T_1188 = _T_1182 | out_11_aw_valid; // @[Xbar.scala 258:23]
  wire  _T_1190 = _T_1188 | reset; // @[Xbar.scala 258:12]
  wire  _T_1191 = ~_T_1190; // @[Xbar.scala 258:12]
  wire  _T_1203 = ~out_11_ar_valid; // @[Xbar.scala 256:60]
  wire  _T_1209 = _T_1203 | out_11_ar_valid; // @[Xbar.scala 258:23]
  wire  _T_1211 = _T_1209 | reset; // @[Xbar.scala 258:12]
  wire  _T_1212 = ~_T_1211; // @[Xbar.scala 258:12]
  wire  _T_1226 = ~out_12_aw_valid; // @[Xbar.scala 256:60]
  wire  _T_1232 = _T_1226 | out_12_aw_valid; // @[Xbar.scala 258:23]
  wire  _T_1234 = _T_1232 | reset; // @[Xbar.scala 258:12]
  wire  _T_1235 = ~_T_1234; // @[Xbar.scala 258:12]
  wire  _T_1247 = ~out_12_ar_valid; // @[Xbar.scala 256:60]
  wire  _T_1253 = _T_1247 | out_12_ar_valid; // @[Xbar.scala 258:23]
  wire  _T_1255 = _T_1253 | reset; // @[Xbar.scala 258:12]
  wire  _T_1256 = ~_T_1255; // @[Xbar.scala 258:12]
  wire  _T_1270 = ~out_13_aw_valid; // @[Xbar.scala 256:60]
  wire  _T_1276 = _T_1270 | out_13_aw_valid; // @[Xbar.scala 258:23]
  wire  _T_1278 = _T_1276 | reset; // @[Xbar.scala 258:12]
  wire  _T_1279 = ~_T_1278; // @[Xbar.scala 258:12]
  wire  _T_1291 = ~out_13_ar_valid; // @[Xbar.scala 256:60]
  wire  _T_1297 = _T_1291 | out_13_ar_valid; // @[Xbar.scala 258:23]
  wire  _T_1299 = _T_1297 | reset; // @[Xbar.scala 258:12]
  wire  _T_1300 = ~_T_1299; // @[Xbar.scala 258:12]
  wire  _T_1314 = ~out_14_aw_valid; // @[Xbar.scala 256:60]
  wire  _T_1320 = _T_1314 | out_14_aw_valid; // @[Xbar.scala 258:23]
  wire  _T_1322 = _T_1320 | reset; // @[Xbar.scala 258:12]
  wire  _T_1323 = ~_T_1322; // @[Xbar.scala 258:12]
  wire  _T_1335 = ~out_14_ar_valid; // @[Xbar.scala 256:60]
  wire  _T_1341 = _T_1335 | out_14_ar_valid; // @[Xbar.scala 258:23]
  wire  _T_1343 = _T_1341 | reset; // @[Xbar.scala 258:12]
  wire  _T_1344 = ~_T_1343; // @[Xbar.scala 258:12]
  wire  _T_1358 = ~out_15_aw_valid; // @[Xbar.scala 256:60]
  wire  _T_1364 = _T_1358 | out_15_aw_valid; // @[Xbar.scala 258:23]
  wire  _T_1366 = _T_1364 | reset; // @[Xbar.scala 258:12]
  wire  _T_1367 = ~_T_1366; // @[Xbar.scala 258:12]
  wire  _T_1379 = ~out_15_ar_valid; // @[Xbar.scala 256:60]
  wire  _T_1385 = _T_1379 | out_15_ar_valid; // @[Xbar.scala 258:23]
  wire  _T_1387 = _T_1385 | reset; // @[Xbar.scala 258:12]
  wire  _T_1388 = ~_T_1387; // @[Xbar.scala 258:12]
  wire  _T_1402 = ~out_16_aw_valid; // @[Xbar.scala 256:60]
  wire  _T_1408 = _T_1402 | out_16_aw_valid; // @[Xbar.scala 258:23]
  wire  _T_1410 = _T_1408 | reset; // @[Xbar.scala 258:12]
  wire  _T_1411 = ~_T_1410; // @[Xbar.scala 258:12]
  wire  _T_1423 = ~out_16_ar_valid; // @[Xbar.scala 256:60]
  wire  _T_1429 = _T_1423 | out_16_ar_valid; // @[Xbar.scala 258:23]
  wire  _T_1431 = _T_1429 | reset; // @[Xbar.scala 258:12]
  wire  _T_1432 = ~_T_1431; // @[Xbar.scala 258:12]
  wire  _T_1446 = ~out_17_aw_valid; // @[Xbar.scala 256:60]
  wire  _T_1452 = _T_1446 | out_17_aw_valid; // @[Xbar.scala 258:23]
  wire  _T_1454 = _T_1452 | reset; // @[Xbar.scala 258:12]
  wire  _T_1455 = ~_T_1454; // @[Xbar.scala 258:12]
  wire  _T_1467 = ~out_17_ar_valid; // @[Xbar.scala 256:60]
  wire  _T_1473 = _T_1467 | out_17_ar_valid; // @[Xbar.scala 258:23]
  wire  _T_1475 = _T_1473 | reset; // @[Xbar.scala 258:12]
  wire  _T_1476 = ~_T_1475; // @[Xbar.scala 258:12]
  wire  _T_1490 = ~out_18_aw_valid; // @[Xbar.scala 256:60]
  wire  _T_1496 = _T_1490 | out_18_aw_valid; // @[Xbar.scala 258:23]
  wire  _T_1498 = _T_1496 | reset; // @[Xbar.scala 258:12]
  wire  _T_1499 = ~_T_1498; // @[Xbar.scala 258:12]
  wire  _T_1511 = ~out_18_ar_valid; // @[Xbar.scala 256:60]
  wire  _T_1517 = _T_1511 | out_18_ar_valid; // @[Xbar.scala 258:23]
  wire  _T_1519 = _T_1517 | reset; // @[Xbar.scala 258:12]
  wire  _T_1520 = ~_T_1519; // @[Xbar.scala 258:12]
  wire  _T_1534 = ~out_19_aw_valid; // @[Xbar.scala 256:60]
  wire  _T_1540 = _T_1534 | out_19_aw_valid; // @[Xbar.scala 258:23]
  wire  _T_1542 = _T_1540 | reset; // @[Xbar.scala 258:12]
  wire  _T_1543 = ~_T_1542; // @[Xbar.scala 258:12]
  wire  _T_1555 = ~out_19_ar_valid; // @[Xbar.scala 256:60]
  wire  _T_1561 = _T_1555 | out_19_ar_valid; // @[Xbar.scala 258:23]
  wire  _T_1563 = _T_1561 | reset; // @[Xbar.scala 258:12]
  wire  _T_1564 = ~_T_1563; // @[Xbar.scala 258:12]
  wire  _T_1578 = ~out_20_aw_valid; // @[Xbar.scala 256:60]
  wire  _T_1584 = _T_1578 | out_20_aw_valid; // @[Xbar.scala 258:23]
  wire  _T_1586 = _T_1584 | reset; // @[Xbar.scala 258:12]
  wire  _T_1587 = ~_T_1586; // @[Xbar.scala 258:12]
  wire  _T_1599 = ~out_20_ar_valid; // @[Xbar.scala 256:60]
  wire  _T_1605 = _T_1599 | out_20_ar_valid; // @[Xbar.scala 258:23]
  wire  _T_1607 = _T_1605 | reset; // @[Xbar.scala 258:12]
  wire  _T_1608 = ~_T_1607; // @[Xbar.scala 258:12]
  wire  _T_1685 = _T_1656 != 21'h0; // @[Arbiter.scala 24:27]
  wire  _T_1686 = _T_1616 & _T_1685; // @[Arbiter.scala 24:18]
  wire [20:0] _T_1687 = _T_1684 & _T_1656; // @[Arbiter.scala 25:29]
  wire [21:0] _T_1688 = {_T_1687, 1'h0}; // @[package.scala 199:48]
  wire [20:0] _T_1690 = _T_1687 | _T_1688[20:0]; // @[package.scala 199:43]
  wire [22:0] _T_1691 = {_T_1690, 2'h0}; // @[package.scala 199:48]
  wire [20:0] _T_1693 = _T_1690 | _T_1691[20:0]; // @[package.scala 199:43]
  wire [24:0] _T_1694 = {_T_1693, 4'h0}; // @[package.scala 199:48]
  wire [20:0] _T_1696 = _T_1693 | _T_1694[20:0]; // @[package.scala 199:43]
  wire [28:0] _T_1697 = {_T_1696, 8'h0}; // @[package.scala 199:48]
  wire [20:0] _T_1699 = _T_1696 | _T_1697[20:0]; // @[package.scala 199:43]
  wire [36:0] _T_1700 = {_T_1699, 16'h0}; // @[package.scala 199:48]
  wire [20:0] _T_1702 = _T_1699 | _T_1700[20:0]; // @[package.scala 199:43]
  wire  _T_1750 = _T_1727 | _T_1728; // @[Xbar.scala 255:50]
  wire  _T_1751 = _T_1750 | _T_1729; // @[Xbar.scala 255:50]
  wire  _T_1752 = _T_1751 | _T_1730; // @[Xbar.scala 255:50]
  wire  _T_1753 = _T_1752 | _T_1731; // @[Xbar.scala 255:50]
  wire  _T_1754 = _T_1753 | _T_1732; // @[Xbar.scala 255:50]
  wire  _T_1755 = _T_1754 | _T_1733; // @[Xbar.scala 255:50]
  wire  _T_1756 = _T_1755 | _T_1734; // @[Xbar.scala 255:50]
  wire  _T_1757 = _T_1756 | _T_1735; // @[Xbar.scala 255:50]
  wire  _T_1758 = _T_1757 | _T_1736; // @[Xbar.scala 255:50]
  wire  _T_1759 = _T_1758 | _T_1737; // @[Xbar.scala 255:50]
  wire  _T_1760 = _T_1759 | _T_1738; // @[Xbar.scala 255:50]
  wire  _T_1761 = _T_1760 | _T_1739; // @[Xbar.scala 255:50]
  wire  _T_1762 = _T_1761 | _T_1740; // @[Xbar.scala 255:50]
  wire  _T_1763 = _T_1762 | _T_1741; // @[Xbar.scala 255:50]
  wire  _T_1764 = _T_1763 | _T_1742; // @[Xbar.scala 255:50]
  wire  _T_1765 = _T_1764 | _T_1743; // @[Xbar.scala 255:50]
  wire  _T_1766 = _T_1765 | _T_1744; // @[Xbar.scala 255:50]
  wire  _T_1767 = _T_1766 | _T_1745; // @[Xbar.scala 255:50]
  wire  _T_1768 = _T_1767 | _T_1746; // @[Xbar.scala 255:50]
  wire  _T_1769 = _T_1768 | _T_1747; // @[Xbar.scala 255:50]
  wire  _T_1771 = ~_T_1727; // @[Xbar.scala 256:60]
  wire  _T_1774 = ~_T_1728; // @[Xbar.scala 256:60]
  wire  _T_1775 = _T_1771 | _T_1774; // @[Xbar.scala 256:57]
  wire  _T_1776 = ~_T_1750; // @[Xbar.scala 256:54]
  wire  _T_1777 = ~_T_1729; // @[Xbar.scala 256:60]
  wire  _T_1778 = _T_1776 | _T_1777; // @[Xbar.scala 256:57]
  wire  _T_1779 = ~_T_1751; // @[Xbar.scala 256:54]
  wire  _T_1780 = ~_T_1730; // @[Xbar.scala 256:60]
  wire  _T_1781 = _T_1779 | _T_1780; // @[Xbar.scala 256:57]
  wire  _T_1782 = ~_T_1752; // @[Xbar.scala 256:54]
  wire  _T_1783 = ~_T_1731; // @[Xbar.scala 256:60]
  wire  _T_1784 = _T_1782 | _T_1783; // @[Xbar.scala 256:57]
  wire  _T_1785 = ~_T_1753; // @[Xbar.scala 256:54]
  wire  _T_1786 = ~_T_1732; // @[Xbar.scala 256:60]
  wire  _T_1787 = _T_1785 | _T_1786; // @[Xbar.scala 256:57]
  wire  _T_1788 = ~_T_1754; // @[Xbar.scala 256:54]
  wire  _T_1789 = ~_T_1733; // @[Xbar.scala 256:60]
  wire  _T_1790 = _T_1788 | _T_1789; // @[Xbar.scala 256:57]
  wire  _T_1791 = ~_T_1755; // @[Xbar.scala 256:54]
  wire  _T_1792 = ~_T_1734; // @[Xbar.scala 256:60]
  wire  _T_1793 = _T_1791 | _T_1792; // @[Xbar.scala 256:57]
  wire  _T_1794 = ~_T_1756; // @[Xbar.scala 256:54]
  wire  _T_1795 = ~_T_1735; // @[Xbar.scala 256:60]
  wire  _T_1796 = _T_1794 | _T_1795; // @[Xbar.scala 256:57]
  wire  _T_1797 = ~_T_1757; // @[Xbar.scala 256:54]
  wire  _T_1798 = ~_T_1736; // @[Xbar.scala 256:60]
  wire  _T_1799 = _T_1797 | _T_1798; // @[Xbar.scala 256:57]
  wire  _T_1800 = ~_T_1758; // @[Xbar.scala 256:54]
  wire  _T_1801 = ~_T_1737; // @[Xbar.scala 256:60]
  wire  _T_1802 = _T_1800 | _T_1801; // @[Xbar.scala 256:57]
  wire  _T_1803 = ~_T_1759; // @[Xbar.scala 256:54]
  wire  _T_1804 = ~_T_1738; // @[Xbar.scala 256:60]
  wire  _T_1805 = _T_1803 | _T_1804; // @[Xbar.scala 256:57]
  wire  _T_1806 = ~_T_1760; // @[Xbar.scala 256:54]
  wire  _T_1807 = ~_T_1739; // @[Xbar.scala 256:60]
  wire  _T_1808 = _T_1806 | _T_1807; // @[Xbar.scala 256:57]
  wire  _T_1809 = ~_T_1761; // @[Xbar.scala 256:54]
  wire  _T_1810 = ~_T_1740; // @[Xbar.scala 256:60]
  wire  _T_1811 = _T_1809 | _T_1810; // @[Xbar.scala 256:57]
  wire  _T_1812 = ~_T_1762; // @[Xbar.scala 256:54]
  wire  _T_1813 = ~_T_1741; // @[Xbar.scala 256:60]
  wire  _T_1814 = _T_1812 | _T_1813; // @[Xbar.scala 256:57]
  wire  _T_1815 = ~_T_1763; // @[Xbar.scala 256:54]
  wire  _T_1816 = ~_T_1742; // @[Xbar.scala 256:60]
  wire  _T_1817 = _T_1815 | _T_1816; // @[Xbar.scala 256:57]
  wire  _T_1818 = ~_T_1764; // @[Xbar.scala 256:54]
  wire  _T_1819 = ~_T_1743; // @[Xbar.scala 256:60]
  wire  _T_1820 = _T_1818 | _T_1819; // @[Xbar.scala 256:57]
  wire  _T_1821 = ~_T_1765; // @[Xbar.scala 256:54]
  wire  _T_1822 = ~_T_1744; // @[Xbar.scala 256:60]
  wire  _T_1823 = _T_1821 | _T_1822; // @[Xbar.scala 256:57]
  wire  _T_1824 = ~_T_1766; // @[Xbar.scala 256:54]
  wire  _T_1825 = ~_T_1745; // @[Xbar.scala 256:60]
  wire  _T_1826 = _T_1824 | _T_1825; // @[Xbar.scala 256:57]
  wire  _T_1827 = ~_T_1767; // @[Xbar.scala 256:54]
  wire  _T_1828 = ~_T_1746; // @[Xbar.scala 256:60]
  wire  _T_1829 = _T_1827 | _T_1828; // @[Xbar.scala 256:57]
  wire  _T_1830 = ~_T_1768; // @[Xbar.scala 256:54]
  wire  _T_1831 = ~_T_1747; // @[Xbar.scala 256:60]
  wire  _T_1832 = _T_1830 | _T_1831; // @[Xbar.scala 256:57]
  wire  _T_1834 = _T_1775 & _T_1778; // @[Xbar.scala 256:75]
  wire  _T_1835 = _T_1834 & _T_1781; // @[Xbar.scala 256:75]
  wire  _T_1836 = _T_1835 & _T_1784; // @[Xbar.scala 256:75]
  wire  _T_1837 = _T_1836 & _T_1787; // @[Xbar.scala 256:75]
  wire  _T_1838 = _T_1837 & _T_1790; // @[Xbar.scala 256:75]
  wire  _T_1839 = _T_1838 & _T_1793; // @[Xbar.scala 256:75]
  wire  _T_1840 = _T_1839 & _T_1796; // @[Xbar.scala 256:75]
  wire  _T_1841 = _T_1840 & _T_1799; // @[Xbar.scala 256:75]
  wire  _T_1842 = _T_1841 & _T_1802; // @[Xbar.scala 256:75]
  wire  _T_1843 = _T_1842 & _T_1805; // @[Xbar.scala 256:75]
  wire  _T_1844 = _T_1843 & _T_1808; // @[Xbar.scala 256:75]
  wire  _T_1845 = _T_1844 & _T_1811; // @[Xbar.scala 256:75]
  wire  _T_1846 = _T_1845 & _T_1814; // @[Xbar.scala 256:75]
  wire  _T_1847 = _T_1846 & _T_1817; // @[Xbar.scala 256:75]
  wire  _T_1848 = _T_1847 & _T_1820; // @[Xbar.scala 256:75]
  wire  _T_1849 = _T_1848 & _T_1823; // @[Xbar.scala 256:75]
  wire  _T_1850 = _T_1849 & _T_1826; // @[Xbar.scala 256:75]
  wire  _T_1851 = _T_1850 & _T_1829; // @[Xbar.scala 256:75]
  wire  _T_1852 = _T_1851 & _T_1832; // @[Xbar.scala 256:75]
  wire  _T_1854 = _T_1852 | reset; // @[Xbar.scala 256:11]
  wire  _T_1855 = ~_T_1854; // @[Xbar.scala 256:11]
  wire  _T_1856 = ~_T_1636; // @[Xbar.scala 258:13]
  wire  _T_1877 = _T_1856 | _T_1769; // @[Xbar.scala 258:23]
  wire  _T_1879 = _T_1877 | reset; // @[Xbar.scala 258:12]
  wire  _T_1880 = ~_T_1879; // @[Xbar.scala 258:12]
  wire  _GEN_89 = _T_1636 ? 1'h0 : _T_1616; // @[Xbar.scala 266:21]
  wire  _GEN_90 = _T_344 | _GEN_89; // @[Xbar.scala 267:24]
  wire  _T_1885_0 = _T_1616 ? _T_1684[0] : _T_1882_0; // @[Xbar.scala 270:24]
  wire  _T_1885_1 = _T_1616 ? _T_1684[1] : _T_1882_1; // @[Xbar.scala 270:24]
  wire  _T_1885_2 = _T_1616 ? _T_1684[2] : _T_1882_2; // @[Xbar.scala 270:24]
  wire  _T_1885_3 = _T_1616 ? _T_1684[3] : _T_1882_3; // @[Xbar.scala 270:24]
  wire  _T_1885_4 = _T_1616 ? _T_1684[4] : _T_1882_4; // @[Xbar.scala 270:24]
  wire  _T_1885_5 = _T_1616 ? _T_1684[5] : _T_1882_5; // @[Xbar.scala 270:24]
  wire  _T_1885_6 = _T_1616 ? _T_1684[6] : _T_1882_6; // @[Xbar.scala 270:24]
  wire  _T_1885_7 = _T_1616 ? _T_1684[7] : _T_1882_7; // @[Xbar.scala 270:24]
  wire  _T_1885_8 = _T_1616 ? _T_1684[8] : _T_1882_8; // @[Xbar.scala 270:24]
  wire  _T_1885_9 = _T_1616 ? _T_1684[9] : _T_1882_9; // @[Xbar.scala 270:24]
  wire  _T_1885_10 = _T_1616 ? _T_1684[10] : _T_1882_10; // @[Xbar.scala 270:24]
  wire  _T_1885_11 = _T_1616 ? _T_1684[11] : _T_1882_11; // @[Xbar.scala 270:24]
  wire  _T_1885_12 = _T_1616 ? _T_1684[12] : _T_1882_12; // @[Xbar.scala 270:24]
  wire  _T_1885_13 = _T_1616 ? _T_1684[13] : _T_1882_13; // @[Xbar.scala 270:24]
  wire  _T_1885_14 = _T_1616 ? _T_1684[14] : _T_1882_14; // @[Xbar.scala 270:24]
  wire  _T_1885_15 = _T_1616 ? _T_1684[15] : _T_1882_15; // @[Xbar.scala 270:24]
  wire  _T_1885_16 = _T_1616 ? _T_1684[16] : _T_1882_16; // @[Xbar.scala 270:24]
  wire  _T_1885_17 = _T_1616 ? _T_1684[17] : _T_1882_17; // @[Xbar.scala 270:24]
  wire  _T_1885_18 = _T_1616 ? _T_1684[18] : _T_1882_18; // @[Xbar.scala 270:24]
  wire  _T_1885_19 = _T_1616 ? _T_1684[19] : _T_1882_19; // @[Xbar.scala 270:24]
  wire  _T_1885_20 = _T_1616 ? _T_1684[20] : _T_1882_20; // @[Xbar.scala 270:24]
  wire [9:0] _T_2089 = {_T_669,_T_667,_T_665,_T_663,_T_661,_T_659,_T_657,_T_655,_T_653,_T_651}; // @[Cat.scala 29:58]
  wire [4:0] _T_2093 = {_T_679,_T_677,_T_675,_T_673,_T_671}; // @[Cat.scala 29:58]
  wire [20:0] _T_2100 = {auto_out_20_b_valid,_T_689,_T_687,_T_685,_T_683,_T_681,_T_2093,_T_2089}; // @[Cat.scala 29:58]
  reg [20:0] _T_2107; // @[Arbiter.scala 20:23]
  reg [31:0] _RAND_50;
  wire [20:0] _T_2108 = ~_T_2107; // @[Arbiter.scala 21:30]
  wire [20:0] _T_2109 = _T_2100 & _T_2108; // @[Arbiter.scala 21:28]
  wire [41:0] _T_2110 = {_T_2109,auto_out_20_b_valid,_T_689,_T_687,_T_685,_T_683,_T_681,_T_2093,_T_2089}; // @[Cat.scala 29:58]
  wire [41:0] _GEN_106 = {{1'd0}, _T_2110[41:1]}; // @[package.scala 208:43]
  wire [41:0] _T_2112 = _T_2110 | _GEN_106; // @[package.scala 208:43]
  wire [41:0] _GEN_107 = {{2'd0}, _T_2112[41:2]}; // @[package.scala 208:43]
  wire [41:0] _T_2114 = _T_2112 | _GEN_107; // @[package.scala 208:43]
  wire [41:0] _GEN_108 = {{4'd0}, _T_2114[41:4]}; // @[package.scala 208:43]
  wire [41:0] _T_2116 = _T_2114 | _GEN_108; // @[package.scala 208:43]
  wire [41:0] _GEN_109 = {{8'd0}, _T_2116[41:8]}; // @[package.scala 208:43]
  wire [41:0] _T_2118 = _T_2116 | _GEN_109; // @[package.scala 208:43]
  wire [41:0] _GEN_110 = {{16'd0}, _T_2118[41:16]}; // @[package.scala 208:43]
  wire [41:0] _T_2120 = _T_2118 | _GEN_110; // @[package.scala 208:43]
  wire [41:0] _T_2123 = {_T_2107, 21'h0}; // @[Arbiter.scala 22:66]
  wire [41:0] _GEN_111 = {{1'd0}, _T_2120[41:1]}; // @[Arbiter.scala 22:58]
  wire [41:0] _T_2124 = _GEN_111 | _T_2123; // @[Arbiter.scala 22:58]
  wire [20:0] _T_2127 = _T_2124[41:21] & _T_2124[20:0]; // @[Arbiter.scala 23:39]
  wire [20:0] _T_2128 = ~_T_2127; // @[Arbiter.scala 23:18]
  wire  _T_2129 = _T_2100 != 21'h0; // @[Arbiter.scala 24:27]
  wire  _T_2130 = _T_2060 & _T_2129; // @[Arbiter.scala 24:18]
  wire [20:0] _T_2131 = _T_2128 & _T_2100; // @[Arbiter.scala 25:29]
  wire [21:0] _T_2132 = {_T_2131, 1'h0}; // @[package.scala 199:48]
  wire [20:0] _T_2134 = _T_2131 | _T_2132[20:0]; // @[package.scala 199:43]
  wire [22:0] _T_2135 = {_T_2134, 2'h0}; // @[package.scala 199:48]
  wire [20:0] _T_2137 = _T_2134 | _T_2135[20:0]; // @[package.scala 199:43]
  wire [24:0] _T_2138 = {_T_2137, 4'h0}; // @[package.scala 199:48]
  wire [20:0] _T_2140 = _T_2137 | _T_2138[20:0]; // @[package.scala 199:43]
  wire [28:0] _T_2141 = {_T_2140, 8'h0}; // @[package.scala 199:48]
  wire [20:0] _T_2143 = _T_2140 | _T_2141[20:0]; // @[package.scala 199:43]
  wire [36:0] _T_2144 = {_T_2143, 16'h0}; // @[package.scala 199:48]
  wire [20:0] _T_2146 = _T_2143 | _T_2144[20:0]; // @[package.scala 199:43]
  wire  _T_2171 = _T_2128[0] & _T_651; // @[Xbar.scala 250:63]
  wire  _T_2172 = _T_2128[1] & _T_653; // @[Xbar.scala 250:63]
  wire  _T_2173 = _T_2128[2] & _T_655; // @[Xbar.scala 250:63]
  wire  _T_2174 = _T_2128[3] & _T_657; // @[Xbar.scala 250:63]
  wire  _T_2175 = _T_2128[4] & _T_659; // @[Xbar.scala 250:63]
  wire  _T_2176 = _T_2128[5] & _T_661; // @[Xbar.scala 250:63]
  wire  _T_2177 = _T_2128[6] & _T_663; // @[Xbar.scala 250:63]
  wire  _T_2178 = _T_2128[7] & _T_665; // @[Xbar.scala 250:63]
  wire  _T_2179 = _T_2128[8] & _T_667; // @[Xbar.scala 250:63]
  wire  _T_2180 = _T_2128[9] & _T_669; // @[Xbar.scala 250:63]
  wire  _T_2181 = _T_2128[10] & _T_671; // @[Xbar.scala 250:63]
  wire  _T_2182 = _T_2128[11] & _T_673; // @[Xbar.scala 250:63]
  wire  _T_2183 = _T_2128[12] & _T_675; // @[Xbar.scala 250:63]
  wire  _T_2184 = _T_2128[13] & _T_677; // @[Xbar.scala 250:63]
  wire  _T_2185 = _T_2128[14] & _T_679; // @[Xbar.scala 250:63]
  wire  _T_2186 = _T_2128[15] & _T_681; // @[Xbar.scala 250:63]
  wire  _T_2187 = _T_2128[16] & _T_683; // @[Xbar.scala 250:63]
  wire  _T_2188 = _T_2128[17] & _T_685; // @[Xbar.scala 250:63]
  wire  _T_2189 = _T_2128[18] & _T_687; // @[Xbar.scala 250:63]
  wire  _T_2190 = _T_2128[19] & _T_689; // @[Xbar.scala 250:63]
  wire  _T_2191 = _T_2128[20] & auto_out_20_b_valid; // @[Xbar.scala 250:63]
  wire  _T_2194 = _T_2171 | _T_2172; // @[Xbar.scala 255:50]
  wire  _T_2195 = _T_2194 | _T_2173; // @[Xbar.scala 255:50]
  wire  _T_2196 = _T_2195 | _T_2174; // @[Xbar.scala 255:50]
  wire  _T_2197 = _T_2196 | _T_2175; // @[Xbar.scala 255:50]
  wire  _T_2198 = _T_2197 | _T_2176; // @[Xbar.scala 255:50]
  wire  _T_2199 = _T_2198 | _T_2177; // @[Xbar.scala 255:50]
  wire  _T_2200 = _T_2199 | _T_2178; // @[Xbar.scala 255:50]
  wire  _T_2201 = _T_2200 | _T_2179; // @[Xbar.scala 255:50]
  wire  _T_2202 = _T_2201 | _T_2180; // @[Xbar.scala 255:50]
  wire  _T_2203 = _T_2202 | _T_2181; // @[Xbar.scala 255:50]
  wire  _T_2204 = _T_2203 | _T_2182; // @[Xbar.scala 255:50]
  wire  _T_2205 = _T_2204 | _T_2183; // @[Xbar.scala 255:50]
  wire  _T_2206 = _T_2205 | _T_2184; // @[Xbar.scala 255:50]
  wire  _T_2207 = _T_2206 | _T_2185; // @[Xbar.scala 255:50]
  wire  _T_2208 = _T_2207 | _T_2186; // @[Xbar.scala 255:50]
  wire  _T_2209 = _T_2208 | _T_2187; // @[Xbar.scala 255:50]
  wire  _T_2210 = _T_2209 | _T_2188; // @[Xbar.scala 255:50]
  wire  _T_2211 = _T_2210 | _T_2189; // @[Xbar.scala 255:50]
  wire  _T_2212 = _T_2211 | _T_2190; // @[Xbar.scala 255:50]
  wire  _T_2213 = _T_2212 | _T_2191; // @[Xbar.scala 255:50]
  wire  _T_2215 = ~_T_2171; // @[Xbar.scala 256:60]
  wire  _T_2218 = ~_T_2172; // @[Xbar.scala 256:60]
  wire  _T_2219 = _T_2215 | _T_2218; // @[Xbar.scala 256:57]
  wire  _T_2220 = ~_T_2194; // @[Xbar.scala 256:54]
  wire  _T_2221 = ~_T_2173; // @[Xbar.scala 256:60]
  wire  _T_2222 = _T_2220 | _T_2221; // @[Xbar.scala 256:57]
  wire  _T_2223 = ~_T_2195; // @[Xbar.scala 256:54]
  wire  _T_2224 = ~_T_2174; // @[Xbar.scala 256:60]
  wire  _T_2225 = _T_2223 | _T_2224; // @[Xbar.scala 256:57]
  wire  _T_2226 = ~_T_2196; // @[Xbar.scala 256:54]
  wire  _T_2227 = ~_T_2175; // @[Xbar.scala 256:60]
  wire  _T_2228 = _T_2226 | _T_2227; // @[Xbar.scala 256:57]
  wire  _T_2229 = ~_T_2197; // @[Xbar.scala 256:54]
  wire  _T_2230 = ~_T_2176; // @[Xbar.scala 256:60]
  wire  _T_2231 = _T_2229 | _T_2230; // @[Xbar.scala 256:57]
  wire  _T_2232 = ~_T_2198; // @[Xbar.scala 256:54]
  wire  _T_2233 = ~_T_2177; // @[Xbar.scala 256:60]
  wire  _T_2234 = _T_2232 | _T_2233; // @[Xbar.scala 256:57]
  wire  _T_2235 = ~_T_2199; // @[Xbar.scala 256:54]
  wire  _T_2236 = ~_T_2178; // @[Xbar.scala 256:60]
  wire  _T_2237 = _T_2235 | _T_2236; // @[Xbar.scala 256:57]
  wire  _T_2238 = ~_T_2200; // @[Xbar.scala 256:54]
  wire  _T_2239 = ~_T_2179; // @[Xbar.scala 256:60]
  wire  _T_2240 = _T_2238 | _T_2239; // @[Xbar.scala 256:57]
  wire  _T_2241 = ~_T_2201; // @[Xbar.scala 256:54]
  wire  _T_2242 = ~_T_2180; // @[Xbar.scala 256:60]
  wire  _T_2243 = _T_2241 | _T_2242; // @[Xbar.scala 256:57]
  wire  _T_2244 = ~_T_2202; // @[Xbar.scala 256:54]
  wire  _T_2245 = ~_T_2181; // @[Xbar.scala 256:60]
  wire  _T_2246 = _T_2244 | _T_2245; // @[Xbar.scala 256:57]
  wire  _T_2247 = ~_T_2203; // @[Xbar.scala 256:54]
  wire  _T_2248 = ~_T_2182; // @[Xbar.scala 256:60]
  wire  _T_2249 = _T_2247 | _T_2248; // @[Xbar.scala 256:57]
  wire  _T_2250 = ~_T_2204; // @[Xbar.scala 256:54]
  wire  _T_2251 = ~_T_2183; // @[Xbar.scala 256:60]
  wire  _T_2252 = _T_2250 | _T_2251; // @[Xbar.scala 256:57]
  wire  _T_2253 = ~_T_2205; // @[Xbar.scala 256:54]
  wire  _T_2254 = ~_T_2184; // @[Xbar.scala 256:60]
  wire  _T_2255 = _T_2253 | _T_2254; // @[Xbar.scala 256:57]
  wire  _T_2256 = ~_T_2206; // @[Xbar.scala 256:54]
  wire  _T_2257 = ~_T_2185; // @[Xbar.scala 256:60]
  wire  _T_2258 = _T_2256 | _T_2257; // @[Xbar.scala 256:57]
  wire  _T_2259 = ~_T_2207; // @[Xbar.scala 256:54]
  wire  _T_2260 = ~_T_2186; // @[Xbar.scala 256:60]
  wire  _T_2261 = _T_2259 | _T_2260; // @[Xbar.scala 256:57]
  wire  _T_2262 = ~_T_2208; // @[Xbar.scala 256:54]
  wire  _T_2263 = ~_T_2187; // @[Xbar.scala 256:60]
  wire  _T_2264 = _T_2262 | _T_2263; // @[Xbar.scala 256:57]
  wire  _T_2265 = ~_T_2209; // @[Xbar.scala 256:54]
  wire  _T_2266 = ~_T_2188; // @[Xbar.scala 256:60]
  wire  _T_2267 = _T_2265 | _T_2266; // @[Xbar.scala 256:57]
  wire  _T_2268 = ~_T_2210; // @[Xbar.scala 256:54]
  wire  _T_2269 = ~_T_2189; // @[Xbar.scala 256:60]
  wire  _T_2270 = _T_2268 | _T_2269; // @[Xbar.scala 256:57]
  wire  _T_2271 = ~_T_2211; // @[Xbar.scala 256:54]
  wire  _T_2272 = ~_T_2190; // @[Xbar.scala 256:60]
  wire  _T_2273 = _T_2271 | _T_2272; // @[Xbar.scala 256:57]
  wire  _T_2274 = ~_T_2212; // @[Xbar.scala 256:54]
  wire  _T_2275 = ~_T_2191; // @[Xbar.scala 256:60]
  wire  _T_2276 = _T_2274 | _T_2275; // @[Xbar.scala 256:57]
  wire  _T_2278 = _T_2219 & _T_2222; // @[Xbar.scala 256:75]
  wire  _T_2279 = _T_2278 & _T_2225; // @[Xbar.scala 256:75]
  wire  _T_2280 = _T_2279 & _T_2228; // @[Xbar.scala 256:75]
  wire  _T_2281 = _T_2280 & _T_2231; // @[Xbar.scala 256:75]
  wire  _T_2282 = _T_2281 & _T_2234; // @[Xbar.scala 256:75]
  wire  _T_2283 = _T_2282 & _T_2237; // @[Xbar.scala 256:75]
  wire  _T_2284 = _T_2283 & _T_2240; // @[Xbar.scala 256:75]
  wire  _T_2285 = _T_2284 & _T_2243; // @[Xbar.scala 256:75]
  wire  _T_2286 = _T_2285 & _T_2246; // @[Xbar.scala 256:75]
  wire  _T_2287 = _T_2286 & _T_2249; // @[Xbar.scala 256:75]
  wire  _T_2288 = _T_2287 & _T_2252; // @[Xbar.scala 256:75]
  wire  _T_2289 = _T_2288 & _T_2255; // @[Xbar.scala 256:75]
  wire  _T_2290 = _T_2289 & _T_2258; // @[Xbar.scala 256:75]
  wire  _T_2291 = _T_2290 & _T_2261; // @[Xbar.scala 256:75]
  wire  _T_2292 = _T_2291 & _T_2264; // @[Xbar.scala 256:75]
  wire  _T_2293 = _T_2292 & _T_2267; // @[Xbar.scala 256:75]
  wire  _T_2294 = _T_2293 & _T_2270; // @[Xbar.scala 256:75]
  wire  _T_2295 = _T_2294 & _T_2273; // @[Xbar.scala 256:75]
  wire  _T_2296 = _T_2295 & _T_2276; // @[Xbar.scala 256:75]
  wire  _T_2298 = _T_2296 | reset; // @[Xbar.scala 256:11]
  wire  _T_2299 = ~_T_2298; // @[Xbar.scala 256:11]
  wire  _T_2300 = ~_T_2080; // @[Xbar.scala 258:13]
  wire  _T_2321 = _T_2300 | _T_2213; // @[Xbar.scala 258:23]
  wire  _T_2323 = _T_2321 | reset; // @[Xbar.scala 258:12]
  wire  _T_2324 = ~_T_2323; // @[Xbar.scala 258:12]
  wire  _T_2327_0 = _T_2060 ? _T_2171 : _T_2326_0; // @[Xbar.scala 262:23]
  wire  _T_2327_1 = _T_2060 ? _T_2172 : _T_2326_1; // @[Xbar.scala 262:23]
  wire  _T_2327_2 = _T_2060 ? _T_2173 : _T_2326_2; // @[Xbar.scala 262:23]
  wire  _T_2327_3 = _T_2060 ? _T_2174 : _T_2326_3; // @[Xbar.scala 262:23]
  wire  _T_2327_4 = _T_2060 ? _T_2175 : _T_2326_4; // @[Xbar.scala 262:23]
  wire  _T_2327_5 = _T_2060 ? _T_2176 : _T_2326_5; // @[Xbar.scala 262:23]
  wire  _T_2327_6 = _T_2060 ? _T_2177 : _T_2326_6; // @[Xbar.scala 262:23]
  wire  _T_2327_7 = _T_2060 ? _T_2178 : _T_2326_7; // @[Xbar.scala 262:23]
  wire  _T_2327_8 = _T_2060 ? _T_2179 : _T_2326_8; // @[Xbar.scala 262:23]
  wire  _T_2327_9 = _T_2060 ? _T_2180 : _T_2326_9; // @[Xbar.scala 262:23]
  wire  _T_2327_10 = _T_2060 ? _T_2181 : _T_2326_10; // @[Xbar.scala 262:23]
  wire  _T_2327_11 = _T_2060 ? _T_2182 : _T_2326_11; // @[Xbar.scala 262:23]
  wire  _T_2327_12 = _T_2060 ? _T_2183 : _T_2326_12; // @[Xbar.scala 262:23]
  wire  _T_2327_13 = _T_2060 ? _T_2184 : _T_2326_13; // @[Xbar.scala 262:23]
  wire  _T_2327_14 = _T_2060 ? _T_2185 : _T_2326_14; // @[Xbar.scala 262:23]
  wire  _T_2327_15 = _T_2060 ? _T_2186 : _T_2326_15; // @[Xbar.scala 262:23]
  wire  _T_2327_16 = _T_2060 ? _T_2187 : _T_2326_16; // @[Xbar.scala 262:23]
  wire  _T_2327_17 = _T_2060 ? _T_2188 : _T_2326_17; // @[Xbar.scala 262:23]
  wire  _T_2327_18 = _T_2060 ? _T_2189 : _T_2326_18; // @[Xbar.scala 262:23]
  wire  _T_2327_19 = _T_2060 ? _T_2190 : _T_2326_19; // @[Xbar.scala 262:23]
  wire  _T_2327_20 = _T_2060 ? _T_2191 : _T_2326_20; // @[Xbar.scala 262:23]
  wire  _GEN_92 = _T_2080 ? 1'h0 : _T_2060; // @[Xbar.scala 266:21]
  wire  _GEN_93 = _T_373 | _GEN_92; // @[Xbar.scala 267:24]
  wire  _T_2329_0 = _T_2060 ? _T_2128[0] : _T_2326_0; // @[Xbar.scala 270:24]
  wire  _T_2329_1 = _T_2060 ? _T_2128[1] : _T_2326_1; // @[Xbar.scala 270:24]
  wire  _T_2329_2 = _T_2060 ? _T_2128[2] : _T_2326_2; // @[Xbar.scala 270:24]
  wire  _T_2329_3 = _T_2060 ? _T_2128[3] : _T_2326_3; // @[Xbar.scala 270:24]
  wire  _T_2329_4 = _T_2060 ? _T_2128[4] : _T_2326_4; // @[Xbar.scala 270:24]
  wire  _T_2329_5 = _T_2060 ? _T_2128[5] : _T_2326_5; // @[Xbar.scala 270:24]
  wire  _T_2329_6 = _T_2060 ? _T_2128[6] : _T_2326_6; // @[Xbar.scala 270:24]
  wire  _T_2329_7 = _T_2060 ? _T_2128[7] : _T_2326_7; // @[Xbar.scala 270:24]
  wire  _T_2329_8 = _T_2060 ? _T_2128[8] : _T_2326_8; // @[Xbar.scala 270:24]
  wire  _T_2329_9 = _T_2060 ? _T_2128[9] : _T_2326_9; // @[Xbar.scala 270:24]
  wire  _T_2329_10 = _T_2060 ? _T_2128[10] : _T_2326_10; // @[Xbar.scala 270:24]
  wire  _T_2329_11 = _T_2060 ? _T_2128[11] : _T_2326_11; // @[Xbar.scala 270:24]
  wire  _T_2329_12 = _T_2060 ? _T_2128[12] : _T_2326_12; // @[Xbar.scala 270:24]
  wire  _T_2329_13 = _T_2060 ? _T_2128[13] : _T_2326_13; // @[Xbar.scala 270:24]
  wire  _T_2329_14 = _T_2060 ? _T_2128[14] : _T_2326_14; // @[Xbar.scala 270:24]
  wire  _T_2329_15 = _T_2060 ? _T_2128[15] : _T_2326_15; // @[Xbar.scala 270:24]
  wire  _T_2329_16 = _T_2060 ? _T_2128[16] : _T_2326_16; // @[Xbar.scala 270:24]
  wire  _T_2329_17 = _T_2060 ? _T_2128[17] : _T_2326_17; // @[Xbar.scala 270:24]
  wire  _T_2329_18 = _T_2060 ? _T_2128[18] : _T_2326_18; // @[Xbar.scala 270:24]
  wire  _T_2329_19 = _T_2060 ? _T_2128[19] : _T_2326_19; // @[Xbar.scala 270:24]
  wire  _T_2329_20 = _T_2060 ? _T_2128[20] : _T_2326_20; // @[Xbar.scala 270:24]
  wire [2:0] _T_2394 = {auto_out_0_b_bits_id,auto_out_0_b_bits_resp}; // @[Mux.scala 27:72]
  wire [2:0] _T_2395 = _T_2327_0 ? _T_2394 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_2396 = {auto_out_1_b_bits_id,auto_out_1_b_bits_resp}; // @[Mux.scala 27:72]
  wire [2:0] _T_2397 = _T_2327_1 ? _T_2396 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_2398 = {auto_out_2_b_bits_id,auto_out_2_b_bits_resp}; // @[Mux.scala 27:72]
  wire [2:0] _T_2399 = _T_2327_2 ? _T_2398 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_2400 = {auto_out_3_b_bits_id,auto_out_3_b_bits_resp}; // @[Mux.scala 27:72]
  wire [2:0] _T_2401 = _T_2327_3 ? _T_2400 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_2402 = {auto_out_4_b_bits_id,auto_out_4_b_bits_resp}; // @[Mux.scala 27:72]
  wire [2:0] _T_2403 = _T_2327_4 ? _T_2402 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_2404 = {auto_out_5_b_bits_id,auto_out_5_b_bits_resp}; // @[Mux.scala 27:72]
  wire [2:0] _T_2405 = _T_2327_5 ? _T_2404 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_2406 = {auto_out_6_b_bits_id,auto_out_6_b_bits_resp}; // @[Mux.scala 27:72]
  wire [2:0] _T_2407 = _T_2327_6 ? _T_2406 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_2408 = {auto_out_7_b_bits_id,auto_out_7_b_bits_resp}; // @[Mux.scala 27:72]
  wire [2:0] _T_2409 = _T_2327_7 ? _T_2408 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_2410 = {auto_out_8_b_bits_id,auto_out_8_b_bits_resp}; // @[Mux.scala 27:72]
  wire [2:0] _T_2411 = _T_2327_8 ? _T_2410 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_2412 = {auto_out_9_b_bits_id,auto_out_9_b_bits_resp}; // @[Mux.scala 27:72]
  wire [2:0] _T_2413 = _T_2327_9 ? _T_2412 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_2414 = {auto_out_10_b_bits_id,auto_out_10_b_bits_resp}; // @[Mux.scala 27:72]
  wire [2:0] _T_2415 = _T_2327_10 ? _T_2414 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_2416 = {auto_out_11_b_bits_id,auto_out_11_b_bits_resp}; // @[Mux.scala 27:72]
  wire [2:0] _T_2417 = _T_2327_11 ? _T_2416 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_2418 = {auto_out_12_b_bits_id,auto_out_12_b_bits_resp}; // @[Mux.scala 27:72]
  wire [2:0] _T_2419 = _T_2327_12 ? _T_2418 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_2420 = {auto_out_13_b_bits_id,auto_out_13_b_bits_resp}; // @[Mux.scala 27:72]
  wire [2:0] _T_2421 = _T_2327_13 ? _T_2420 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_2422 = {auto_out_14_b_bits_id,auto_out_14_b_bits_resp}; // @[Mux.scala 27:72]
  wire [2:0] _T_2423 = _T_2327_14 ? _T_2422 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_2424 = {auto_out_15_b_bits_id,auto_out_15_b_bits_resp}; // @[Mux.scala 27:72]
  wire [2:0] _T_2425 = _T_2327_15 ? _T_2424 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_2426 = {auto_out_16_b_bits_id,auto_out_16_b_bits_resp}; // @[Mux.scala 27:72]
  wire [2:0] _T_2427 = _T_2327_16 ? _T_2426 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_2428 = {auto_out_17_b_bits_id,auto_out_17_b_bits_resp}; // @[Mux.scala 27:72]
  wire [2:0] _T_2429 = _T_2327_17 ? _T_2428 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_2430 = {auto_out_18_b_bits_id,auto_out_18_b_bits_resp}; // @[Mux.scala 27:72]
  wire [2:0] _T_2431 = _T_2327_18 ? _T_2430 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_2432 = {auto_out_19_b_bits_id,auto_out_19_b_bits_resp}; // @[Mux.scala 27:72]
  wire [2:0] _T_2433 = _T_2327_19 ? _T_2432 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_2434 = {1'h0,auto_out_20_b_bits_resp}; // @[Mux.scala 27:72]
  wire [2:0] _T_2435 = _T_2327_20 ? _T_2434 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_2436 = _T_2395 | _T_2397; // @[Mux.scala 27:72]
  wire [2:0] _T_2437 = _T_2436 | _T_2399; // @[Mux.scala 27:72]
  wire [2:0] _T_2438 = _T_2437 | _T_2401; // @[Mux.scala 27:72]
  wire [2:0] _T_2439 = _T_2438 | _T_2403; // @[Mux.scala 27:72]
  wire [2:0] _T_2440 = _T_2439 | _T_2405; // @[Mux.scala 27:72]
  wire [2:0] _T_2441 = _T_2440 | _T_2407; // @[Mux.scala 27:72]
  wire [2:0] _T_2442 = _T_2441 | _T_2409; // @[Mux.scala 27:72]
  wire [2:0] _T_2443 = _T_2442 | _T_2411; // @[Mux.scala 27:72]
  wire [2:0] _T_2444 = _T_2443 | _T_2413; // @[Mux.scala 27:72]
  wire [2:0] _T_2445 = _T_2444 | _T_2415; // @[Mux.scala 27:72]
  wire [2:0] _T_2446 = _T_2445 | _T_2417; // @[Mux.scala 27:72]
  wire [2:0] _T_2447 = _T_2446 | _T_2419; // @[Mux.scala 27:72]
  wire [2:0] _T_2448 = _T_2447 | _T_2421; // @[Mux.scala 27:72]
  wire [2:0] _T_2449 = _T_2448 | _T_2423; // @[Mux.scala 27:72]
  wire [2:0] _T_2450 = _T_2449 | _T_2425; // @[Mux.scala 27:72]
  wire [2:0] _T_2451 = _T_2450 | _T_2427; // @[Mux.scala 27:72]
  wire [2:0] _T_2452 = _T_2451 | _T_2429; // @[Mux.scala 27:72]
  wire [2:0] _T_2453 = _T_2452 | _T_2431; // @[Mux.scala 27:72]
  wire [2:0] _T_2454 = _T_2453 | _T_2433; // @[Mux.scala 27:72]
  wire [2:0] _T_2455 = _T_2454 | _T_2435; // @[Mux.scala 27:72]
  QueueCompatibility_8 awIn_0 ( // @[Xbar.scala 55:47]
    .clock(awIn_0_clock),
    .reset(awIn_0_reset),
    .io_enq_ready(awIn_0_io_enq_ready),
    .io_enq_valid(awIn_0_io_enq_valid),
    .io_enq_bits(awIn_0_io_enq_bits),
    .io_deq_ready(awIn_0_io_deq_ready),
    .io_deq_valid(awIn_0_io_deq_valid),
    .io_deq_bits(awIn_0_io_deq_bits)
  );
  assign auto_in_aw_ready = _T_406 & _T_398; // @[LazyModule.scala 173:31]
  assign auto_in_w_ready = in_0_w_ready & awIn_0_io_deq_valid; // @[LazyModule.scala 173:31]
  assign auto_in_b_valid = _T_2060 ? _T_2080 : _T_2391; // @[LazyModule.scala 173:31]
  assign auto_in_b_bits_resp = _T_2455[1:0]; // @[LazyModule.scala 173:31]
  assign auto_in_ar_ready = in_0_ar_ready & _T_370; // @[LazyModule.scala 173:31]
  assign auto_in_r_valid = _T_1616 ? _T_1636 : _T_1947; // @[LazyModule.scala 173:31]
  assign auto_in_r_bits_data = _T_2053[34:3]; // @[LazyModule.scala 173:31]
  assign auto_in_r_bits_resp = _T_2053[2:1]; // @[LazyModule.scala 173:31]
  assign auto_in_r_bits_last = _T_2053[0]; // @[LazyModule.scala 173:31]
  assign auto_out_20_aw_valid = in_0_aw_valid & requestAWIO_0_20; // @[LazyModule.scala 173:49]
  assign auto_out_20_aw_bits_id = auto_in_aw_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_20_aw_bits_addr = auto_in_aw_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_20_aw_bits_size = auto_in_aw_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_20_w_valid = in_0_w_valid & requestWIO_0_20; // @[LazyModule.scala 173:49]
  assign auto_out_20_w_bits_data = auto_in_w_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_20_w_bits_strb = auto_in_w_bits_strb; // @[LazyModule.scala 173:49]
  assign auto_out_20_w_bits_last = auto_in_w_bits_last; // @[LazyModule.scala 173:49]
  assign auto_out_20_b_ready = auto_in_b_ready & _T_2329_20; // @[LazyModule.scala 173:49]
  assign auto_out_20_ar_valid = in_0_ar_valid & requestARIO_0_20; // @[LazyModule.scala 173:49]
  assign auto_out_20_ar_bits_id = auto_in_ar_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_20_ar_bits_addr = auto_in_ar_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_20_ar_bits_size = auto_in_ar_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_20_r_ready = auto_in_r_ready & _T_1885_20; // @[LazyModule.scala 173:49]
  assign auto_out_19_aw_valid = in_0_aw_valid & requestAWIO_0_19; // @[LazyModule.scala 173:49]
  assign auto_out_19_aw_bits_id = auto_in_aw_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_19_aw_bits_addr = auto_in_aw_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_19_aw_bits_size = auto_in_aw_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_19_w_valid = in_0_w_valid & requestWIO_0_19; // @[LazyModule.scala 173:49]
  assign auto_out_19_w_bits_data = auto_in_w_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_19_w_bits_strb = auto_in_w_bits_strb; // @[LazyModule.scala 173:49]
  assign auto_out_19_w_bits_last = auto_in_w_bits_last; // @[LazyModule.scala 173:49]
  assign auto_out_19_b_ready = auto_in_b_ready & _T_2329_19; // @[LazyModule.scala 173:49]
  assign auto_out_19_ar_valid = in_0_ar_valid & requestARIO_0_19; // @[LazyModule.scala 173:49]
  assign auto_out_19_ar_bits_id = auto_in_ar_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_19_ar_bits_addr = auto_in_ar_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_19_ar_bits_size = auto_in_ar_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_19_r_ready = auto_in_r_ready & _T_1885_19; // @[LazyModule.scala 173:49]
  assign auto_out_18_aw_valid = in_0_aw_valid & requestAWIO_0_18; // @[LazyModule.scala 173:49]
  assign auto_out_18_aw_bits_id = auto_in_aw_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_18_aw_bits_addr = auto_in_aw_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_18_aw_bits_size = auto_in_aw_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_18_w_valid = in_0_w_valid & requestWIO_0_18; // @[LazyModule.scala 173:49]
  assign auto_out_18_w_bits_data = auto_in_w_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_18_w_bits_strb = auto_in_w_bits_strb; // @[LazyModule.scala 173:49]
  assign auto_out_18_w_bits_last = auto_in_w_bits_last; // @[LazyModule.scala 173:49]
  assign auto_out_18_b_ready = auto_in_b_ready & _T_2329_18; // @[LazyModule.scala 173:49]
  assign auto_out_18_ar_valid = in_0_ar_valid & requestARIO_0_18; // @[LazyModule.scala 173:49]
  assign auto_out_18_ar_bits_id = auto_in_ar_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_18_ar_bits_addr = auto_in_ar_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_18_ar_bits_size = auto_in_ar_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_18_r_ready = auto_in_r_ready & _T_1885_18; // @[LazyModule.scala 173:49]
  assign auto_out_17_aw_valid = in_0_aw_valid & requestAWIO_0_17; // @[LazyModule.scala 173:49]
  assign auto_out_17_aw_bits_id = auto_in_aw_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_17_aw_bits_addr = auto_in_aw_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_17_aw_bits_size = auto_in_aw_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_17_w_valid = in_0_w_valid & requestWIO_0_17; // @[LazyModule.scala 173:49]
  assign auto_out_17_w_bits_data = auto_in_w_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_17_w_bits_strb = auto_in_w_bits_strb; // @[LazyModule.scala 173:49]
  assign auto_out_17_w_bits_last = auto_in_w_bits_last; // @[LazyModule.scala 173:49]
  assign auto_out_17_b_ready = auto_in_b_ready & _T_2329_17; // @[LazyModule.scala 173:49]
  assign auto_out_17_ar_valid = in_0_ar_valid & requestARIO_0_17; // @[LazyModule.scala 173:49]
  assign auto_out_17_ar_bits_id = auto_in_ar_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_17_ar_bits_addr = auto_in_ar_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_17_ar_bits_size = auto_in_ar_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_17_r_ready = auto_in_r_ready & _T_1885_17; // @[LazyModule.scala 173:49]
  assign auto_out_16_aw_valid = in_0_aw_valid & requestAWIO_0_16; // @[LazyModule.scala 173:49]
  assign auto_out_16_aw_bits_id = auto_in_aw_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_16_aw_bits_addr = auto_in_aw_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_16_aw_bits_size = auto_in_aw_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_16_w_valid = in_0_w_valid & requestWIO_0_16; // @[LazyModule.scala 173:49]
  assign auto_out_16_w_bits_data = auto_in_w_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_16_w_bits_strb = auto_in_w_bits_strb; // @[LazyModule.scala 173:49]
  assign auto_out_16_w_bits_last = auto_in_w_bits_last; // @[LazyModule.scala 173:49]
  assign auto_out_16_b_ready = auto_in_b_ready & _T_2329_16; // @[LazyModule.scala 173:49]
  assign auto_out_16_ar_valid = in_0_ar_valid & requestARIO_0_16; // @[LazyModule.scala 173:49]
  assign auto_out_16_ar_bits_id = auto_in_ar_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_16_ar_bits_addr = auto_in_ar_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_16_ar_bits_size = auto_in_ar_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_16_r_ready = auto_in_r_ready & _T_1885_16; // @[LazyModule.scala 173:49]
  assign auto_out_15_aw_valid = in_0_aw_valid & requestAWIO_0_15; // @[LazyModule.scala 173:49]
  assign auto_out_15_aw_bits_id = auto_in_aw_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_15_aw_bits_addr = auto_in_aw_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_15_aw_bits_size = auto_in_aw_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_15_w_valid = in_0_w_valid & requestWIO_0_15; // @[LazyModule.scala 173:49]
  assign auto_out_15_w_bits_data = auto_in_w_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_15_w_bits_strb = auto_in_w_bits_strb; // @[LazyModule.scala 173:49]
  assign auto_out_15_w_bits_last = auto_in_w_bits_last; // @[LazyModule.scala 173:49]
  assign auto_out_15_b_ready = auto_in_b_ready & _T_2329_15; // @[LazyModule.scala 173:49]
  assign auto_out_15_ar_valid = in_0_ar_valid & requestARIO_0_15; // @[LazyModule.scala 173:49]
  assign auto_out_15_ar_bits_id = auto_in_ar_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_15_ar_bits_addr = auto_in_ar_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_15_ar_bits_size = auto_in_ar_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_15_r_ready = auto_in_r_ready & _T_1885_15; // @[LazyModule.scala 173:49]
  assign auto_out_14_aw_valid = in_0_aw_valid & requestAWIO_0_14; // @[LazyModule.scala 173:49]
  assign auto_out_14_aw_bits_id = auto_in_aw_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_14_aw_bits_addr = auto_in_aw_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_14_aw_bits_size = auto_in_aw_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_14_w_valid = in_0_w_valid & requestWIO_0_14; // @[LazyModule.scala 173:49]
  assign auto_out_14_w_bits_data = auto_in_w_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_14_w_bits_strb = auto_in_w_bits_strb; // @[LazyModule.scala 173:49]
  assign auto_out_14_w_bits_last = auto_in_w_bits_last; // @[LazyModule.scala 173:49]
  assign auto_out_14_b_ready = auto_in_b_ready & _T_2329_14; // @[LazyModule.scala 173:49]
  assign auto_out_14_ar_valid = in_0_ar_valid & requestARIO_0_14; // @[LazyModule.scala 173:49]
  assign auto_out_14_ar_bits_id = auto_in_ar_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_14_ar_bits_addr = auto_in_ar_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_14_ar_bits_size = auto_in_ar_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_14_r_ready = auto_in_r_ready & _T_1885_14; // @[LazyModule.scala 173:49]
  assign auto_out_13_aw_valid = in_0_aw_valid & requestAWIO_0_13; // @[LazyModule.scala 173:49]
  assign auto_out_13_aw_bits_id = auto_in_aw_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_13_aw_bits_addr = auto_in_aw_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_13_aw_bits_size = auto_in_aw_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_13_w_valid = in_0_w_valid & requestWIO_0_13; // @[LazyModule.scala 173:49]
  assign auto_out_13_w_bits_data = auto_in_w_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_13_w_bits_strb = auto_in_w_bits_strb; // @[LazyModule.scala 173:49]
  assign auto_out_13_w_bits_last = auto_in_w_bits_last; // @[LazyModule.scala 173:49]
  assign auto_out_13_b_ready = auto_in_b_ready & _T_2329_13; // @[LazyModule.scala 173:49]
  assign auto_out_13_ar_valid = in_0_ar_valid & requestARIO_0_13; // @[LazyModule.scala 173:49]
  assign auto_out_13_ar_bits_id = auto_in_ar_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_13_ar_bits_addr = auto_in_ar_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_13_ar_bits_size = auto_in_ar_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_13_r_ready = auto_in_r_ready & _T_1885_13; // @[LazyModule.scala 173:49]
  assign auto_out_12_aw_valid = in_0_aw_valid & requestAWIO_0_12; // @[LazyModule.scala 173:49]
  assign auto_out_12_aw_bits_id = auto_in_aw_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_12_aw_bits_addr = auto_in_aw_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_12_aw_bits_size = auto_in_aw_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_12_w_valid = in_0_w_valid & requestWIO_0_12; // @[LazyModule.scala 173:49]
  assign auto_out_12_w_bits_data = auto_in_w_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_12_w_bits_strb = auto_in_w_bits_strb; // @[LazyModule.scala 173:49]
  assign auto_out_12_w_bits_last = auto_in_w_bits_last; // @[LazyModule.scala 173:49]
  assign auto_out_12_b_ready = auto_in_b_ready & _T_2329_12; // @[LazyModule.scala 173:49]
  assign auto_out_12_ar_valid = in_0_ar_valid & requestARIO_0_12; // @[LazyModule.scala 173:49]
  assign auto_out_12_ar_bits_id = auto_in_ar_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_12_ar_bits_addr = auto_in_ar_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_12_ar_bits_size = auto_in_ar_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_12_r_ready = auto_in_r_ready & _T_1885_12; // @[LazyModule.scala 173:49]
  assign auto_out_11_aw_valid = in_0_aw_valid & requestAWIO_0_11; // @[LazyModule.scala 173:49]
  assign auto_out_11_aw_bits_id = auto_in_aw_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_11_aw_bits_addr = auto_in_aw_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_11_aw_bits_size = auto_in_aw_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_11_w_valid = in_0_w_valid & requestWIO_0_11; // @[LazyModule.scala 173:49]
  assign auto_out_11_w_bits_data = auto_in_w_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_11_w_bits_strb = auto_in_w_bits_strb; // @[LazyModule.scala 173:49]
  assign auto_out_11_w_bits_last = auto_in_w_bits_last; // @[LazyModule.scala 173:49]
  assign auto_out_11_b_ready = auto_in_b_ready & _T_2329_11; // @[LazyModule.scala 173:49]
  assign auto_out_11_ar_valid = in_0_ar_valid & requestARIO_0_11; // @[LazyModule.scala 173:49]
  assign auto_out_11_ar_bits_id = auto_in_ar_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_11_ar_bits_addr = auto_in_ar_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_11_ar_bits_size = auto_in_ar_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_11_r_ready = auto_in_r_ready & _T_1885_11; // @[LazyModule.scala 173:49]
  assign auto_out_10_aw_valid = in_0_aw_valid & requestAWIO_0_10; // @[LazyModule.scala 173:49]
  assign auto_out_10_aw_bits_id = auto_in_aw_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_10_aw_bits_addr = auto_in_aw_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_10_aw_bits_size = auto_in_aw_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_10_w_valid = in_0_w_valid & requestWIO_0_10; // @[LazyModule.scala 173:49]
  assign auto_out_10_w_bits_data = auto_in_w_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_10_w_bits_strb = auto_in_w_bits_strb; // @[LazyModule.scala 173:49]
  assign auto_out_10_w_bits_last = auto_in_w_bits_last; // @[LazyModule.scala 173:49]
  assign auto_out_10_b_ready = auto_in_b_ready & _T_2329_10; // @[LazyModule.scala 173:49]
  assign auto_out_10_ar_valid = in_0_ar_valid & requestARIO_0_10; // @[LazyModule.scala 173:49]
  assign auto_out_10_ar_bits_id = auto_in_ar_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_10_ar_bits_addr = auto_in_ar_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_10_ar_bits_size = auto_in_ar_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_10_r_ready = auto_in_r_ready & _T_1885_10; // @[LazyModule.scala 173:49]
  assign auto_out_9_aw_valid = in_0_aw_valid & requestAWIO_0_9; // @[LazyModule.scala 173:49]
  assign auto_out_9_aw_bits_id = auto_in_aw_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_9_aw_bits_addr = auto_in_aw_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_9_aw_bits_size = auto_in_aw_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_9_w_valid = in_0_w_valid & requestWIO_0_9; // @[LazyModule.scala 173:49]
  assign auto_out_9_w_bits_data = auto_in_w_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_9_w_bits_strb = auto_in_w_bits_strb; // @[LazyModule.scala 173:49]
  assign auto_out_9_w_bits_last = auto_in_w_bits_last; // @[LazyModule.scala 173:49]
  assign auto_out_9_b_ready = auto_in_b_ready & _T_2329_9; // @[LazyModule.scala 173:49]
  assign auto_out_9_ar_valid = in_0_ar_valid & requestARIO_0_9; // @[LazyModule.scala 173:49]
  assign auto_out_9_ar_bits_id = auto_in_ar_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_9_ar_bits_addr = auto_in_ar_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_9_ar_bits_size = auto_in_ar_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_9_r_ready = auto_in_r_ready & _T_1885_9; // @[LazyModule.scala 173:49]
  assign auto_out_8_aw_valid = in_0_aw_valid & requestAWIO_0_8; // @[LazyModule.scala 173:49]
  assign auto_out_8_aw_bits_id = auto_in_aw_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_8_aw_bits_addr = auto_in_aw_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_8_aw_bits_size = auto_in_aw_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_8_w_valid = in_0_w_valid & requestWIO_0_8; // @[LazyModule.scala 173:49]
  assign auto_out_8_w_bits_data = auto_in_w_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_8_w_bits_strb = auto_in_w_bits_strb; // @[LazyModule.scala 173:49]
  assign auto_out_8_w_bits_last = auto_in_w_bits_last; // @[LazyModule.scala 173:49]
  assign auto_out_8_b_ready = auto_in_b_ready & _T_2329_8; // @[LazyModule.scala 173:49]
  assign auto_out_8_ar_valid = in_0_ar_valid & requestARIO_0_8; // @[LazyModule.scala 173:49]
  assign auto_out_8_ar_bits_id = auto_in_ar_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_8_ar_bits_addr = auto_in_ar_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_8_ar_bits_size = auto_in_ar_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_8_r_ready = auto_in_r_ready & _T_1885_8; // @[LazyModule.scala 173:49]
  assign auto_out_7_aw_valid = in_0_aw_valid & requestAWIO_0_7; // @[LazyModule.scala 173:49]
  assign auto_out_7_aw_bits_id = auto_in_aw_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_7_aw_bits_addr = auto_in_aw_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_7_aw_bits_size = auto_in_aw_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_7_w_valid = in_0_w_valid & requestWIO_0_7; // @[LazyModule.scala 173:49]
  assign auto_out_7_w_bits_data = auto_in_w_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_7_w_bits_strb = auto_in_w_bits_strb; // @[LazyModule.scala 173:49]
  assign auto_out_7_w_bits_last = auto_in_w_bits_last; // @[LazyModule.scala 173:49]
  assign auto_out_7_b_ready = auto_in_b_ready & _T_2329_7; // @[LazyModule.scala 173:49]
  assign auto_out_7_ar_valid = in_0_ar_valid & requestARIO_0_7; // @[LazyModule.scala 173:49]
  assign auto_out_7_ar_bits_id = auto_in_ar_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_7_ar_bits_addr = auto_in_ar_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_7_ar_bits_size = auto_in_ar_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_7_r_ready = auto_in_r_ready & _T_1885_7; // @[LazyModule.scala 173:49]
  assign auto_out_6_aw_valid = in_0_aw_valid & requestAWIO_0_6; // @[LazyModule.scala 173:49]
  assign auto_out_6_aw_bits_id = auto_in_aw_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_6_aw_bits_addr = auto_in_aw_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_6_aw_bits_size = auto_in_aw_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_6_w_valid = in_0_w_valid & requestWIO_0_6; // @[LazyModule.scala 173:49]
  assign auto_out_6_w_bits_data = auto_in_w_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_6_w_bits_strb = auto_in_w_bits_strb; // @[LazyModule.scala 173:49]
  assign auto_out_6_w_bits_last = auto_in_w_bits_last; // @[LazyModule.scala 173:49]
  assign auto_out_6_b_ready = auto_in_b_ready & _T_2329_6; // @[LazyModule.scala 173:49]
  assign auto_out_6_ar_valid = in_0_ar_valid & requestARIO_0_6; // @[LazyModule.scala 173:49]
  assign auto_out_6_ar_bits_id = auto_in_ar_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_6_ar_bits_addr = auto_in_ar_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_6_ar_bits_size = auto_in_ar_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_6_r_ready = auto_in_r_ready & _T_1885_6; // @[LazyModule.scala 173:49]
  assign auto_out_5_aw_valid = in_0_aw_valid & requestAWIO_0_5; // @[LazyModule.scala 173:49]
  assign auto_out_5_aw_bits_id = auto_in_aw_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_5_aw_bits_addr = auto_in_aw_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_5_aw_bits_size = auto_in_aw_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_5_w_valid = in_0_w_valid & requestWIO_0_5; // @[LazyModule.scala 173:49]
  assign auto_out_5_w_bits_data = auto_in_w_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_5_w_bits_strb = auto_in_w_bits_strb; // @[LazyModule.scala 173:49]
  assign auto_out_5_w_bits_last = auto_in_w_bits_last; // @[LazyModule.scala 173:49]
  assign auto_out_5_b_ready = auto_in_b_ready & _T_2329_5; // @[LazyModule.scala 173:49]
  assign auto_out_5_ar_valid = in_0_ar_valid & requestARIO_0_5; // @[LazyModule.scala 173:49]
  assign auto_out_5_ar_bits_id = auto_in_ar_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_5_ar_bits_addr = auto_in_ar_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_5_ar_bits_size = auto_in_ar_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_5_r_ready = auto_in_r_ready & _T_1885_5; // @[LazyModule.scala 173:49]
  assign auto_out_4_aw_valid = in_0_aw_valid & requestAWIO_0_4; // @[LazyModule.scala 173:49]
  assign auto_out_4_aw_bits_id = auto_in_aw_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_4_aw_bits_addr = auto_in_aw_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_4_aw_bits_size = auto_in_aw_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_4_w_valid = in_0_w_valid & requestWIO_0_4; // @[LazyModule.scala 173:49]
  assign auto_out_4_w_bits_data = auto_in_w_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_4_w_bits_strb = auto_in_w_bits_strb; // @[LazyModule.scala 173:49]
  assign auto_out_4_w_bits_last = auto_in_w_bits_last; // @[LazyModule.scala 173:49]
  assign auto_out_4_b_ready = auto_in_b_ready & _T_2329_4; // @[LazyModule.scala 173:49]
  assign auto_out_4_ar_valid = in_0_ar_valid & requestARIO_0_4; // @[LazyModule.scala 173:49]
  assign auto_out_4_ar_bits_id = auto_in_ar_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_4_ar_bits_addr = auto_in_ar_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_4_ar_bits_size = auto_in_ar_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_4_r_ready = auto_in_r_ready & _T_1885_4; // @[LazyModule.scala 173:49]
  assign auto_out_3_aw_valid = in_0_aw_valid & requestAWIO_0_3; // @[LazyModule.scala 173:49]
  assign auto_out_3_aw_bits_id = auto_in_aw_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_3_aw_bits_addr = auto_in_aw_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_3_aw_bits_size = auto_in_aw_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_3_w_valid = in_0_w_valid & requestWIO_0_3; // @[LazyModule.scala 173:49]
  assign auto_out_3_w_bits_data = auto_in_w_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_3_w_bits_strb = auto_in_w_bits_strb; // @[LazyModule.scala 173:49]
  assign auto_out_3_w_bits_last = auto_in_w_bits_last; // @[LazyModule.scala 173:49]
  assign auto_out_3_b_ready = auto_in_b_ready & _T_2329_3; // @[LazyModule.scala 173:49]
  assign auto_out_3_ar_valid = in_0_ar_valid & requestARIO_0_3; // @[LazyModule.scala 173:49]
  assign auto_out_3_ar_bits_id = auto_in_ar_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_3_ar_bits_addr = auto_in_ar_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_3_ar_bits_size = auto_in_ar_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_3_r_ready = auto_in_r_ready & _T_1885_3; // @[LazyModule.scala 173:49]
  assign auto_out_2_aw_valid = in_0_aw_valid & requestAWIO_0_2; // @[LazyModule.scala 173:49]
  assign auto_out_2_aw_bits_id = auto_in_aw_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_2_aw_bits_addr = auto_in_aw_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_2_aw_bits_size = auto_in_aw_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_2_w_valid = in_0_w_valid & requestWIO_0_2; // @[LazyModule.scala 173:49]
  assign auto_out_2_w_bits_data = auto_in_w_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_2_w_bits_strb = auto_in_w_bits_strb; // @[LazyModule.scala 173:49]
  assign auto_out_2_w_bits_last = auto_in_w_bits_last; // @[LazyModule.scala 173:49]
  assign auto_out_2_b_ready = auto_in_b_ready & _T_2329_2; // @[LazyModule.scala 173:49]
  assign auto_out_2_ar_valid = in_0_ar_valid & requestARIO_0_2; // @[LazyModule.scala 173:49]
  assign auto_out_2_ar_bits_id = auto_in_ar_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_2_ar_bits_addr = auto_in_ar_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_2_ar_bits_size = auto_in_ar_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_2_r_ready = auto_in_r_ready & _T_1885_2; // @[LazyModule.scala 173:49]
  assign auto_out_1_aw_valid = in_0_aw_valid & requestAWIO_0_1; // @[LazyModule.scala 173:49]
  assign auto_out_1_aw_bits_id = auto_in_aw_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_1_aw_bits_addr = auto_in_aw_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_1_aw_bits_size = auto_in_aw_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_1_w_valid = in_0_w_valid & requestWIO_0_1; // @[LazyModule.scala 173:49]
  assign auto_out_1_w_bits_data = auto_in_w_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_1_w_bits_strb = auto_in_w_bits_strb; // @[LazyModule.scala 173:49]
  assign auto_out_1_w_bits_last = auto_in_w_bits_last; // @[LazyModule.scala 173:49]
  assign auto_out_1_b_ready = auto_in_b_ready & _T_2329_1; // @[LazyModule.scala 173:49]
  assign auto_out_1_ar_valid = in_0_ar_valid & requestARIO_0_1; // @[LazyModule.scala 173:49]
  assign auto_out_1_ar_bits_id = auto_in_ar_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_1_ar_bits_addr = auto_in_ar_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_1_ar_bits_size = auto_in_ar_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_1_r_ready = auto_in_r_ready & _T_1885_1; // @[LazyModule.scala 173:49]
  assign auto_out_0_aw_valid = in_0_aw_valid & requestAWIO_0_0; // @[LazyModule.scala 173:49]
  assign auto_out_0_aw_bits_id = auto_in_aw_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_0_aw_bits_addr = auto_in_aw_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_0_aw_bits_size = auto_in_aw_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_0_w_valid = in_0_w_valid & requestWIO_0_0; // @[LazyModule.scala 173:49]
  assign auto_out_0_w_bits_data = auto_in_w_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_0_w_bits_strb = auto_in_w_bits_strb; // @[LazyModule.scala 173:49]
  assign auto_out_0_w_bits_last = auto_in_w_bits_last; // @[LazyModule.scala 173:49]
  assign auto_out_0_b_ready = auto_in_b_ready & _T_2329_0; // @[LazyModule.scala 173:49]
  assign auto_out_0_ar_valid = in_0_ar_valid & requestARIO_0_0; // @[LazyModule.scala 173:49]
  assign auto_out_0_ar_bits_id = auto_in_ar_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_0_ar_bits_addr = auto_in_ar_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_0_ar_bits_size = auto_in_ar_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_0_r_ready = auto_in_r_ready & _T_1885_0; // @[LazyModule.scala 173:49]
  assign awIn_0_clock = clock;
  assign awIn_0_reset = reset;
  assign awIn_0_io_enq_valid = auto_in_aw_valid & _T_408; // @[Xbar.scala 140:30]
  assign awIn_0_io_enq_bits = {_T_252,_T_242}; // @[Xbar.scala 64:57]
  assign awIn_0_io_deq_ready = _T_414 & in_0_w_ready; // @[Xbar.scala 147:30]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_347 = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_348 = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_1616 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_1882_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_1882_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_1882_2 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_1882_3 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_1882_4 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_1882_5 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_1882_6 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_1882_7 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_1882_8 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_1882_9 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_1882_10 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_1882_11 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_1882_12 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_1882_13 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_1882_14 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_1882_15 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_1882_16 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_1882_17 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_1882_18 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_1882_19 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_1882_20 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_1663 = _RAND_24[20:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_401 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_375 = _RAND_26[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T_376 = _RAND_27[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_2060 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_2326_0 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_2326_1 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T_2326_2 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _T_2326_3 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _T_2326_4 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _T_2326_5 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _T_2326_6 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _T_2326_7 = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _T_2326_8 = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _T_2326_9 = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _T_2326_10 = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _T_2326_11 = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  _T_2326_12 = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  _T_2326_13 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  _T_2326_14 = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  _T_2326_15 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  _T_2326_16 = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  _T_2326_17 = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  _T_2326_18 = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  _T_2326_19 = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  _T_2326_20 = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  _T_2107 = _RAND_50[20:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      _T_347 <= 3'h0;
    end else begin
      _T_347 <= _T_352;
    end
    if (_T_342) begin
      _T_348 <= _T_300;
    end
    _T_1616 <= reset | _GEN_90;
    if (reset) begin
      _T_1882_0 <= 1'h0;
    end else if (_T_1616) begin
      _T_1882_0 <= _T_1727;
    end
    if (reset) begin
      _T_1882_1 <= 1'h0;
    end else if (_T_1616) begin
      _T_1882_1 <= _T_1728;
    end
    if (reset) begin
      _T_1882_2 <= 1'h0;
    end else if (_T_1616) begin
      _T_1882_2 <= _T_1729;
    end
    if (reset) begin
      _T_1882_3 <= 1'h0;
    end else if (_T_1616) begin
      _T_1882_3 <= _T_1730;
    end
    if (reset) begin
      _T_1882_4 <= 1'h0;
    end else if (_T_1616) begin
      _T_1882_4 <= _T_1731;
    end
    if (reset) begin
      _T_1882_5 <= 1'h0;
    end else if (_T_1616) begin
      _T_1882_5 <= _T_1732;
    end
    if (reset) begin
      _T_1882_6 <= 1'h0;
    end else if (_T_1616) begin
      _T_1882_6 <= _T_1733;
    end
    if (reset) begin
      _T_1882_7 <= 1'h0;
    end else if (_T_1616) begin
      _T_1882_7 <= _T_1734;
    end
    if (reset) begin
      _T_1882_8 <= 1'h0;
    end else if (_T_1616) begin
      _T_1882_8 <= _T_1735;
    end
    if (reset) begin
      _T_1882_9 <= 1'h0;
    end else if (_T_1616) begin
      _T_1882_9 <= _T_1736;
    end
    if (reset) begin
      _T_1882_10 <= 1'h0;
    end else if (_T_1616) begin
      _T_1882_10 <= _T_1737;
    end
    if (reset) begin
      _T_1882_11 <= 1'h0;
    end else if (_T_1616) begin
      _T_1882_11 <= _T_1738;
    end
    if (reset) begin
      _T_1882_12 <= 1'h0;
    end else if (_T_1616) begin
      _T_1882_12 <= _T_1739;
    end
    if (reset) begin
      _T_1882_13 <= 1'h0;
    end else if (_T_1616) begin
      _T_1882_13 <= _T_1740;
    end
    if (reset) begin
      _T_1882_14 <= 1'h0;
    end else if (_T_1616) begin
      _T_1882_14 <= _T_1741;
    end
    if (reset) begin
      _T_1882_15 <= 1'h0;
    end else if (_T_1616) begin
      _T_1882_15 <= _T_1742;
    end
    if (reset) begin
      _T_1882_16 <= 1'h0;
    end else if (_T_1616) begin
      _T_1882_16 <= _T_1743;
    end
    if (reset) begin
      _T_1882_17 <= 1'h0;
    end else if (_T_1616) begin
      _T_1882_17 <= _T_1744;
    end
    if (reset) begin
      _T_1882_18 <= 1'h0;
    end else if (_T_1616) begin
      _T_1882_18 <= _T_1745;
    end
    if (reset) begin
      _T_1882_19 <= 1'h0;
    end else if (_T_1616) begin
      _T_1882_19 <= _T_1746;
    end
    if (reset) begin
      _T_1882_20 <= 1'h0;
    end else if (_T_1616) begin
      _T_1882_20 <= _T_1747;
    end
    if (reset) begin
      _T_1663 <= 21'h1fffff;
    end else if (_T_1686) begin
      _T_1663 <= _T_1702;
    end
    if (reset) begin
      _T_401 <= 1'h0;
    end else if (_T_411) begin
      _T_401 <= 1'h0;
    end else begin
      _T_401 <= _GEN_2;
    end
    if (reset) begin
      _T_375 <= 3'h0;
    end else begin
      _T_375 <= _T_380;
    end
    if (_T_371) begin
      _T_376 <= _T_341;
    end
    _T_2060 <= reset | _GEN_93;
    if (reset) begin
      _T_2326_0 <= 1'h0;
    end else if (_T_2060) begin
      _T_2326_0 <= _T_2171;
    end
    if (reset) begin
      _T_2326_1 <= 1'h0;
    end else if (_T_2060) begin
      _T_2326_1 <= _T_2172;
    end
    if (reset) begin
      _T_2326_2 <= 1'h0;
    end else if (_T_2060) begin
      _T_2326_2 <= _T_2173;
    end
    if (reset) begin
      _T_2326_3 <= 1'h0;
    end else if (_T_2060) begin
      _T_2326_3 <= _T_2174;
    end
    if (reset) begin
      _T_2326_4 <= 1'h0;
    end else if (_T_2060) begin
      _T_2326_4 <= _T_2175;
    end
    if (reset) begin
      _T_2326_5 <= 1'h0;
    end else if (_T_2060) begin
      _T_2326_5 <= _T_2176;
    end
    if (reset) begin
      _T_2326_6 <= 1'h0;
    end else if (_T_2060) begin
      _T_2326_6 <= _T_2177;
    end
    if (reset) begin
      _T_2326_7 <= 1'h0;
    end else if (_T_2060) begin
      _T_2326_7 <= _T_2178;
    end
    if (reset) begin
      _T_2326_8 <= 1'h0;
    end else if (_T_2060) begin
      _T_2326_8 <= _T_2179;
    end
    if (reset) begin
      _T_2326_9 <= 1'h0;
    end else if (_T_2060) begin
      _T_2326_9 <= _T_2180;
    end
    if (reset) begin
      _T_2326_10 <= 1'h0;
    end else if (_T_2060) begin
      _T_2326_10 <= _T_2181;
    end
    if (reset) begin
      _T_2326_11 <= 1'h0;
    end else if (_T_2060) begin
      _T_2326_11 <= _T_2182;
    end
    if (reset) begin
      _T_2326_12 <= 1'h0;
    end else if (_T_2060) begin
      _T_2326_12 <= _T_2183;
    end
    if (reset) begin
      _T_2326_13 <= 1'h0;
    end else if (_T_2060) begin
      _T_2326_13 <= _T_2184;
    end
    if (reset) begin
      _T_2326_14 <= 1'h0;
    end else if (_T_2060) begin
      _T_2326_14 <= _T_2185;
    end
    if (reset) begin
      _T_2326_15 <= 1'h0;
    end else if (_T_2060) begin
      _T_2326_15 <= _T_2186;
    end
    if (reset) begin
      _T_2326_16 <= 1'h0;
    end else if (_T_2060) begin
      _T_2326_16 <= _T_2187;
    end
    if (reset) begin
      _T_2326_17 <= 1'h0;
    end else if (_T_2060) begin
      _T_2326_17 <= _T_2188;
    end
    if (reset) begin
      _T_2326_18 <= 1'h0;
    end else if (_T_2060) begin
      _T_2326_18 <= _T_2189;
    end
    if (reset) begin
      _T_2326_19 <= 1'h0;
    end else if (_T_2060) begin
      _T_2326_19 <= _T_2190;
    end
    if (reset) begin
      _T_2326_20 <= 1'h0;
    end else if (_T_2060) begin
      _T_2326_20 <= _T_2191;
    end
    if (reset) begin
      _T_2107 <= 21'h1fffff;
    end else if (_T_2130) begin
      _T_2107 <= _T_2146;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_358) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:107 assert (!resp_fire || count =/= UInt(0))\n"); // @[Xbar.scala 107:22]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_358) begin
          $fatal; // @[Xbar.scala 107:22]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_364) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:108 assert (!req_fire  || count =/= UInt(flight))\n"); // @[Xbar.scala 108:22]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_364) begin
          $fatal; // @[Xbar.scala 108:22]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_386) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:107 assert (!resp_fire || count =/= UInt(0))\n"); // @[Xbar.scala 107:22]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_386) begin
          $fatal; // @[Xbar.scala 107:22]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_392) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:108 assert (!req_fire  || count =/= UInt(flight))\n"); // @[Xbar.scala 108:22]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_392) begin
          $fatal; // @[Xbar.scala 108:22]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_707) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_707) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_728) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_728) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_751) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_751) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_772) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_772) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_795) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_795) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_816) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_816) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_839) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_839) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_860) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_860) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_883) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_883) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_904) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_904) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_927) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_927) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_948) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_948) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_971) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_971) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_992) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_992) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1015) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1015) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1036) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1036) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1059) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1059) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1080) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1080) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1103) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1103) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1124) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1124) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1147) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1147) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1168) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1168) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1191) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1191) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1212) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1212) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1235) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1235) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1256) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1256) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1279) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1279) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1300) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1300) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1323) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1323) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1344) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1344) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1367) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1367) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1388) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1388) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1411) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1411) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1432) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1432) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1455) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1455) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1476) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1476) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1499) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1499) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1520) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1520) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1543) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1543) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1564) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1564) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1587) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1587) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1608) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1608) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1855) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:256 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n"); // @[Xbar.scala 256:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1855) begin
          $fatal; // @[Xbar.scala 256:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1880) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1880) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2299) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:256 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n"); // @[Xbar.scala 256:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2299) begin
          $fatal; // @[Xbar.scala 256:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2324) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2324) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module Queue_141(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [31:0] io_enq_bits_data,
  input         io_enq_bits_last,
  input         io_deq_ready,
  output        io_deq_valid,
  output [31:0] io_deq_bits_data,
  output        io_deq_bits_last
);
  reg [31:0] _T_data [0:1]; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_0;
  wire [31:0] _T_data__T_18_data; // @[Decoupled.scala 218:24]
  wire  _T_data__T_18_addr; // @[Decoupled.scala 218:24]
  wire [31:0] _T_data__T_10_data; // @[Decoupled.scala 218:24]
  wire  _T_data__T_10_addr; // @[Decoupled.scala 218:24]
  wire  _T_data__T_10_mask; // @[Decoupled.scala 218:24]
  wire  _T_data__T_10_en; // @[Decoupled.scala 218:24]
  reg  _T_last [0:1]; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_1;
  wire  _T_last__T_18_data; // @[Decoupled.scala 218:24]
  wire  _T_last__T_18_addr; // @[Decoupled.scala 218:24]
  wire  _T_last__T_10_data; // @[Decoupled.scala 218:24]
  wire  _T_last__T_10_addr; // @[Decoupled.scala 218:24]
  wire  _T_last__T_10_mask; // @[Decoupled.scala 218:24]
  wire  _T_last__T_10_en; // @[Decoupled.scala 218:24]
  reg  value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_2;
  reg  value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_3;
  reg  _T_1; // @[Decoupled.scala 221:35]
  reg [31:0] _RAND_4;
  wire  _T_2 = value == value_1; // @[Decoupled.scala 223:41]
  wire  _T_3 = ~_T_1; // @[Decoupled.scala 224:36]
  wire  _T_4 = _T_2 & _T_3; // @[Decoupled.scala 224:33]
  wire  _T_5 = _T_2 & _T_1; // @[Decoupled.scala 225:32]
  wire  _T_6 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  _T_8 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire  _T_12 = value + 1'h1; // @[Counter.scala 39:22]
  wire  _T_14 = value_1 + 1'h1; // @[Counter.scala 39:22]
  wire  _T_15 = _T_6 != _T_8; // @[Decoupled.scala 236:16]
  assign _T_data__T_18_addr = value_1;
  assign _T_data__T_18_data = _T_data[_T_data__T_18_addr]; // @[Decoupled.scala 218:24]
  assign _T_data__T_10_data = io_enq_bits_data;
  assign _T_data__T_10_addr = value;
  assign _T_data__T_10_mask = 1'h1;
  assign _T_data__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_last__T_18_addr = value_1;
  assign _T_last__T_18_data = _T_last[_T_last__T_18_addr]; // @[Decoupled.scala 218:24]
  assign _T_last__T_10_data = io_enq_bits_last;
  assign _T_last__T_10_addr = value;
  assign _T_last__T_10_mask = 1'h1;
  assign _T_last__T_10_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~_T_5; // @[Decoupled.scala 241:16]
  assign io_deq_valid = ~_T_4; // @[Decoupled.scala 240:16]
  assign io_deq_bits_data = _T_data__T_18_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_last = _T_last__T_18_data; // @[Decoupled.scala 242:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_data[initvar] = _RAND_0[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_last[initvar] = _RAND_1[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  value = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  value_1 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T_data__T_10_en & _T_data__T_10_mask) begin
      _T_data[_T_data__T_10_addr] <= _T_data__T_10_data; // @[Decoupled.scala 218:24]
    end
    if(_T_last__T_10_en & _T_last__T_10_mask) begin
      _T_last[_T_last__T_10_addr] <= _T_last__T_10_data; // @[Decoupled.scala 218:24]
    end
    if (reset) begin
      value <= 1'h0;
    end else if (_T_6) begin
      value <= _T_12;
    end
    if (reset) begin
      value_1 <= 1'h0;
    end else if (_T_8) begin
      value_1 <= _T_14;
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else if (_T_15) begin
      _T_1 <= _T_6;
    end
  end
endmodule
module AXI4StreamBuffer(
  input         clock,
  input         reset,
  output        auto_in_ready,
  input         auto_in_valid,
  input  [31:0] auto_in_bits_data,
  input         auto_in_bits_last,
  input         auto_out_ready,
  output        auto_out_valid,
  output [31:0] auto_out_bits_data,
  output        auto_out_bits_last
);
  wire  Queue_clock; // @[Decoupled.scala 296:21]
  wire  Queue_reset; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [31:0] Queue_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_bits_last; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [31:0] Queue_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_bits_last; // @[Decoupled.scala 296:21]
  Queue_141 Queue ( // @[Decoupled.scala 296:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_last(Queue_io_enq_bits_last),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_last(Queue_io_deq_bits_last)
  );
  assign auto_in_ready = Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_out_valid = Queue_io_deq_valid; // @[LazyModule.scala 173:49]
  assign auto_out_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_bits_last = Queue_io_deq_bits_last; // @[LazyModule.scala 173:49]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_in_valid; // @[Decoupled.scala 297:22]
  assign Queue_io_enq_bits_data = auto_in_bits_data; // @[Decoupled.scala 298:21]
  assign Queue_io_enq_bits_last = auto_in_bits_last; // @[Decoupled.scala 298:21]
  assign Queue_io_deq_ready = auto_out_ready; // @[Decoupled.scala 320:15]
endmodule
module Queue_142(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [31:0] io_enq_bits_data,
  input         io_enq_bits_last,
  input         io_deq_ready,
  output        io_deq_valid,
  output [31:0] io_deq_bits_data,
  output        io_deq_bits_last
);
  reg [31:0] _T_data [0:1]; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_0;
  wire [31:0] _T_data__T_18_data; // @[Decoupled.scala 218:24]
  wire  _T_data__T_18_addr; // @[Decoupled.scala 218:24]
  wire [31:0] _T_data__T_10_data; // @[Decoupled.scala 218:24]
  wire  _T_data__T_10_addr; // @[Decoupled.scala 218:24]
  wire  _T_data__T_10_mask; // @[Decoupled.scala 218:24]
  wire  _T_data__T_10_en; // @[Decoupled.scala 218:24]
  reg  _T_last [0:1]; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_1;
  wire  _T_last__T_18_data; // @[Decoupled.scala 218:24]
  wire  _T_last__T_18_addr; // @[Decoupled.scala 218:24]
  wire  _T_last__T_10_data; // @[Decoupled.scala 218:24]
  wire  _T_last__T_10_addr; // @[Decoupled.scala 218:24]
  wire  _T_last__T_10_mask; // @[Decoupled.scala 218:24]
  wire  _T_last__T_10_en; // @[Decoupled.scala 218:24]
  reg  value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_2;
  reg  value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_3;
  reg  _T_1; // @[Decoupled.scala 221:35]
  reg [31:0] _RAND_4;
  wire  _T_2 = value == value_1; // @[Decoupled.scala 223:41]
  wire  _T_3 = ~_T_1; // @[Decoupled.scala 224:36]
  wire  _T_4 = _T_2 & _T_3; // @[Decoupled.scala 224:33]
  wire  _T_5 = _T_2 & _T_1; // @[Decoupled.scala 225:32]
  wire  _T_6 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  _T_8 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire  _T_12 = value + 1'h1; // @[Counter.scala 39:22]
  wire  _T_14 = value_1 + 1'h1; // @[Counter.scala 39:22]
  wire  _T_15 = _T_6 != _T_8; // @[Decoupled.scala 236:16]
  assign _T_data__T_18_addr = value_1;
  assign _T_data__T_18_data = _T_data[_T_data__T_18_addr]; // @[Decoupled.scala 218:24]
  assign _T_data__T_10_data = io_enq_bits_data;
  assign _T_data__T_10_addr = value;
  assign _T_data__T_10_mask = 1'h1;
  assign _T_data__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_last__T_18_addr = value_1;
  assign _T_last__T_18_data = _T_last[_T_last__T_18_addr]; // @[Decoupled.scala 218:24]
  assign _T_last__T_10_data = io_enq_bits_last;
  assign _T_last__T_10_addr = value;
  assign _T_last__T_10_mask = 1'h1;
  assign _T_last__T_10_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~_T_5; // @[Decoupled.scala 241:16]
  assign io_deq_valid = ~_T_4; // @[Decoupled.scala 240:16]
  assign io_deq_bits_data = _T_data__T_18_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_last = _T_last__T_18_data; // @[Decoupled.scala 242:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_data[initvar] = _RAND_0[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_last[initvar] = _RAND_1[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  value = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  value_1 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T_data__T_10_en & _T_data__T_10_mask) begin
      _T_data[_T_data__T_10_addr] <= _T_data__T_10_data; // @[Decoupled.scala 218:24]
    end
    if(_T_last__T_10_en & _T_last__T_10_mask) begin
      _T_last[_T_last__T_10_addr] <= _T_last__T_10_data; // @[Decoupled.scala 218:24]
    end
    if (reset) begin
      value <= 1'h0;
    end else if (_T_6) begin
      value <= _T_12;
    end
    if (reset) begin
      value_1 <= 1'h0;
    end else if (_T_8) begin
      value_1 <= _T_14;
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else if (_T_15) begin
      _T_1 <= _T_6;
    end
  end
endmodule
module AXI4StreamBuffer_1(
  input         clock,
  input         reset,
  output        auto_in_ready,
  input         auto_in_valid,
  input  [31:0] auto_in_bits_data,
  input         auto_in_bits_last,
  input         auto_out_ready,
  output        auto_out_valid,
  output [31:0] auto_out_bits_data,
  output        auto_out_bits_last
);
  wire  Queue_clock; // @[Decoupled.scala 296:21]
  wire  Queue_reset; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [31:0] Queue_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_bits_last; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [31:0] Queue_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_bits_last; // @[Decoupled.scala 296:21]
  Queue_142 Queue ( // @[Decoupled.scala 296:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_last(Queue_io_enq_bits_last),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_last(Queue_io_deq_bits_last)
  );
  assign auto_in_ready = Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_out_valid = Queue_io_deq_valid; // @[LazyModule.scala 173:49]
  assign auto_out_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_bits_last = Queue_io_deq_bits_last; // @[LazyModule.scala 173:49]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_in_valid; // @[Decoupled.scala 297:22]
  assign Queue_io_enq_bits_data = auto_in_bits_data; // @[Decoupled.scala 298:21]
  assign Queue_io_enq_bits_last = auto_in_bits_last; // @[Decoupled.scala 298:21]
  assign Queue_io_deq_ready = auto_out_ready; // @[Decoupled.scala 320:15]
endmodule
module Queue_143(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [31:0] io_enq_bits_data,
  input         io_enq_bits_last,
  input         io_deq_ready,
  output        io_deq_valid,
  output [31:0] io_deq_bits_data,
  output        io_deq_bits_last
);
  reg [31:0] _T_data [0:1]; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_0;
  wire [31:0] _T_data__T_18_data; // @[Decoupled.scala 218:24]
  wire  _T_data__T_18_addr; // @[Decoupled.scala 218:24]
  wire [31:0] _T_data__T_10_data; // @[Decoupled.scala 218:24]
  wire  _T_data__T_10_addr; // @[Decoupled.scala 218:24]
  wire  _T_data__T_10_mask; // @[Decoupled.scala 218:24]
  wire  _T_data__T_10_en; // @[Decoupled.scala 218:24]
  reg  _T_last [0:1]; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_1;
  wire  _T_last__T_18_data; // @[Decoupled.scala 218:24]
  wire  _T_last__T_18_addr; // @[Decoupled.scala 218:24]
  wire  _T_last__T_10_data; // @[Decoupled.scala 218:24]
  wire  _T_last__T_10_addr; // @[Decoupled.scala 218:24]
  wire  _T_last__T_10_mask; // @[Decoupled.scala 218:24]
  wire  _T_last__T_10_en; // @[Decoupled.scala 218:24]
  reg  value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_2;
  reg  value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_3;
  reg  _T_1; // @[Decoupled.scala 221:35]
  reg [31:0] _RAND_4;
  wire  _T_2 = value == value_1; // @[Decoupled.scala 223:41]
  wire  _T_3 = ~_T_1; // @[Decoupled.scala 224:36]
  wire  _T_4 = _T_2 & _T_3; // @[Decoupled.scala 224:33]
  wire  _T_5 = _T_2 & _T_1; // @[Decoupled.scala 225:32]
  wire  _T_6 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  _T_8 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire  _T_12 = value + 1'h1; // @[Counter.scala 39:22]
  wire  _T_14 = value_1 + 1'h1; // @[Counter.scala 39:22]
  wire  _T_15 = _T_6 != _T_8; // @[Decoupled.scala 236:16]
  assign _T_data__T_18_addr = value_1;
  assign _T_data__T_18_data = _T_data[_T_data__T_18_addr]; // @[Decoupled.scala 218:24]
  assign _T_data__T_10_data = io_enq_bits_data;
  assign _T_data__T_10_addr = value;
  assign _T_data__T_10_mask = 1'h1;
  assign _T_data__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_last__T_18_addr = value_1;
  assign _T_last__T_18_data = _T_last[_T_last__T_18_addr]; // @[Decoupled.scala 218:24]
  assign _T_last__T_10_data = io_enq_bits_last;
  assign _T_last__T_10_addr = value;
  assign _T_last__T_10_mask = 1'h1;
  assign _T_last__T_10_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~_T_5; // @[Decoupled.scala 241:16]
  assign io_deq_valid = ~_T_4; // @[Decoupled.scala 240:16]
  assign io_deq_bits_data = _T_data__T_18_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_last = _T_last__T_18_data; // @[Decoupled.scala 242:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_data[initvar] = _RAND_0[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_last[initvar] = _RAND_1[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  value = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  value_1 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T_data__T_10_en & _T_data__T_10_mask) begin
      _T_data[_T_data__T_10_addr] <= _T_data__T_10_data; // @[Decoupled.scala 218:24]
    end
    if(_T_last__T_10_en & _T_last__T_10_mask) begin
      _T_last[_T_last__T_10_addr] <= _T_last__T_10_data; // @[Decoupled.scala 218:24]
    end
    if (reset) begin
      value <= 1'h0;
    end else if (_T_6) begin
      value <= _T_12;
    end
    if (reset) begin
      value_1 <= 1'h0;
    end else if (_T_8) begin
      value_1 <= _T_14;
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else if (_T_15) begin
      _T_1 <= _T_6;
    end
  end
endmodule
module AXI4StreamBuffer_2(
  input         clock,
  input         reset,
  output        auto_in_ready,
  input         auto_in_valid,
  input  [31:0] auto_in_bits_data,
  input         auto_in_bits_last,
  input         auto_out_ready,
  output        auto_out_valid,
  output [31:0] auto_out_bits_data,
  output        auto_out_bits_last
);
  wire  Queue_clock; // @[Decoupled.scala 296:21]
  wire  Queue_reset; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [31:0] Queue_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_bits_last; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [31:0] Queue_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_bits_last; // @[Decoupled.scala 296:21]
  Queue_143 Queue ( // @[Decoupled.scala 296:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_last(Queue_io_enq_bits_last),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_last(Queue_io_deq_bits_last)
  );
  assign auto_in_ready = Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_out_valid = Queue_io_deq_valid; // @[LazyModule.scala 173:49]
  assign auto_out_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_bits_last = Queue_io_deq_bits_last; // @[LazyModule.scala 173:49]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_in_valid; // @[Decoupled.scala 297:22]
  assign Queue_io_enq_bits_data = auto_in_bits_data; // @[Decoupled.scala 298:21]
  assign Queue_io_enq_bits_last = auto_in_bits_last; // @[Decoupled.scala 298:21]
  assign Queue_io_deq_ready = auto_out_ready; // @[Decoupled.scala 320:15]
endmodule
module Queue_145(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [31:0] io_enq_bits_data,
  input         io_enq_bits_last,
  input         io_deq_ready,
  output        io_deq_valid,
  output [31:0] io_deq_bits_data,
  output        io_deq_bits_last
);
  reg [31:0] _T_data [0:1]; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_0;
  wire [31:0] _T_data__T_18_data; // @[Decoupled.scala 218:24]
  wire  _T_data__T_18_addr; // @[Decoupled.scala 218:24]
  wire [31:0] _T_data__T_10_data; // @[Decoupled.scala 218:24]
  wire  _T_data__T_10_addr; // @[Decoupled.scala 218:24]
  wire  _T_data__T_10_mask; // @[Decoupled.scala 218:24]
  wire  _T_data__T_10_en; // @[Decoupled.scala 218:24]
  reg  _T_last [0:1]; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_1;
  wire  _T_last__T_18_data; // @[Decoupled.scala 218:24]
  wire  _T_last__T_18_addr; // @[Decoupled.scala 218:24]
  wire  _T_last__T_10_data; // @[Decoupled.scala 218:24]
  wire  _T_last__T_10_addr; // @[Decoupled.scala 218:24]
  wire  _T_last__T_10_mask; // @[Decoupled.scala 218:24]
  wire  _T_last__T_10_en; // @[Decoupled.scala 218:24]
  reg  value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_2;
  reg  value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_3;
  reg  _T_1; // @[Decoupled.scala 221:35]
  reg [31:0] _RAND_4;
  wire  _T_2 = value == value_1; // @[Decoupled.scala 223:41]
  wire  _T_3 = ~_T_1; // @[Decoupled.scala 224:36]
  wire  _T_4 = _T_2 & _T_3; // @[Decoupled.scala 224:33]
  wire  _T_5 = _T_2 & _T_1; // @[Decoupled.scala 225:32]
  wire  _T_6 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  _T_8 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire  _T_12 = value + 1'h1; // @[Counter.scala 39:22]
  wire  _T_14 = value_1 + 1'h1; // @[Counter.scala 39:22]
  wire  _T_15 = _T_6 != _T_8; // @[Decoupled.scala 236:16]
  assign _T_data__T_18_addr = value_1;
  assign _T_data__T_18_data = _T_data[_T_data__T_18_addr]; // @[Decoupled.scala 218:24]
  assign _T_data__T_10_data = io_enq_bits_data;
  assign _T_data__T_10_addr = value;
  assign _T_data__T_10_mask = 1'h1;
  assign _T_data__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_last__T_18_addr = value_1;
  assign _T_last__T_18_data = _T_last[_T_last__T_18_addr]; // @[Decoupled.scala 218:24]
  assign _T_last__T_10_data = io_enq_bits_last;
  assign _T_last__T_10_addr = value;
  assign _T_last__T_10_mask = 1'h1;
  assign _T_last__T_10_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~_T_5; // @[Decoupled.scala 241:16]
  assign io_deq_valid = ~_T_4; // @[Decoupled.scala 240:16]
  assign io_deq_bits_data = _T_data__T_18_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_last = _T_last__T_18_data; // @[Decoupled.scala 242:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_data[initvar] = _RAND_0[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_last[initvar] = _RAND_1[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  value = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  value_1 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T_data__T_10_en & _T_data__T_10_mask) begin
      _T_data[_T_data__T_10_addr] <= _T_data__T_10_data; // @[Decoupled.scala 218:24]
    end
    if(_T_last__T_10_en & _T_last__T_10_mask) begin
      _T_last[_T_last__T_10_addr] <= _T_last__T_10_data; // @[Decoupled.scala 218:24]
    end
    if (reset) begin
      value <= 1'h0;
    end else if (_T_6) begin
      value <= _T_12;
    end
    if (reset) begin
      value_1 <= 1'h0;
    end else if (_T_8) begin
      value_1 <= _T_14;
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else if (_T_15) begin
      _T_1 <= _T_6;
    end
  end
endmodule
module AXI4StreamBuffer_4(
  input         clock,
  input         reset,
  output        auto_in_ready,
  input         auto_in_valid,
  input  [31:0] auto_in_bits_data,
  input         auto_in_bits_last,
  input         auto_out_ready,
  output        auto_out_valid,
  output [31:0] auto_out_bits_data,
  output        auto_out_bits_last
);
  wire  Queue_clock; // @[Decoupled.scala 296:21]
  wire  Queue_reset; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [31:0] Queue_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_bits_last; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [31:0] Queue_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_bits_last; // @[Decoupled.scala 296:21]
  Queue_145 Queue ( // @[Decoupled.scala 296:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_last(Queue_io_enq_bits_last),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_last(Queue_io_deq_bits_last)
  );
  assign auto_in_ready = Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_out_valid = Queue_io_deq_valid; // @[LazyModule.scala 173:49]
  assign auto_out_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_bits_last = Queue_io_deq_bits_last; // @[LazyModule.scala 173:49]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_in_valid; // @[Decoupled.scala 297:22]
  assign Queue_io_enq_bits_data = auto_in_bits_data; // @[Decoupled.scala 298:21]
  assign Queue_io_enq_bits_last = auto_in_bits_last; // @[Decoupled.scala 298:21]
  assign Queue_io_deq_ready = auto_out_ready; // @[Decoupled.scala 320:15]
endmodule
module Queue_146(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [31:0] io_enq_bits_data,
  input         io_enq_bits_last,
  input         io_deq_ready,
  output        io_deq_valid,
  output [31:0] io_deq_bits_data,
  output        io_deq_bits_last
);
  reg [31:0] _T_data [0:1]; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_0;
  wire [31:0] _T_data__T_18_data; // @[Decoupled.scala 218:24]
  wire  _T_data__T_18_addr; // @[Decoupled.scala 218:24]
  wire [31:0] _T_data__T_10_data; // @[Decoupled.scala 218:24]
  wire  _T_data__T_10_addr; // @[Decoupled.scala 218:24]
  wire  _T_data__T_10_mask; // @[Decoupled.scala 218:24]
  wire  _T_data__T_10_en; // @[Decoupled.scala 218:24]
  reg  _T_last [0:1]; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_1;
  wire  _T_last__T_18_data; // @[Decoupled.scala 218:24]
  wire  _T_last__T_18_addr; // @[Decoupled.scala 218:24]
  wire  _T_last__T_10_data; // @[Decoupled.scala 218:24]
  wire  _T_last__T_10_addr; // @[Decoupled.scala 218:24]
  wire  _T_last__T_10_mask; // @[Decoupled.scala 218:24]
  wire  _T_last__T_10_en; // @[Decoupled.scala 218:24]
  reg  value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_2;
  reg  value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_3;
  reg  _T_1; // @[Decoupled.scala 221:35]
  reg [31:0] _RAND_4;
  wire  _T_2 = value == value_1; // @[Decoupled.scala 223:41]
  wire  _T_3 = ~_T_1; // @[Decoupled.scala 224:36]
  wire  _T_4 = _T_2 & _T_3; // @[Decoupled.scala 224:33]
  wire  _T_5 = _T_2 & _T_1; // @[Decoupled.scala 225:32]
  wire  _T_6 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  _T_8 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire  _T_12 = value + 1'h1; // @[Counter.scala 39:22]
  wire  _T_14 = value_1 + 1'h1; // @[Counter.scala 39:22]
  wire  _T_15 = _T_6 != _T_8; // @[Decoupled.scala 236:16]
  assign _T_data__T_18_addr = value_1;
  assign _T_data__T_18_data = _T_data[_T_data__T_18_addr]; // @[Decoupled.scala 218:24]
  assign _T_data__T_10_data = io_enq_bits_data;
  assign _T_data__T_10_addr = value;
  assign _T_data__T_10_mask = 1'h1;
  assign _T_data__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_last__T_18_addr = value_1;
  assign _T_last__T_18_data = _T_last[_T_last__T_18_addr]; // @[Decoupled.scala 218:24]
  assign _T_last__T_10_data = io_enq_bits_last;
  assign _T_last__T_10_addr = value;
  assign _T_last__T_10_mask = 1'h1;
  assign _T_last__T_10_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~_T_5; // @[Decoupled.scala 241:16]
  assign io_deq_valid = ~_T_4; // @[Decoupled.scala 240:16]
  assign io_deq_bits_data = _T_data__T_18_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_last = _T_last__T_18_data; // @[Decoupled.scala 242:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_data[initvar] = _RAND_0[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_last[initvar] = _RAND_1[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  value = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  value_1 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T_data__T_10_en & _T_data__T_10_mask) begin
      _T_data[_T_data__T_10_addr] <= _T_data__T_10_data; // @[Decoupled.scala 218:24]
    end
    if(_T_last__T_10_en & _T_last__T_10_mask) begin
      _T_last[_T_last__T_10_addr] <= _T_last__T_10_data; // @[Decoupled.scala 218:24]
    end
    if (reset) begin
      value <= 1'h0;
    end else if (_T_6) begin
      value <= _T_12;
    end
    if (reset) begin
      value_1 <= 1'h0;
    end else if (_T_8) begin
      value_1 <= _T_14;
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else if (_T_15) begin
      _T_1 <= _T_6;
    end
  end
endmodule
module AXI4StreamBuffer_5(
  input         clock,
  input         reset,
  output        auto_in_ready,
  input         auto_in_valid,
  input  [31:0] auto_in_bits_data,
  input         auto_in_bits_last,
  input         auto_out_ready,
  output        auto_out_valid,
  output [31:0] auto_out_bits_data,
  output        auto_out_bits_last
);
  wire  Queue_clock; // @[Decoupled.scala 296:21]
  wire  Queue_reset; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [31:0] Queue_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_bits_last; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [31:0] Queue_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_bits_last; // @[Decoupled.scala 296:21]
  Queue_146 Queue ( // @[Decoupled.scala 296:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_last(Queue_io_enq_bits_last),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_last(Queue_io_deq_bits_last)
  );
  assign auto_in_ready = Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_out_valid = Queue_io_deq_valid; // @[LazyModule.scala 173:49]
  assign auto_out_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_bits_last = Queue_io_deq_bits_last; // @[LazyModule.scala 173:49]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_in_valid; // @[Decoupled.scala 297:22]
  assign Queue_io_enq_bits_data = auto_in_bits_data; // @[Decoupled.scala 298:21]
  assign Queue_io_enq_bits_last = auto_in_bits_last; // @[Decoupled.scala 298:21]
  assign Queue_io_deq_ready = auto_out_ready; // @[Decoupled.scala 320:15]
endmodule
module Queue_150(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [31:0] io_enq_bits_data,
  input         io_enq_bits_last,
  input         io_deq_ready,
  output        io_deq_valid,
  output [31:0] io_deq_bits_data,
  output        io_deq_bits_last
);
  reg [31:0] _T_data [0:1]; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_0;
  wire [31:0] _T_data__T_18_data; // @[Decoupled.scala 218:24]
  wire  _T_data__T_18_addr; // @[Decoupled.scala 218:24]
  wire [31:0] _T_data__T_10_data; // @[Decoupled.scala 218:24]
  wire  _T_data__T_10_addr; // @[Decoupled.scala 218:24]
  wire  _T_data__T_10_mask; // @[Decoupled.scala 218:24]
  wire  _T_data__T_10_en; // @[Decoupled.scala 218:24]
  reg  _T_last [0:1]; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_1;
  wire  _T_last__T_18_data; // @[Decoupled.scala 218:24]
  wire  _T_last__T_18_addr; // @[Decoupled.scala 218:24]
  wire  _T_last__T_10_data; // @[Decoupled.scala 218:24]
  wire  _T_last__T_10_addr; // @[Decoupled.scala 218:24]
  wire  _T_last__T_10_mask; // @[Decoupled.scala 218:24]
  wire  _T_last__T_10_en; // @[Decoupled.scala 218:24]
  reg  value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_2;
  reg  value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_3;
  reg  _T_1; // @[Decoupled.scala 221:35]
  reg [31:0] _RAND_4;
  wire  _T_2 = value == value_1; // @[Decoupled.scala 223:41]
  wire  _T_3 = ~_T_1; // @[Decoupled.scala 224:36]
  wire  _T_4 = _T_2 & _T_3; // @[Decoupled.scala 224:33]
  wire  _T_5 = _T_2 & _T_1; // @[Decoupled.scala 225:32]
  wire  _T_6 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  _T_8 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire  _T_12 = value + 1'h1; // @[Counter.scala 39:22]
  wire  _T_14 = value_1 + 1'h1; // @[Counter.scala 39:22]
  wire  _T_15 = _T_6 != _T_8; // @[Decoupled.scala 236:16]
  assign _T_data__T_18_addr = value_1;
  assign _T_data__T_18_data = _T_data[_T_data__T_18_addr]; // @[Decoupled.scala 218:24]
  assign _T_data__T_10_data = io_enq_bits_data;
  assign _T_data__T_10_addr = value;
  assign _T_data__T_10_mask = 1'h1;
  assign _T_data__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_last__T_18_addr = value_1;
  assign _T_last__T_18_data = _T_last[_T_last__T_18_addr]; // @[Decoupled.scala 218:24]
  assign _T_last__T_10_data = io_enq_bits_last;
  assign _T_last__T_10_addr = value;
  assign _T_last__T_10_mask = 1'h1;
  assign _T_last__T_10_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~_T_5; // @[Decoupled.scala 241:16]
  assign io_deq_valid = ~_T_4; // @[Decoupled.scala 240:16]
  assign io_deq_bits_data = _T_data__T_18_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_last = _T_last__T_18_data; // @[Decoupled.scala 242:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_data[initvar] = _RAND_0[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_last[initvar] = _RAND_1[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  value = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  value_1 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T_data__T_10_en & _T_data__T_10_mask) begin
      _T_data[_T_data__T_10_addr] <= _T_data__T_10_data; // @[Decoupled.scala 218:24]
    end
    if(_T_last__T_10_en & _T_last__T_10_mask) begin
      _T_last[_T_last__T_10_addr] <= _T_last__T_10_data; // @[Decoupled.scala 218:24]
    end
    if (reset) begin
      value <= 1'h0;
    end else if (_T_6) begin
      value <= _T_12;
    end
    if (reset) begin
      value_1 <= 1'h0;
    end else if (_T_8) begin
      value_1 <= _T_14;
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else if (_T_15) begin
      _T_1 <= _T_6;
    end
  end
endmodule
module AXI4StreamBuffer_9(
  input         clock,
  input         reset,
  output        auto_in_ready,
  input         auto_in_valid,
  input  [31:0] auto_in_bits_data,
  input         auto_in_bits_last,
  input         auto_out_ready,
  output        auto_out_valid,
  output [31:0] auto_out_bits_data,
  output        auto_out_bits_last
);
  wire  Queue_clock; // @[Decoupled.scala 296:21]
  wire  Queue_reset; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [31:0] Queue_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire  Queue_io_enq_bits_last; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [31:0] Queue_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire  Queue_io_deq_bits_last; // @[Decoupled.scala 296:21]
  Queue_150 Queue ( // @[Decoupled.scala 296:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_last(Queue_io_enq_bits_last),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_last(Queue_io_deq_bits_last)
  );
  assign auto_in_ready = Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_out_valid = Queue_io_deq_valid; // @[LazyModule.scala 173:49]
  assign auto_out_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_bits_last = Queue_io_deq_bits_last; // @[LazyModule.scala 173:49]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_in_valid; // @[Decoupled.scala 297:22]
  assign Queue_io_enq_bits_data = auto_in_bits_data; // @[Decoupled.scala 298:21]
  assign Queue_io_enq_bits_last = auto_in_bits_last; // @[Decoupled.scala 298:21]
  assign Queue_io_deq_ready = auto_out_ready; // @[Decoupled.scala 320:15]
endmodule
module BundleBridgeToAXI4(
  output        auto_in_aw_ready,
  input         auto_in_aw_valid,
  input         auto_in_aw_bits_id,
  input  [31:0] auto_in_aw_bits_addr,
  input  [2:0]  auto_in_aw_bits_size,
  output        auto_in_w_ready,
  input         auto_in_w_valid,
  input  [31:0] auto_in_w_bits_data,
  input  [3:0]  auto_in_w_bits_strb,
  input         auto_in_w_bits_last,
  input         auto_in_b_ready,
  output        auto_in_b_valid,
  output [1:0]  auto_in_b_bits_resp,
  output        auto_in_ar_ready,
  input         auto_in_ar_valid,
  input         auto_in_ar_bits_id,
  input  [31:0] auto_in_ar_bits_addr,
  input  [2:0]  auto_in_ar_bits_size,
  input         auto_in_r_ready,
  output        auto_in_r_valid,
  output [31:0] auto_in_r_bits_data,
  output [1:0]  auto_in_r_bits_resp,
  output        auto_in_r_bits_last,
  input         auto_out_aw_ready,
  output        auto_out_aw_valid,
  output        auto_out_aw_bits_id,
  output [29:0] auto_out_aw_bits_addr,
  output [2:0]  auto_out_aw_bits_size,
  input         auto_out_w_ready,
  output        auto_out_w_valid,
  output [31:0] auto_out_w_bits_data,
  output [3:0]  auto_out_w_bits_strb,
  output        auto_out_w_bits_last,
  output        auto_out_b_ready,
  input         auto_out_b_valid,
  input  [1:0]  auto_out_b_bits_resp,
  input         auto_out_ar_ready,
  output        auto_out_ar_valid,
  output        auto_out_ar_bits_id,
  output [29:0] auto_out_ar_bits_addr,
  output [2:0]  auto_out_ar_bits_size,
  output        auto_out_r_ready,
  input         auto_out_r_valid,
  input  [31:0] auto_out_r_bits_data,
  input  [1:0]  auto_out_r_bits_resp,
  input         auto_out_r_bits_last
);
  assign auto_in_aw_ready = auto_out_aw_ready; // @[LazyModule.scala 173:31]
  assign auto_in_w_ready = auto_out_w_ready; // @[LazyModule.scala 173:31]
  assign auto_in_b_valid = auto_out_b_valid; // @[LazyModule.scala 173:31]
  assign auto_in_b_bits_resp = auto_out_b_bits_resp; // @[LazyModule.scala 173:31]
  assign auto_in_ar_ready = auto_out_ar_ready; // @[LazyModule.scala 173:31]
  assign auto_in_r_valid = auto_out_r_valid; // @[LazyModule.scala 173:31]
  assign auto_in_r_bits_data = auto_out_r_bits_data; // @[LazyModule.scala 173:31]
  assign auto_in_r_bits_resp = auto_out_r_bits_resp; // @[LazyModule.scala 173:31]
  assign auto_in_r_bits_last = auto_out_r_bits_last; // @[LazyModule.scala 173:31]
  assign auto_out_aw_valid = auto_in_aw_valid; // @[LazyModule.scala 173:49]
  assign auto_out_aw_bits_id = auto_in_aw_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_aw_bits_addr = auto_in_aw_bits_addr[29:0]; // @[LazyModule.scala 173:49]
  assign auto_out_aw_bits_size = auto_in_aw_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_w_valid = auto_in_w_valid; // @[LazyModule.scala 173:49]
  assign auto_out_w_bits_data = auto_in_w_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_w_bits_strb = auto_in_w_bits_strb; // @[LazyModule.scala 173:49]
  assign auto_out_w_bits_last = auto_in_w_bits_last; // @[LazyModule.scala 173:49]
  assign auto_out_b_ready = auto_in_b_ready; // @[LazyModule.scala 173:49]
  assign auto_out_ar_valid = auto_in_ar_valid; // @[LazyModule.scala 173:49]
  assign auto_out_ar_bits_id = auto_in_ar_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_ar_bits_addr = auto_in_ar_bits_addr[29:0]; // @[LazyModule.scala 173:49]
  assign auto_out_ar_bits_size = auto_in_ar_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_r_ready = auto_in_r_ready; // @[LazyModule.scala 173:49]
endmodule
module AXI4StreamToBundleBridge(
  output       auto_in_ready,
  input        auto_in_valid,
  input  [7:0] auto_in_bits_data,
  input        auto_in_bits_last,
  input        auto_out_ready,
  output       auto_out_valid,
  output [7:0] auto_out_bits_data,
  output       auto_out_bits_last
);
  assign auto_in_ready = auto_out_ready; // @[LazyModule.scala 173:31]
  assign auto_out_valid = auto_in_valid; // @[LazyModule.scala 173:49]
  assign auto_out_bits_data = auto_in_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_bits_last = auto_in_bits_last; // @[LazyModule.scala 173:49]
endmodule
module SpectrometerTest(
  input         clock,
  input         reset,
  output        ioMem_0_aw_ready,
  input         ioMem_0_aw_valid,
  input         ioMem_0_aw_bits_id,
  input  [31:0] ioMem_0_aw_bits_addr,
  input  [7:0]  ioMem_0_aw_bits_len,
  input  [2:0]  ioMem_0_aw_bits_size,
  input  [1:0]  ioMem_0_aw_bits_burst,
  input         ioMem_0_aw_bits_lock,
  input  [3:0]  ioMem_0_aw_bits_cache,
  input  [2:0]  ioMem_0_aw_bits_prot,
  input  [3:0]  ioMem_0_aw_bits_qos,
  output        ioMem_0_w_ready,
  input         ioMem_0_w_valid,
  input  [31:0] ioMem_0_w_bits_data,
  input  [3:0]  ioMem_0_w_bits_strb,
  input         ioMem_0_w_bits_last,
  input         ioMem_0_b_ready,
  output        ioMem_0_b_valid,
  output        ioMem_0_b_bits_id,
  output [1:0]  ioMem_0_b_bits_resp,
  output        ioMem_0_ar_ready,
  input         ioMem_0_ar_valid,
  input         ioMem_0_ar_bits_id,
  input  [31:0] ioMem_0_ar_bits_addr,
  input  [7:0]  ioMem_0_ar_bits_len,
  input  [2:0]  ioMem_0_ar_bits_size,
  input  [1:0]  ioMem_0_ar_bits_burst,
  input         ioMem_0_ar_bits_lock,
  input  [3:0]  ioMem_0_ar_bits_cache,
  input  [2:0]  ioMem_0_ar_bits_prot,
  input  [3:0]  ioMem_0_ar_bits_qos,
  input         ioMem_0_r_ready,
  output        ioMem_0_r_valid,
  output        ioMem_0_r_bits_id,
  output [31:0] ioMem_0_r_bits_data,
  output [1:0]  ioMem_0_r_bits_resp,
  output        ioMem_0_r_bits_last,
  input         outStream_0_ready,
  output        outStream_0_valid,
  output [7:0]  outStream_0_bits_data,
  output        outStream_0_bits_last,
  output        inStream_0_ready,
  input         inStream_0_valid,
  input  [7:0]  inStream_0_bits_data,
  input         inStream_0_bits_last,
  output        int_0,
  output        uTx,
  input         uRx
);
  wire  widthAdapter_clock; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_reset; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_auto_in_ready; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_auto_in_valid; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire [7:0] widthAdapter_auto_in_bits_data; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_auto_in_bits_last; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_auto_out_ready; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_auto_out_valid; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire [31:0] widthAdapter_auto_out_bits_data; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_auto_out_bits_last; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  in_split_clock; // @[SpectrometerTest.scala 114:29]
  wire  in_split_reset; // @[SpectrometerTest.scala 114:29]
  wire  in_split_auto_mem_in_aw_ready; // @[SpectrometerTest.scala 114:29]
  wire  in_split_auto_mem_in_aw_valid; // @[SpectrometerTest.scala 114:29]
  wire  in_split_auto_mem_in_aw_bits_id; // @[SpectrometerTest.scala 114:29]
  wire [29:0] in_split_auto_mem_in_aw_bits_addr; // @[SpectrometerTest.scala 114:29]
  wire  in_split_auto_mem_in_w_ready; // @[SpectrometerTest.scala 114:29]
  wire  in_split_auto_mem_in_w_valid; // @[SpectrometerTest.scala 114:29]
  wire [31:0] in_split_auto_mem_in_w_bits_data; // @[SpectrometerTest.scala 114:29]
  wire [3:0] in_split_auto_mem_in_w_bits_strb; // @[SpectrometerTest.scala 114:29]
  wire  in_split_auto_mem_in_b_ready; // @[SpectrometerTest.scala 114:29]
  wire  in_split_auto_mem_in_b_valid; // @[SpectrometerTest.scala 114:29]
  wire  in_split_auto_mem_in_b_bits_id; // @[SpectrometerTest.scala 114:29]
  wire  in_split_auto_mem_in_ar_ready; // @[SpectrometerTest.scala 114:29]
  wire  in_split_auto_mem_in_ar_valid; // @[SpectrometerTest.scala 114:29]
  wire  in_split_auto_mem_in_ar_bits_id; // @[SpectrometerTest.scala 114:29]
  wire [29:0] in_split_auto_mem_in_ar_bits_addr; // @[SpectrometerTest.scala 114:29]
  wire [2:0] in_split_auto_mem_in_ar_bits_size; // @[SpectrometerTest.scala 114:29]
  wire  in_split_auto_mem_in_r_ready; // @[SpectrometerTest.scala 114:29]
  wire  in_split_auto_mem_in_r_valid; // @[SpectrometerTest.scala 114:29]
  wire  in_split_auto_mem_in_r_bits_id; // @[SpectrometerTest.scala 114:29]
  wire [31:0] in_split_auto_mem_in_r_bits_data; // @[SpectrometerTest.scala 114:29]
  wire  in_split_auto_stream_in_ready; // @[SpectrometerTest.scala 114:29]
  wire  in_split_auto_stream_in_valid; // @[SpectrometerTest.scala 114:29]
  wire [31:0] in_split_auto_stream_in_bits_data; // @[SpectrometerTest.scala 114:29]
  wire  in_split_auto_stream_in_bits_last; // @[SpectrometerTest.scala 114:29]
  wire  in_split_auto_stream_out_4_ready; // @[SpectrometerTest.scala 114:29]
  wire  in_split_auto_stream_out_4_valid; // @[SpectrometerTest.scala 114:29]
  wire [31:0] in_split_auto_stream_out_4_bits_data; // @[SpectrometerTest.scala 114:29]
  wire  in_split_auto_stream_out_4_bits_last; // @[SpectrometerTest.scala 114:29]
  wire  in_split_auto_stream_out_3_ready; // @[SpectrometerTest.scala 114:29]
  wire  in_split_auto_stream_out_3_valid; // @[SpectrometerTest.scala 114:29]
  wire [31:0] in_split_auto_stream_out_3_bits_data; // @[SpectrometerTest.scala 114:29]
  wire  in_split_auto_stream_out_3_bits_last; // @[SpectrometerTest.scala 114:29]
  wire  in_split_auto_stream_out_2_ready; // @[SpectrometerTest.scala 114:29]
  wire  in_split_auto_stream_out_2_valid; // @[SpectrometerTest.scala 114:29]
  wire [31:0] in_split_auto_stream_out_2_bits_data; // @[SpectrometerTest.scala 114:29]
  wire  in_split_auto_stream_out_2_bits_last; // @[SpectrometerTest.scala 114:29]
  wire  in_split_auto_stream_out_1_ready; // @[SpectrometerTest.scala 114:29]
  wire  in_split_auto_stream_out_1_valid; // @[SpectrometerTest.scala 114:29]
  wire [31:0] in_split_auto_stream_out_1_bits_data; // @[SpectrometerTest.scala 114:29]
  wire  in_split_auto_stream_out_1_bits_last; // @[SpectrometerTest.scala 114:29]
  wire  in_split_auto_stream_out_0_ready; // @[SpectrometerTest.scala 114:29]
  wire  in_split_auto_stream_out_0_valid; // @[SpectrometerTest.scala 114:29]
  wire [31:0] in_split_auto_stream_out_0_bits_data; // @[SpectrometerTest.scala 114:29]
  wire  in_split_auto_stream_out_0_bits_last; // @[SpectrometerTest.scala 114:29]
  wire  in_queue_clock; // @[SpectrometerTest.scala 115:29]
  wire  in_queue_reset; // @[SpectrometerTest.scala 115:29]
  wire  in_queue_auto_out_out_ready; // @[SpectrometerTest.scala 115:29]
  wire  in_queue_auto_out_out_valid; // @[SpectrometerTest.scala 115:29]
  wire [7:0] in_queue_auto_out_out_bits_data; // @[SpectrometerTest.scala 115:29]
  wire  in_queue_auto_out_out_bits_last; // @[SpectrometerTest.scala 115:29]
  wire  in_queue_auto_in_in_ready; // @[SpectrometerTest.scala 115:29]
  wire  in_queue_auto_in_in_valid; // @[SpectrometerTest.scala 115:29]
  wire [7:0] in_queue_auto_in_in_bits_data; // @[SpectrometerTest.scala 115:29]
  wire  in_queue_auto_in_in_bits_last; // @[SpectrometerTest.scala 115:29]
  wire  plfg_clock; // @[SpectrometerTest.scala 117:30]
  wire  plfg_reset; // @[SpectrometerTest.scala 117:30]
  wire  plfg_auto_mem_in_aw_ready; // @[SpectrometerTest.scala 117:30]
  wire  plfg_auto_mem_in_aw_valid; // @[SpectrometerTest.scala 117:30]
  wire  plfg_auto_mem_in_aw_bits_id; // @[SpectrometerTest.scala 117:30]
  wire [29:0] plfg_auto_mem_in_aw_bits_addr; // @[SpectrometerTest.scala 117:30]
  wire  plfg_auto_mem_in_w_ready; // @[SpectrometerTest.scala 117:30]
  wire  plfg_auto_mem_in_w_valid; // @[SpectrometerTest.scala 117:30]
  wire [31:0] plfg_auto_mem_in_w_bits_data; // @[SpectrometerTest.scala 117:30]
  wire [3:0] plfg_auto_mem_in_w_bits_strb; // @[SpectrometerTest.scala 117:30]
  wire  plfg_auto_mem_in_w_bits_last; // @[SpectrometerTest.scala 117:30]
  wire  plfg_auto_mem_in_b_ready; // @[SpectrometerTest.scala 117:30]
  wire  plfg_auto_mem_in_b_valid; // @[SpectrometerTest.scala 117:30]
  wire [1:0] plfg_auto_mem_in_b_bits_resp; // @[SpectrometerTest.scala 117:30]
  wire  plfg_auto_mem_in_ar_ready; // @[SpectrometerTest.scala 117:30]
  wire  plfg_auto_mem_in_ar_valid; // @[SpectrometerTest.scala 117:30]
  wire  plfg_auto_mem_in_ar_bits_id; // @[SpectrometerTest.scala 117:30]
  wire [29:0] plfg_auto_mem_in_ar_bits_addr; // @[SpectrometerTest.scala 117:30]
  wire [2:0] plfg_auto_mem_in_ar_bits_size; // @[SpectrometerTest.scala 117:30]
  wire  plfg_auto_mem_in_r_ready; // @[SpectrometerTest.scala 117:30]
  wire  plfg_auto_mem_in_r_valid; // @[SpectrometerTest.scala 117:30]
  wire [31:0] plfg_auto_mem_in_r_bits_data; // @[SpectrometerTest.scala 117:30]
  wire [1:0] plfg_auto_mem_in_r_bits_resp; // @[SpectrometerTest.scala 117:30]
  wire  plfg_auto_mem_in_r_bits_last; // @[SpectrometerTest.scala 117:30]
  wire  plfg_auto_stream_out_ready; // @[SpectrometerTest.scala 117:30]
  wire  plfg_auto_stream_out_valid; // @[SpectrometerTest.scala 117:30]
  wire [31:0] plfg_auto_stream_out_bits_data; // @[SpectrometerTest.scala 117:30]
  wire  plfg_auto_stream_out_bits_last; // @[SpectrometerTest.scala 117:30]
  wire  plfg_split_clock; // @[SpectrometerTest.scala 118:30]
  wire  plfg_split_reset; // @[SpectrometerTest.scala 118:30]
  wire  plfg_split_auto_mem_in_aw_ready; // @[SpectrometerTest.scala 118:30]
  wire  plfg_split_auto_mem_in_aw_valid; // @[SpectrometerTest.scala 118:30]
  wire  plfg_split_auto_mem_in_aw_bits_id; // @[SpectrometerTest.scala 118:30]
  wire [29:0] plfg_split_auto_mem_in_aw_bits_addr; // @[SpectrometerTest.scala 118:30]
  wire  plfg_split_auto_mem_in_w_ready; // @[SpectrometerTest.scala 118:30]
  wire  plfg_split_auto_mem_in_w_valid; // @[SpectrometerTest.scala 118:30]
  wire [31:0] plfg_split_auto_mem_in_w_bits_data; // @[SpectrometerTest.scala 118:30]
  wire [3:0] plfg_split_auto_mem_in_w_bits_strb; // @[SpectrometerTest.scala 118:30]
  wire  plfg_split_auto_mem_in_b_ready; // @[SpectrometerTest.scala 118:30]
  wire  plfg_split_auto_mem_in_b_valid; // @[SpectrometerTest.scala 118:30]
  wire  plfg_split_auto_mem_in_b_bits_id; // @[SpectrometerTest.scala 118:30]
  wire  plfg_split_auto_mem_in_ar_ready; // @[SpectrometerTest.scala 118:30]
  wire  plfg_split_auto_mem_in_ar_valid; // @[SpectrometerTest.scala 118:30]
  wire  plfg_split_auto_mem_in_ar_bits_id; // @[SpectrometerTest.scala 118:30]
  wire [29:0] plfg_split_auto_mem_in_ar_bits_addr; // @[SpectrometerTest.scala 118:30]
  wire [2:0] plfg_split_auto_mem_in_ar_bits_size; // @[SpectrometerTest.scala 118:30]
  wire  plfg_split_auto_mem_in_r_ready; // @[SpectrometerTest.scala 118:30]
  wire  plfg_split_auto_mem_in_r_valid; // @[SpectrometerTest.scala 118:30]
  wire  plfg_split_auto_mem_in_r_bits_id; // @[SpectrometerTest.scala 118:30]
  wire [31:0] plfg_split_auto_mem_in_r_bits_data; // @[SpectrometerTest.scala 118:30]
  wire  plfg_split_auto_stream_in_ready; // @[SpectrometerTest.scala 118:30]
  wire  plfg_split_auto_stream_in_valid; // @[SpectrometerTest.scala 118:30]
  wire [31:0] plfg_split_auto_stream_in_bits_data; // @[SpectrometerTest.scala 118:30]
  wire  plfg_split_auto_stream_in_bits_last; // @[SpectrometerTest.scala 118:30]
  wire  plfg_split_auto_stream_out_1_ready; // @[SpectrometerTest.scala 118:30]
  wire  plfg_split_auto_stream_out_1_valid; // @[SpectrometerTest.scala 118:30]
  wire [31:0] plfg_split_auto_stream_out_1_bits_data; // @[SpectrometerTest.scala 118:30]
  wire  plfg_split_auto_stream_out_1_bits_last; // @[SpectrometerTest.scala 118:30]
  wire  plfg_split_auto_stream_out_0_ready; // @[SpectrometerTest.scala 118:30]
  wire  plfg_split_auto_stream_out_0_valid; // @[SpectrometerTest.scala 118:30]
  wire [31:0] plfg_split_auto_stream_out_0_bits_data; // @[SpectrometerTest.scala 118:30]
  wire  plfg_split_auto_stream_out_0_bits_last; // @[SpectrometerTest.scala 118:30]
  wire  plfg_mux_0_clock; // @[SpectrometerTest.scala 119:30]
  wire  plfg_mux_0_reset; // @[SpectrometerTest.scala 119:30]
  wire  plfg_mux_0_auto_register_in_aw_ready; // @[SpectrometerTest.scala 119:30]
  wire  plfg_mux_0_auto_register_in_aw_valid; // @[SpectrometerTest.scala 119:30]
  wire  plfg_mux_0_auto_register_in_aw_bits_id; // @[SpectrometerTest.scala 119:30]
  wire [29:0] plfg_mux_0_auto_register_in_aw_bits_addr; // @[SpectrometerTest.scala 119:30]
  wire  plfg_mux_0_auto_register_in_w_ready; // @[SpectrometerTest.scala 119:30]
  wire  plfg_mux_0_auto_register_in_w_valid; // @[SpectrometerTest.scala 119:30]
  wire [31:0] plfg_mux_0_auto_register_in_w_bits_data; // @[SpectrometerTest.scala 119:30]
  wire [3:0] plfg_mux_0_auto_register_in_w_bits_strb; // @[SpectrometerTest.scala 119:30]
  wire  plfg_mux_0_auto_register_in_b_ready; // @[SpectrometerTest.scala 119:30]
  wire  plfg_mux_0_auto_register_in_b_valid; // @[SpectrometerTest.scala 119:30]
  wire  plfg_mux_0_auto_register_in_b_bits_id; // @[SpectrometerTest.scala 119:30]
  wire  plfg_mux_0_auto_register_in_ar_ready; // @[SpectrometerTest.scala 119:30]
  wire  plfg_mux_0_auto_register_in_ar_valid; // @[SpectrometerTest.scala 119:30]
  wire  plfg_mux_0_auto_register_in_ar_bits_id; // @[SpectrometerTest.scala 119:30]
  wire [29:0] plfg_mux_0_auto_register_in_ar_bits_addr; // @[SpectrometerTest.scala 119:30]
  wire [2:0] plfg_mux_0_auto_register_in_ar_bits_size; // @[SpectrometerTest.scala 119:30]
  wire  plfg_mux_0_auto_register_in_r_ready; // @[SpectrometerTest.scala 119:30]
  wire  plfg_mux_0_auto_register_in_r_valid; // @[SpectrometerTest.scala 119:30]
  wire  plfg_mux_0_auto_register_in_r_bits_id; // @[SpectrometerTest.scala 119:30]
  wire [31:0] plfg_mux_0_auto_register_in_r_bits_data; // @[SpectrometerTest.scala 119:30]
  wire  plfg_mux_0_auto_stream_in_2_ready; // @[SpectrometerTest.scala 119:30]
  wire  plfg_mux_0_auto_stream_in_2_valid; // @[SpectrometerTest.scala 119:30]
  wire [31:0] plfg_mux_0_auto_stream_in_2_bits_data; // @[SpectrometerTest.scala 119:30]
  wire  plfg_mux_0_auto_stream_in_2_bits_last; // @[SpectrometerTest.scala 119:30]
  wire  plfg_mux_0_auto_stream_in_1_ready; // @[SpectrometerTest.scala 119:30]
  wire  plfg_mux_0_auto_stream_in_1_valid; // @[SpectrometerTest.scala 119:30]
  wire [31:0] plfg_mux_0_auto_stream_in_1_bits_data; // @[SpectrometerTest.scala 119:30]
  wire  plfg_mux_0_auto_stream_in_1_bits_last; // @[SpectrometerTest.scala 119:30]
  wire  plfg_mux_0_auto_stream_in_0_ready; // @[SpectrometerTest.scala 119:30]
  wire  plfg_mux_0_auto_stream_in_0_valid; // @[SpectrometerTest.scala 119:30]
  wire [31:0] plfg_mux_0_auto_stream_in_0_bits_data; // @[SpectrometerTest.scala 119:30]
  wire  plfg_mux_0_auto_stream_in_0_bits_last; // @[SpectrometerTest.scala 119:30]
  wire  plfg_mux_0_auto_stream_out_0_ready; // @[SpectrometerTest.scala 119:30]
  wire  plfg_mux_0_auto_stream_out_0_valid; // @[SpectrometerTest.scala 119:30]
  wire [31:0] plfg_mux_0_auto_stream_out_0_bits_data; // @[SpectrometerTest.scala 119:30]
  wire  plfg_mux_0_auto_stream_out_0_bits_last; // @[SpectrometerTest.scala 119:30]
  wire  plfg_mux_1_clock; // @[SpectrometerTest.scala 120:30]
  wire  plfg_mux_1_reset; // @[SpectrometerTest.scala 120:30]
  wire  plfg_mux_1_auto_register_in_aw_ready; // @[SpectrometerTest.scala 120:30]
  wire  plfg_mux_1_auto_register_in_aw_valid; // @[SpectrometerTest.scala 120:30]
  wire  plfg_mux_1_auto_register_in_aw_bits_id; // @[SpectrometerTest.scala 120:30]
  wire [29:0] plfg_mux_1_auto_register_in_aw_bits_addr; // @[SpectrometerTest.scala 120:30]
  wire  plfg_mux_1_auto_register_in_w_ready; // @[SpectrometerTest.scala 120:30]
  wire  plfg_mux_1_auto_register_in_w_valid; // @[SpectrometerTest.scala 120:30]
  wire [31:0] plfg_mux_1_auto_register_in_w_bits_data; // @[SpectrometerTest.scala 120:30]
  wire [3:0] plfg_mux_1_auto_register_in_w_bits_strb; // @[SpectrometerTest.scala 120:30]
  wire  plfg_mux_1_auto_register_in_b_ready; // @[SpectrometerTest.scala 120:30]
  wire  plfg_mux_1_auto_register_in_b_valid; // @[SpectrometerTest.scala 120:30]
  wire  plfg_mux_1_auto_register_in_b_bits_id; // @[SpectrometerTest.scala 120:30]
  wire  plfg_mux_1_auto_register_in_ar_ready; // @[SpectrometerTest.scala 120:30]
  wire  plfg_mux_1_auto_register_in_ar_valid; // @[SpectrometerTest.scala 120:30]
  wire  plfg_mux_1_auto_register_in_ar_bits_id; // @[SpectrometerTest.scala 120:30]
  wire [29:0] plfg_mux_1_auto_register_in_ar_bits_addr; // @[SpectrometerTest.scala 120:30]
  wire [2:0] plfg_mux_1_auto_register_in_ar_bits_size; // @[SpectrometerTest.scala 120:30]
  wire  plfg_mux_1_auto_register_in_r_ready; // @[SpectrometerTest.scala 120:30]
  wire  plfg_mux_1_auto_register_in_r_valid; // @[SpectrometerTest.scala 120:30]
  wire  plfg_mux_1_auto_register_in_r_bits_id; // @[SpectrometerTest.scala 120:30]
  wire [31:0] plfg_mux_1_auto_register_in_r_bits_data; // @[SpectrometerTest.scala 120:30]
  wire  plfg_mux_1_auto_stream_in_ready; // @[SpectrometerTest.scala 120:30]
  wire  plfg_mux_1_auto_stream_in_valid; // @[SpectrometerTest.scala 120:30]
  wire [31:0] plfg_mux_1_auto_stream_in_bits_data; // @[SpectrometerTest.scala 120:30]
  wire  plfg_mux_1_auto_stream_in_bits_last; // @[SpectrometerTest.scala 120:30]
  wire  plfg_mux_1_auto_stream_out_1_ready; // @[SpectrometerTest.scala 120:30]
  wire  plfg_mux_1_auto_stream_out_1_valid; // @[SpectrometerTest.scala 120:30]
  wire [31:0] plfg_mux_1_auto_stream_out_1_bits_data; // @[SpectrometerTest.scala 120:30]
  wire  plfg_mux_1_auto_stream_out_1_bits_last; // @[SpectrometerTest.scala 120:30]
  wire  nco_clock; // @[SpectrometerTest.scala 126:29]
  wire  nco_reset; // @[SpectrometerTest.scala 126:29]
  wire  nco_auto_stream_out_ready; // @[SpectrometerTest.scala 126:29]
  wire  nco_auto_stream_out_valid; // @[SpectrometerTest.scala 126:29]
  wire [31:0] nco_auto_stream_out_bits_data; // @[SpectrometerTest.scala 126:29]
  wire  nco_auto_stream_out_bits_last; // @[SpectrometerTest.scala 126:29]
  wire  nco_auto_freq_in_ready; // @[SpectrometerTest.scala 126:29]
  wire  nco_auto_freq_in_valid; // @[SpectrometerTest.scala 126:29]
  wire [31:0] nco_auto_freq_in_bits_data; // @[SpectrometerTest.scala 126:29]
  wire  nco_auto_freq_in_bits_last; // @[SpectrometerTest.scala 126:29]
  wire  nco_split_clock; // @[SpectrometerTest.scala 127:29]
  wire  nco_split_reset; // @[SpectrometerTest.scala 127:29]
  wire  nco_split_auto_mem_in_aw_ready; // @[SpectrometerTest.scala 127:29]
  wire  nco_split_auto_mem_in_aw_valid; // @[SpectrometerTest.scala 127:29]
  wire  nco_split_auto_mem_in_aw_bits_id; // @[SpectrometerTest.scala 127:29]
  wire [29:0] nco_split_auto_mem_in_aw_bits_addr; // @[SpectrometerTest.scala 127:29]
  wire  nco_split_auto_mem_in_w_ready; // @[SpectrometerTest.scala 127:29]
  wire  nco_split_auto_mem_in_w_valid; // @[SpectrometerTest.scala 127:29]
  wire [31:0] nco_split_auto_mem_in_w_bits_data; // @[SpectrometerTest.scala 127:29]
  wire [3:0] nco_split_auto_mem_in_w_bits_strb; // @[SpectrometerTest.scala 127:29]
  wire  nco_split_auto_mem_in_b_ready; // @[SpectrometerTest.scala 127:29]
  wire  nco_split_auto_mem_in_b_valid; // @[SpectrometerTest.scala 127:29]
  wire  nco_split_auto_mem_in_b_bits_id; // @[SpectrometerTest.scala 127:29]
  wire  nco_split_auto_mem_in_ar_ready; // @[SpectrometerTest.scala 127:29]
  wire  nco_split_auto_mem_in_ar_valid; // @[SpectrometerTest.scala 127:29]
  wire  nco_split_auto_mem_in_ar_bits_id; // @[SpectrometerTest.scala 127:29]
  wire [29:0] nco_split_auto_mem_in_ar_bits_addr; // @[SpectrometerTest.scala 127:29]
  wire [2:0] nco_split_auto_mem_in_ar_bits_size; // @[SpectrometerTest.scala 127:29]
  wire  nco_split_auto_mem_in_r_ready; // @[SpectrometerTest.scala 127:29]
  wire  nco_split_auto_mem_in_r_valid; // @[SpectrometerTest.scala 127:29]
  wire  nco_split_auto_mem_in_r_bits_id; // @[SpectrometerTest.scala 127:29]
  wire [31:0] nco_split_auto_mem_in_r_bits_data; // @[SpectrometerTest.scala 127:29]
  wire  nco_split_auto_stream_in_ready; // @[SpectrometerTest.scala 127:29]
  wire  nco_split_auto_stream_in_valid; // @[SpectrometerTest.scala 127:29]
  wire [31:0] nco_split_auto_stream_in_bits_data; // @[SpectrometerTest.scala 127:29]
  wire  nco_split_auto_stream_in_bits_last; // @[SpectrometerTest.scala 127:29]
  wire  nco_split_auto_stream_out_1_ready; // @[SpectrometerTest.scala 127:29]
  wire  nco_split_auto_stream_out_1_valid; // @[SpectrometerTest.scala 127:29]
  wire [31:0] nco_split_auto_stream_out_1_bits_data; // @[SpectrometerTest.scala 127:29]
  wire  nco_split_auto_stream_out_1_bits_last; // @[SpectrometerTest.scala 127:29]
  wire  nco_split_auto_stream_out_0_ready; // @[SpectrometerTest.scala 127:29]
  wire  nco_split_auto_stream_out_0_valid; // @[SpectrometerTest.scala 127:29]
  wire [31:0] nco_split_auto_stream_out_0_bits_data; // @[SpectrometerTest.scala 127:29]
  wire  nco_split_auto_stream_out_0_bits_last; // @[SpectrometerTest.scala 127:29]
  wire  nco_mux_0_clock; // @[SpectrometerTest.scala 128:29]
  wire  nco_mux_0_reset; // @[SpectrometerTest.scala 128:29]
  wire  nco_mux_0_auto_register_in_aw_ready; // @[SpectrometerTest.scala 128:29]
  wire  nco_mux_0_auto_register_in_aw_valid; // @[SpectrometerTest.scala 128:29]
  wire  nco_mux_0_auto_register_in_aw_bits_id; // @[SpectrometerTest.scala 128:29]
  wire [29:0] nco_mux_0_auto_register_in_aw_bits_addr; // @[SpectrometerTest.scala 128:29]
  wire  nco_mux_0_auto_register_in_w_ready; // @[SpectrometerTest.scala 128:29]
  wire  nco_mux_0_auto_register_in_w_valid; // @[SpectrometerTest.scala 128:29]
  wire [31:0] nco_mux_0_auto_register_in_w_bits_data; // @[SpectrometerTest.scala 128:29]
  wire [3:0] nco_mux_0_auto_register_in_w_bits_strb; // @[SpectrometerTest.scala 128:29]
  wire  nco_mux_0_auto_register_in_b_ready; // @[SpectrometerTest.scala 128:29]
  wire  nco_mux_0_auto_register_in_b_valid; // @[SpectrometerTest.scala 128:29]
  wire  nco_mux_0_auto_register_in_b_bits_id; // @[SpectrometerTest.scala 128:29]
  wire  nco_mux_0_auto_register_in_ar_ready; // @[SpectrometerTest.scala 128:29]
  wire  nco_mux_0_auto_register_in_ar_valid; // @[SpectrometerTest.scala 128:29]
  wire  nco_mux_0_auto_register_in_ar_bits_id; // @[SpectrometerTest.scala 128:29]
  wire [29:0] nco_mux_0_auto_register_in_ar_bits_addr; // @[SpectrometerTest.scala 128:29]
  wire [2:0] nco_mux_0_auto_register_in_ar_bits_size; // @[SpectrometerTest.scala 128:29]
  wire  nco_mux_0_auto_register_in_r_ready; // @[SpectrometerTest.scala 128:29]
  wire  nco_mux_0_auto_register_in_r_valid; // @[SpectrometerTest.scala 128:29]
  wire  nco_mux_0_auto_register_in_r_bits_id; // @[SpectrometerTest.scala 128:29]
  wire [31:0] nco_mux_0_auto_register_in_r_bits_data; // @[SpectrometerTest.scala 128:29]
  wire  nco_mux_0_auto_stream_in_2_ready; // @[SpectrometerTest.scala 128:29]
  wire  nco_mux_0_auto_stream_in_2_valid; // @[SpectrometerTest.scala 128:29]
  wire [31:0] nco_mux_0_auto_stream_in_2_bits_data; // @[SpectrometerTest.scala 128:29]
  wire  nco_mux_0_auto_stream_in_2_bits_last; // @[SpectrometerTest.scala 128:29]
  wire  nco_mux_0_auto_stream_in_1_ready; // @[SpectrometerTest.scala 128:29]
  wire  nco_mux_0_auto_stream_in_1_valid; // @[SpectrometerTest.scala 128:29]
  wire [31:0] nco_mux_0_auto_stream_in_1_bits_data; // @[SpectrometerTest.scala 128:29]
  wire  nco_mux_0_auto_stream_in_1_bits_last; // @[SpectrometerTest.scala 128:29]
  wire  nco_mux_0_auto_stream_in_0_ready; // @[SpectrometerTest.scala 128:29]
  wire  nco_mux_0_auto_stream_in_0_valid; // @[SpectrometerTest.scala 128:29]
  wire [31:0] nco_mux_0_auto_stream_in_0_bits_data; // @[SpectrometerTest.scala 128:29]
  wire  nco_mux_0_auto_stream_in_0_bits_last; // @[SpectrometerTest.scala 128:29]
  wire  nco_mux_0_auto_stream_out_0_ready; // @[SpectrometerTest.scala 128:29]
  wire  nco_mux_0_auto_stream_out_0_valid; // @[SpectrometerTest.scala 128:29]
  wire [31:0] nco_mux_0_auto_stream_out_0_bits_data; // @[SpectrometerTest.scala 128:29]
  wire  nco_mux_0_auto_stream_out_0_bits_last; // @[SpectrometerTest.scala 128:29]
  wire  nco_mux_1_clock; // @[SpectrometerTest.scala 129:29]
  wire  nco_mux_1_reset; // @[SpectrometerTest.scala 129:29]
  wire  nco_mux_1_auto_register_in_aw_ready; // @[SpectrometerTest.scala 129:29]
  wire  nco_mux_1_auto_register_in_aw_valid; // @[SpectrometerTest.scala 129:29]
  wire  nco_mux_1_auto_register_in_aw_bits_id; // @[SpectrometerTest.scala 129:29]
  wire [29:0] nco_mux_1_auto_register_in_aw_bits_addr; // @[SpectrometerTest.scala 129:29]
  wire  nco_mux_1_auto_register_in_w_ready; // @[SpectrometerTest.scala 129:29]
  wire  nco_mux_1_auto_register_in_w_valid; // @[SpectrometerTest.scala 129:29]
  wire [31:0] nco_mux_1_auto_register_in_w_bits_data; // @[SpectrometerTest.scala 129:29]
  wire [3:0] nco_mux_1_auto_register_in_w_bits_strb; // @[SpectrometerTest.scala 129:29]
  wire  nco_mux_1_auto_register_in_b_ready; // @[SpectrometerTest.scala 129:29]
  wire  nco_mux_1_auto_register_in_b_valid; // @[SpectrometerTest.scala 129:29]
  wire  nco_mux_1_auto_register_in_b_bits_id; // @[SpectrometerTest.scala 129:29]
  wire  nco_mux_1_auto_register_in_ar_ready; // @[SpectrometerTest.scala 129:29]
  wire  nco_mux_1_auto_register_in_ar_valid; // @[SpectrometerTest.scala 129:29]
  wire  nco_mux_1_auto_register_in_ar_bits_id; // @[SpectrometerTest.scala 129:29]
  wire [29:0] nco_mux_1_auto_register_in_ar_bits_addr; // @[SpectrometerTest.scala 129:29]
  wire [2:0] nco_mux_1_auto_register_in_ar_bits_size; // @[SpectrometerTest.scala 129:29]
  wire  nco_mux_1_auto_register_in_r_ready; // @[SpectrometerTest.scala 129:29]
  wire  nco_mux_1_auto_register_in_r_valid; // @[SpectrometerTest.scala 129:29]
  wire  nco_mux_1_auto_register_in_r_bits_id; // @[SpectrometerTest.scala 129:29]
  wire [31:0] nco_mux_1_auto_register_in_r_bits_data; // @[SpectrometerTest.scala 129:29]
  wire  nco_mux_1_auto_stream_in_ready; // @[SpectrometerTest.scala 129:29]
  wire  nco_mux_1_auto_stream_in_valid; // @[SpectrometerTest.scala 129:29]
  wire [31:0] nco_mux_1_auto_stream_in_bits_data; // @[SpectrometerTest.scala 129:29]
  wire  nco_mux_1_auto_stream_in_bits_last; // @[SpectrometerTest.scala 129:29]
  wire  nco_mux_1_auto_stream_out_1_ready; // @[SpectrometerTest.scala 129:29]
  wire  nco_mux_1_auto_stream_out_1_valid; // @[SpectrometerTest.scala 129:29]
  wire [31:0] nco_mux_1_auto_stream_out_1_bits_data; // @[SpectrometerTest.scala 129:29]
  wire  nco_mux_1_auto_stream_out_1_bits_last; // @[SpectrometerTest.scala 129:29]
  wire  fft_clock; // @[SpectrometerTest.scala 135:29]
  wire  fft_reset; // @[SpectrometerTest.scala 135:29]
  wire  fft_auto_mem_in_aw_ready; // @[SpectrometerTest.scala 135:29]
  wire  fft_auto_mem_in_aw_valid; // @[SpectrometerTest.scala 135:29]
  wire  fft_auto_mem_in_aw_bits_id; // @[SpectrometerTest.scala 135:29]
  wire [29:0] fft_auto_mem_in_aw_bits_addr; // @[SpectrometerTest.scala 135:29]
  wire  fft_auto_mem_in_w_ready; // @[SpectrometerTest.scala 135:29]
  wire  fft_auto_mem_in_w_valid; // @[SpectrometerTest.scala 135:29]
  wire [31:0] fft_auto_mem_in_w_bits_data; // @[SpectrometerTest.scala 135:29]
  wire [3:0] fft_auto_mem_in_w_bits_strb; // @[SpectrometerTest.scala 135:29]
  wire  fft_auto_mem_in_b_ready; // @[SpectrometerTest.scala 135:29]
  wire  fft_auto_mem_in_b_valid; // @[SpectrometerTest.scala 135:29]
  wire  fft_auto_mem_in_b_bits_id; // @[SpectrometerTest.scala 135:29]
  wire  fft_auto_mem_in_ar_ready; // @[SpectrometerTest.scala 135:29]
  wire  fft_auto_mem_in_ar_valid; // @[SpectrometerTest.scala 135:29]
  wire  fft_auto_mem_in_ar_bits_id; // @[SpectrometerTest.scala 135:29]
  wire [29:0] fft_auto_mem_in_ar_bits_addr; // @[SpectrometerTest.scala 135:29]
  wire [2:0] fft_auto_mem_in_ar_bits_size; // @[SpectrometerTest.scala 135:29]
  wire  fft_auto_mem_in_r_ready; // @[SpectrometerTest.scala 135:29]
  wire  fft_auto_mem_in_r_valid; // @[SpectrometerTest.scala 135:29]
  wire  fft_auto_mem_in_r_bits_id; // @[SpectrometerTest.scala 135:29]
  wire [31:0] fft_auto_mem_in_r_bits_data; // @[SpectrometerTest.scala 135:29]
  wire  fft_auto_stream_in_ready; // @[SpectrometerTest.scala 135:29]
  wire  fft_auto_stream_in_valid; // @[SpectrometerTest.scala 135:29]
  wire [31:0] fft_auto_stream_in_bits_data; // @[SpectrometerTest.scala 135:29]
  wire  fft_auto_stream_in_bits_last; // @[SpectrometerTest.scala 135:29]
  wire  fft_auto_stream_out_ready; // @[SpectrometerTest.scala 135:29]
  wire  fft_auto_stream_out_valid; // @[SpectrometerTest.scala 135:29]
  wire [31:0] fft_auto_stream_out_bits_data; // @[SpectrometerTest.scala 135:29]
  wire  fft_auto_stream_out_bits_last; // @[SpectrometerTest.scala 135:29]
  wire  fft_split_clock; // @[SpectrometerTest.scala 136:29]
  wire  fft_split_reset; // @[SpectrometerTest.scala 136:29]
  wire  fft_split_auto_mem_in_aw_ready; // @[SpectrometerTest.scala 136:29]
  wire  fft_split_auto_mem_in_aw_valid; // @[SpectrometerTest.scala 136:29]
  wire  fft_split_auto_mem_in_aw_bits_id; // @[SpectrometerTest.scala 136:29]
  wire [29:0] fft_split_auto_mem_in_aw_bits_addr; // @[SpectrometerTest.scala 136:29]
  wire  fft_split_auto_mem_in_w_ready; // @[SpectrometerTest.scala 136:29]
  wire  fft_split_auto_mem_in_w_valid; // @[SpectrometerTest.scala 136:29]
  wire [31:0] fft_split_auto_mem_in_w_bits_data; // @[SpectrometerTest.scala 136:29]
  wire [3:0] fft_split_auto_mem_in_w_bits_strb; // @[SpectrometerTest.scala 136:29]
  wire  fft_split_auto_mem_in_b_ready; // @[SpectrometerTest.scala 136:29]
  wire  fft_split_auto_mem_in_b_valid; // @[SpectrometerTest.scala 136:29]
  wire  fft_split_auto_mem_in_b_bits_id; // @[SpectrometerTest.scala 136:29]
  wire  fft_split_auto_mem_in_ar_ready; // @[SpectrometerTest.scala 136:29]
  wire  fft_split_auto_mem_in_ar_valid; // @[SpectrometerTest.scala 136:29]
  wire  fft_split_auto_mem_in_ar_bits_id; // @[SpectrometerTest.scala 136:29]
  wire [29:0] fft_split_auto_mem_in_ar_bits_addr; // @[SpectrometerTest.scala 136:29]
  wire [2:0] fft_split_auto_mem_in_ar_bits_size; // @[SpectrometerTest.scala 136:29]
  wire  fft_split_auto_mem_in_r_ready; // @[SpectrometerTest.scala 136:29]
  wire  fft_split_auto_mem_in_r_valid; // @[SpectrometerTest.scala 136:29]
  wire  fft_split_auto_mem_in_r_bits_id; // @[SpectrometerTest.scala 136:29]
  wire [31:0] fft_split_auto_mem_in_r_bits_data; // @[SpectrometerTest.scala 136:29]
  wire  fft_split_auto_stream_in_ready; // @[SpectrometerTest.scala 136:29]
  wire  fft_split_auto_stream_in_valid; // @[SpectrometerTest.scala 136:29]
  wire [31:0] fft_split_auto_stream_in_bits_data; // @[SpectrometerTest.scala 136:29]
  wire  fft_split_auto_stream_in_bits_last; // @[SpectrometerTest.scala 136:29]
  wire  fft_split_auto_stream_out_1_ready; // @[SpectrometerTest.scala 136:29]
  wire  fft_split_auto_stream_out_1_valid; // @[SpectrometerTest.scala 136:29]
  wire [31:0] fft_split_auto_stream_out_1_bits_data; // @[SpectrometerTest.scala 136:29]
  wire  fft_split_auto_stream_out_1_bits_last; // @[SpectrometerTest.scala 136:29]
  wire  fft_split_auto_stream_out_0_ready; // @[SpectrometerTest.scala 136:29]
  wire  fft_split_auto_stream_out_0_valid; // @[SpectrometerTest.scala 136:29]
  wire [31:0] fft_split_auto_stream_out_0_bits_data; // @[SpectrometerTest.scala 136:29]
  wire  fft_split_auto_stream_out_0_bits_last; // @[SpectrometerTest.scala 136:29]
  wire  fft_mux_0_clock; // @[SpectrometerTest.scala 137:29]
  wire  fft_mux_0_reset; // @[SpectrometerTest.scala 137:29]
  wire  fft_mux_0_auto_register_in_aw_ready; // @[SpectrometerTest.scala 137:29]
  wire  fft_mux_0_auto_register_in_aw_valid; // @[SpectrometerTest.scala 137:29]
  wire  fft_mux_0_auto_register_in_aw_bits_id; // @[SpectrometerTest.scala 137:29]
  wire [29:0] fft_mux_0_auto_register_in_aw_bits_addr; // @[SpectrometerTest.scala 137:29]
  wire  fft_mux_0_auto_register_in_w_ready; // @[SpectrometerTest.scala 137:29]
  wire  fft_mux_0_auto_register_in_w_valid; // @[SpectrometerTest.scala 137:29]
  wire [31:0] fft_mux_0_auto_register_in_w_bits_data; // @[SpectrometerTest.scala 137:29]
  wire [3:0] fft_mux_0_auto_register_in_w_bits_strb; // @[SpectrometerTest.scala 137:29]
  wire  fft_mux_0_auto_register_in_b_ready; // @[SpectrometerTest.scala 137:29]
  wire  fft_mux_0_auto_register_in_b_valid; // @[SpectrometerTest.scala 137:29]
  wire  fft_mux_0_auto_register_in_b_bits_id; // @[SpectrometerTest.scala 137:29]
  wire  fft_mux_0_auto_register_in_ar_ready; // @[SpectrometerTest.scala 137:29]
  wire  fft_mux_0_auto_register_in_ar_valid; // @[SpectrometerTest.scala 137:29]
  wire  fft_mux_0_auto_register_in_ar_bits_id; // @[SpectrometerTest.scala 137:29]
  wire [29:0] fft_mux_0_auto_register_in_ar_bits_addr; // @[SpectrometerTest.scala 137:29]
  wire [2:0] fft_mux_0_auto_register_in_ar_bits_size; // @[SpectrometerTest.scala 137:29]
  wire  fft_mux_0_auto_register_in_r_ready; // @[SpectrometerTest.scala 137:29]
  wire  fft_mux_0_auto_register_in_r_valid; // @[SpectrometerTest.scala 137:29]
  wire  fft_mux_0_auto_register_in_r_bits_id; // @[SpectrometerTest.scala 137:29]
  wire [31:0] fft_mux_0_auto_register_in_r_bits_data; // @[SpectrometerTest.scala 137:29]
  wire  fft_mux_0_auto_stream_in_2_ready; // @[SpectrometerTest.scala 137:29]
  wire  fft_mux_0_auto_stream_in_2_valid; // @[SpectrometerTest.scala 137:29]
  wire [31:0] fft_mux_0_auto_stream_in_2_bits_data; // @[SpectrometerTest.scala 137:29]
  wire  fft_mux_0_auto_stream_in_2_bits_last; // @[SpectrometerTest.scala 137:29]
  wire  fft_mux_0_auto_stream_in_1_ready; // @[SpectrometerTest.scala 137:29]
  wire  fft_mux_0_auto_stream_in_1_valid; // @[SpectrometerTest.scala 137:29]
  wire [31:0] fft_mux_0_auto_stream_in_1_bits_data; // @[SpectrometerTest.scala 137:29]
  wire  fft_mux_0_auto_stream_in_1_bits_last; // @[SpectrometerTest.scala 137:29]
  wire  fft_mux_0_auto_stream_in_0_ready; // @[SpectrometerTest.scala 137:29]
  wire  fft_mux_0_auto_stream_in_0_valid; // @[SpectrometerTest.scala 137:29]
  wire [31:0] fft_mux_0_auto_stream_in_0_bits_data; // @[SpectrometerTest.scala 137:29]
  wire  fft_mux_0_auto_stream_in_0_bits_last; // @[SpectrometerTest.scala 137:29]
  wire  fft_mux_0_auto_stream_out_0_ready; // @[SpectrometerTest.scala 137:29]
  wire  fft_mux_0_auto_stream_out_0_valid; // @[SpectrometerTest.scala 137:29]
  wire [31:0] fft_mux_0_auto_stream_out_0_bits_data; // @[SpectrometerTest.scala 137:29]
  wire  fft_mux_0_auto_stream_out_0_bits_last; // @[SpectrometerTest.scala 137:29]
  wire  fft_mux_1_clock; // @[SpectrometerTest.scala 138:29]
  wire  fft_mux_1_reset; // @[SpectrometerTest.scala 138:29]
  wire  fft_mux_1_auto_register_in_aw_ready; // @[SpectrometerTest.scala 138:29]
  wire  fft_mux_1_auto_register_in_aw_valid; // @[SpectrometerTest.scala 138:29]
  wire  fft_mux_1_auto_register_in_aw_bits_id; // @[SpectrometerTest.scala 138:29]
  wire [29:0] fft_mux_1_auto_register_in_aw_bits_addr; // @[SpectrometerTest.scala 138:29]
  wire  fft_mux_1_auto_register_in_w_ready; // @[SpectrometerTest.scala 138:29]
  wire  fft_mux_1_auto_register_in_w_valid; // @[SpectrometerTest.scala 138:29]
  wire [31:0] fft_mux_1_auto_register_in_w_bits_data; // @[SpectrometerTest.scala 138:29]
  wire [3:0] fft_mux_1_auto_register_in_w_bits_strb; // @[SpectrometerTest.scala 138:29]
  wire  fft_mux_1_auto_register_in_b_ready; // @[SpectrometerTest.scala 138:29]
  wire  fft_mux_1_auto_register_in_b_valid; // @[SpectrometerTest.scala 138:29]
  wire  fft_mux_1_auto_register_in_b_bits_id; // @[SpectrometerTest.scala 138:29]
  wire  fft_mux_1_auto_register_in_ar_ready; // @[SpectrometerTest.scala 138:29]
  wire  fft_mux_1_auto_register_in_ar_valid; // @[SpectrometerTest.scala 138:29]
  wire  fft_mux_1_auto_register_in_ar_bits_id; // @[SpectrometerTest.scala 138:29]
  wire [29:0] fft_mux_1_auto_register_in_ar_bits_addr; // @[SpectrometerTest.scala 138:29]
  wire [2:0] fft_mux_1_auto_register_in_ar_bits_size; // @[SpectrometerTest.scala 138:29]
  wire  fft_mux_1_auto_register_in_r_ready; // @[SpectrometerTest.scala 138:29]
  wire  fft_mux_1_auto_register_in_r_valid; // @[SpectrometerTest.scala 138:29]
  wire  fft_mux_1_auto_register_in_r_bits_id; // @[SpectrometerTest.scala 138:29]
  wire [31:0] fft_mux_1_auto_register_in_r_bits_data; // @[SpectrometerTest.scala 138:29]
  wire  fft_mux_1_auto_stream_in_ready; // @[SpectrometerTest.scala 138:29]
  wire  fft_mux_1_auto_stream_in_valid; // @[SpectrometerTest.scala 138:29]
  wire [31:0] fft_mux_1_auto_stream_in_bits_data; // @[SpectrometerTest.scala 138:29]
  wire  fft_mux_1_auto_stream_in_bits_last; // @[SpectrometerTest.scala 138:29]
  wire  fft_mux_1_auto_stream_out_1_ready; // @[SpectrometerTest.scala 138:29]
  wire  fft_mux_1_auto_stream_out_1_valid; // @[SpectrometerTest.scala 138:29]
  wire [31:0] fft_mux_1_auto_stream_out_1_bits_data; // @[SpectrometerTest.scala 138:29]
  wire  fft_mux_1_auto_stream_out_1_bits_last; // @[SpectrometerTest.scala 138:29]
  wire  mag_clock; // @[SpectrometerTest.scala 144:29]
  wire  mag_reset; // @[SpectrometerTest.scala 144:29]
  wire  mag_auto_mem_in_aw_ready; // @[SpectrometerTest.scala 144:29]
  wire  mag_auto_mem_in_aw_valid; // @[SpectrometerTest.scala 144:29]
  wire  mag_auto_mem_in_aw_bits_id; // @[SpectrometerTest.scala 144:29]
  wire [29:0] mag_auto_mem_in_aw_bits_addr; // @[SpectrometerTest.scala 144:29]
  wire  mag_auto_mem_in_w_ready; // @[SpectrometerTest.scala 144:29]
  wire  mag_auto_mem_in_w_valid; // @[SpectrometerTest.scala 144:29]
  wire [31:0] mag_auto_mem_in_w_bits_data; // @[SpectrometerTest.scala 144:29]
  wire [3:0] mag_auto_mem_in_w_bits_strb; // @[SpectrometerTest.scala 144:29]
  wire  mag_auto_mem_in_b_ready; // @[SpectrometerTest.scala 144:29]
  wire  mag_auto_mem_in_b_valid; // @[SpectrometerTest.scala 144:29]
  wire  mag_auto_mem_in_b_bits_id; // @[SpectrometerTest.scala 144:29]
  wire  mag_auto_mem_in_ar_ready; // @[SpectrometerTest.scala 144:29]
  wire  mag_auto_mem_in_ar_valid; // @[SpectrometerTest.scala 144:29]
  wire  mag_auto_mem_in_ar_bits_id; // @[SpectrometerTest.scala 144:29]
  wire [29:0] mag_auto_mem_in_ar_bits_addr; // @[SpectrometerTest.scala 144:29]
  wire [2:0] mag_auto_mem_in_ar_bits_size; // @[SpectrometerTest.scala 144:29]
  wire  mag_auto_mem_in_r_ready; // @[SpectrometerTest.scala 144:29]
  wire  mag_auto_mem_in_r_valid; // @[SpectrometerTest.scala 144:29]
  wire  mag_auto_mem_in_r_bits_id; // @[SpectrometerTest.scala 144:29]
  wire [31:0] mag_auto_mem_in_r_bits_data; // @[SpectrometerTest.scala 144:29]
  wire  mag_auto_stream_in_ready; // @[SpectrometerTest.scala 144:29]
  wire  mag_auto_stream_in_valid; // @[SpectrometerTest.scala 144:29]
  wire [31:0] mag_auto_stream_in_bits_data; // @[SpectrometerTest.scala 144:29]
  wire  mag_auto_stream_in_bits_last; // @[SpectrometerTest.scala 144:29]
  wire  mag_auto_stream_out_ready; // @[SpectrometerTest.scala 144:29]
  wire  mag_auto_stream_out_valid; // @[SpectrometerTest.scala 144:29]
  wire [31:0] mag_auto_stream_out_bits_data; // @[SpectrometerTest.scala 144:29]
  wire  mag_auto_stream_out_bits_last; // @[SpectrometerTest.scala 144:29]
  wire  mag_split_clock; // @[SpectrometerTest.scala 145:29]
  wire  mag_split_reset; // @[SpectrometerTest.scala 145:29]
  wire  mag_split_auto_mem_in_aw_ready; // @[SpectrometerTest.scala 145:29]
  wire  mag_split_auto_mem_in_aw_valid; // @[SpectrometerTest.scala 145:29]
  wire  mag_split_auto_mem_in_aw_bits_id; // @[SpectrometerTest.scala 145:29]
  wire [29:0] mag_split_auto_mem_in_aw_bits_addr; // @[SpectrometerTest.scala 145:29]
  wire  mag_split_auto_mem_in_w_ready; // @[SpectrometerTest.scala 145:29]
  wire  mag_split_auto_mem_in_w_valid; // @[SpectrometerTest.scala 145:29]
  wire [31:0] mag_split_auto_mem_in_w_bits_data; // @[SpectrometerTest.scala 145:29]
  wire [3:0] mag_split_auto_mem_in_w_bits_strb; // @[SpectrometerTest.scala 145:29]
  wire  mag_split_auto_mem_in_b_ready; // @[SpectrometerTest.scala 145:29]
  wire  mag_split_auto_mem_in_b_valid; // @[SpectrometerTest.scala 145:29]
  wire  mag_split_auto_mem_in_b_bits_id; // @[SpectrometerTest.scala 145:29]
  wire  mag_split_auto_mem_in_ar_ready; // @[SpectrometerTest.scala 145:29]
  wire  mag_split_auto_mem_in_ar_valid; // @[SpectrometerTest.scala 145:29]
  wire  mag_split_auto_mem_in_ar_bits_id; // @[SpectrometerTest.scala 145:29]
  wire [29:0] mag_split_auto_mem_in_ar_bits_addr; // @[SpectrometerTest.scala 145:29]
  wire [2:0] mag_split_auto_mem_in_ar_bits_size; // @[SpectrometerTest.scala 145:29]
  wire  mag_split_auto_mem_in_r_ready; // @[SpectrometerTest.scala 145:29]
  wire  mag_split_auto_mem_in_r_valid; // @[SpectrometerTest.scala 145:29]
  wire  mag_split_auto_mem_in_r_bits_id; // @[SpectrometerTest.scala 145:29]
  wire [31:0] mag_split_auto_mem_in_r_bits_data; // @[SpectrometerTest.scala 145:29]
  wire  mag_split_auto_stream_in_ready; // @[SpectrometerTest.scala 145:29]
  wire  mag_split_auto_stream_in_valid; // @[SpectrometerTest.scala 145:29]
  wire [31:0] mag_split_auto_stream_in_bits_data; // @[SpectrometerTest.scala 145:29]
  wire  mag_split_auto_stream_in_bits_last; // @[SpectrometerTest.scala 145:29]
  wire  mag_split_auto_stream_out_1_ready; // @[SpectrometerTest.scala 145:29]
  wire  mag_split_auto_stream_out_1_valid; // @[SpectrometerTest.scala 145:29]
  wire [31:0] mag_split_auto_stream_out_1_bits_data; // @[SpectrometerTest.scala 145:29]
  wire  mag_split_auto_stream_out_1_bits_last; // @[SpectrometerTest.scala 145:29]
  wire  mag_split_auto_stream_out_0_ready; // @[SpectrometerTest.scala 145:29]
  wire  mag_split_auto_stream_out_0_valid; // @[SpectrometerTest.scala 145:29]
  wire [31:0] mag_split_auto_stream_out_0_bits_data; // @[SpectrometerTest.scala 145:29]
  wire  mag_split_auto_stream_out_0_bits_last; // @[SpectrometerTest.scala 145:29]
  wire  mag_mux_0_clock; // @[SpectrometerTest.scala 146:29]
  wire  mag_mux_0_reset; // @[SpectrometerTest.scala 146:29]
  wire  mag_mux_0_auto_register_in_aw_ready; // @[SpectrometerTest.scala 146:29]
  wire  mag_mux_0_auto_register_in_aw_valid; // @[SpectrometerTest.scala 146:29]
  wire  mag_mux_0_auto_register_in_aw_bits_id; // @[SpectrometerTest.scala 146:29]
  wire [29:0] mag_mux_0_auto_register_in_aw_bits_addr; // @[SpectrometerTest.scala 146:29]
  wire  mag_mux_0_auto_register_in_w_ready; // @[SpectrometerTest.scala 146:29]
  wire  mag_mux_0_auto_register_in_w_valid; // @[SpectrometerTest.scala 146:29]
  wire [31:0] mag_mux_0_auto_register_in_w_bits_data; // @[SpectrometerTest.scala 146:29]
  wire [3:0] mag_mux_0_auto_register_in_w_bits_strb; // @[SpectrometerTest.scala 146:29]
  wire  mag_mux_0_auto_register_in_b_ready; // @[SpectrometerTest.scala 146:29]
  wire  mag_mux_0_auto_register_in_b_valid; // @[SpectrometerTest.scala 146:29]
  wire  mag_mux_0_auto_register_in_b_bits_id; // @[SpectrometerTest.scala 146:29]
  wire  mag_mux_0_auto_register_in_ar_ready; // @[SpectrometerTest.scala 146:29]
  wire  mag_mux_0_auto_register_in_ar_valid; // @[SpectrometerTest.scala 146:29]
  wire  mag_mux_0_auto_register_in_ar_bits_id; // @[SpectrometerTest.scala 146:29]
  wire [29:0] mag_mux_0_auto_register_in_ar_bits_addr; // @[SpectrometerTest.scala 146:29]
  wire [2:0] mag_mux_0_auto_register_in_ar_bits_size; // @[SpectrometerTest.scala 146:29]
  wire  mag_mux_0_auto_register_in_r_ready; // @[SpectrometerTest.scala 146:29]
  wire  mag_mux_0_auto_register_in_r_valid; // @[SpectrometerTest.scala 146:29]
  wire  mag_mux_0_auto_register_in_r_bits_id; // @[SpectrometerTest.scala 146:29]
  wire [31:0] mag_mux_0_auto_register_in_r_bits_data; // @[SpectrometerTest.scala 146:29]
  wire  mag_mux_0_auto_stream_in_2_ready; // @[SpectrometerTest.scala 146:29]
  wire  mag_mux_0_auto_stream_in_2_valid; // @[SpectrometerTest.scala 146:29]
  wire [31:0] mag_mux_0_auto_stream_in_2_bits_data; // @[SpectrometerTest.scala 146:29]
  wire  mag_mux_0_auto_stream_in_2_bits_last; // @[SpectrometerTest.scala 146:29]
  wire  mag_mux_0_auto_stream_in_1_ready; // @[SpectrometerTest.scala 146:29]
  wire  mag_mux_0_auto_stream_in_1_valid; // @[SpectrometerTest.scala 146:29]
  wire [31:0] mag_mux_0_auto_stream_in_1_bits_data; // @[SpectrometerTest.scala 146:29]
  wire  mag_mux_0_auto_stream_in_1_bits_last; // @[SpectrometerTest.scala 146:29]
  wire  mag_mux_0_auto_stream_in_0_ready; // @[SpectrometerTest.scala 146:29]
  wire  mag_mux_0_auto_stream_in_0_valid; // @[SpectrometerTest.scala 146:29]
  wire [31:0] mag_mux_0_auto_stream_in_0_bits_data; // @[SpectrometerTest.scala 146:29]
  wire  mag_mux_0_auto_stream_in_0_bits_last; // @[SpectrometerTest.scala 146:29]
  wire  mag_mux_0_auto_stream_out_0_ready; // @[SpectrometerTest.scala 146:29]
  wire  mag_mux_0_auto_stream_out_0_valid; // @[SpectrometerTest.scala 146:29]
  wire [31:0] mag_mux_0_auto_stream_out_0_bits_data; // @[SpectrometerTest.scala 146:29]
  wire  mag_mux_0_auto_stream_out_0_bits_last; // @[SpectrometerTest.scala 146:29]
  wire  mag_mux_1_clock; // @[SpectrometerTest.scala 147:29]
  wire  mag_mux_1_reset; // @[SpectrometerTest.scala 147:29]
  wire  mag_mux_1_auto_register_in_aw_ready; // @[SpectrometerTest.scala 147:29]
  wire  mag_mux_1_auto_register_in_aw_valid; // @[SpectrometerTest.scala 147:29]
  wire  mag_mux_1_auto_register_in_aw_bits_id; // @[SpectrometerTest.scala 147:29]
  wire [29:0] mag_mux_1_auto_register_in_aw_bits_addr; // @[SpectrometerTest.scala 147:29]
  wire  mag_mux_1_auto_register_in_w_ready; // @[SpectrometerTest.scala 147:29]
  wire  mag_mux_1_auto_register_in_w_valid; // @[SpectrometerTest.scala 147:29]
  wire [31:0] mag_mux_1_auto_register_in_w_bits_data; // @[SpectrometerTest.scala 147:29]
  wire [3:0] mag_mux_1_auto_register_in_w_bits_strb; // @[SpectrometerTest.scala 147:29]
  wire  mag_mux_1_auto_register_in_b_ready; // @[SpectrometerTest.scala 147:29]
  wire  mag_mux_1_auto_register_in_b_valid; // @[SpectrometerTest.scala 147:29]
  wire  mag_mux_1_auto_register_in_b_bits_id; // @[SpectrometerTest.scala 147:29]
  wire  mag_mux_1_auto_register_in_ar_ready; // @[SpectrometerTest.scala 147:29]
  wire  mag_mux_1_auto_register_in_ar_valid; // @[SpectrometerTest.scala 147:29]
  wire  mag_mux_1_auto_register_in_ar_bits_id; // @[SpectrometerTest.scala 147:29]
  wire [29:0] mag_mux_1_auto_register_in_ar_bits_addr; // @[SpectrometerTest.scala 147:29]
  wire [2:0] mag_mux_1_auto_register_in_ar_bits_size; // @[SpectrometerTest.scala 147:29]
  wire  mag_mux_1_auto_register_in_r_ready; // @[SpectrometerTest.scala 147:29]
  wire  mag_mux_1_auto_register_in_r_valid; // @[SpectrometerTest.scala 147:29]
  wire  mag_mux_1_auto_register_in_r_bits_id; // @[SpectrometerTest.scala 147:29]
  wire [31:0] mag_mux_1_auto_register_in_r_bits_data; // @[SpectrometerTest.scala 147:29]
  wire  mag_mux_1_auto_stream_in_ready; // @[SpectrometerTest.scala 147:29]
  wire  mag_mux_1_auto_stream_in_valid; // @[SpectrometerTest.scala 147:29]
  wire [31:0] mag_mux_1_auto_stream_in_bits_data; // @[SpectrometerTest.scala 147:29]
  wire  mag_mux_1_auto_stream_in_bits_last; // @[SpectrometerTest.scala 147:29]
  wire  mag_mux_1_auto_stream_out_1_ready; // @[SpectrometerTest.scala 147:29]
  wire  mag_mux_1_auto_stream_out_1_valid; // @[SpectrometerTest.scala 147:29]
  wire [31:0] mag_mux_1_auto_stream_out_1_bits_data; // @[SpectrometerTest.scala 147:29]
  wire  mag_mux_1_auto_stream_out_1_bits_last; // @[SpectrometerTest.scala 147:29]
  wire  acc_clock; // @[SpectrometerTest.scala 153:29]
  wire  acc_reset; // @[SpectrometerTest.scala 153:29]
  wire  acc_auto_bus_in_aw_ready; // @[SpectrometerTest.scala 153:29]
  wire  acc_auto_bus_in_aw_valid; // @[SpectrometerTest.scala 153:29]
  wire  acc_auto_bus_in_aw_bits_id; // @[SpectrometerTest.scala 153:29]
  wire [29:0] acc_auto_bus_in_aw_bits_addr; // @[SpectrometerTest.scala 153:29]
  wire [2:0] acc_auto_bus_in_aw_bits_size; // @[SpectrometerTest.scala 153:29]
  wire  acc_auto_bus_in_w_ready; // @[SpectrometerTest.scala 153:29]
  wire  acc_auto_bus_in_w_valid; // @[SpectrometerTest.scala 153:29]
  wire [31:0] acc_auto_bus_in_w_bits_data; // @[SpectrometerTest.scala 153:29]
  wire [3:0] acc_auto_bus_in_w_bits_strb; // @[SpectrometerTest.scala 153:29]
  wire  acc_auto_bus_in_w_bits_last; // @[SpectrometerTest.scala 153:29]
  wire  acc_auto_bus_in_b_ready; // @[SpectrometerTest.scala 153:29]
  wire  acc_auto_bus_in_b_valid; // @[SpectrometerTest.scala 153:29]
  wire [1:0] acc_auto_bus_in_b_bits_resp; // @[SpectrometerTest.scala 153:29]
  wire  acc_auto_bus_in_ar_ready; // @[SpectrometerTest.scala 153:29]
  wire  acc_auto_bus_in_ar_valid; // @[SpectrometerTest.scala 153:29]
  wire  acc_auto_bus_in_ar_bits_id; // @[SpectrometerTest.scala 153:29]
  wire [29:0] acc_auto_bus_in_ar_bits_addr; // @[SpectrometerTest.scala 153:29]
  wire [2:0] acc_auto_bus_in_ar_bits_size; // @[SpectrometerTest.scala 153:29]
  wire  acc_auto_bus_in_r_ready; // @[SpectrometerTest.scala 153:29]
  wire  acc_auto_bus_in_r_valid; // @[SpectrometerTest.scala 153:29]
  wire [31:0] acc_auto_bus_in_r_bits_data; // @[SpectrometerTest.scala 153:29]
  wire [1:0] acc_auto_bus_in_r_bits_resp; // @[SpectrometerTest.scala 153:29]
  wire  acc_auto_bus_in_r_bits_last; // @[SpectrometerTest.scala 153:29]
  wire  acc_auto_dspQueue_stream_out_ready; // @[SpectrometerTest.scala 153:29]
  wire  acc_auto_dspQueue_stream_out_valid; // @[SpectrometerTest.scala 153:29]
  wire [15:0] acc_auto_dspQueue_stream_out_bits_data; // @[SpectrometerTest.scala 153:29]
  wire  acc_auto_dspQueue_stream_out_bits_last; // @[SpectrometerTest.scala 153:29]
  wire  acc_auto_accumulator_slave_in_ready; // @[SpectrometerTest.scala 153:29]
  wire  acc_auto_accumulator_slave_in_valid; // @[SpectrometerTest.scala 153:29]
  wire [31:0] acc_auto_accumulator_slave_in_bits_data; // @[SpectrometerTest.scala 153:29]
  wire  acc_auto_accumulator_slave_in_bits_last; // @[SpectrometerTest.scala 153:29]
  wire  widthAdapter_1_clock; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_1_reset; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_1_auto_in_ready; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_1_auto_in_valid; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire [15:0] widthAdapter_1_auto_in_bits_data; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_1_auto_in_bits_last; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_1_auto_out_ready; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_1_auto_out_valid; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire [31:0] widthAdapter_1_auto_out_bits_data; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_1_auto_out_bits_last; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  acc_queue_clock; // @[SpectrometerTest.scala 155:29]
  wire  acc_queue_reset; // @[SpectrometerTest.scala 155:29]
  wire  acc_queue_auto_out_out_ready; // @[SpectrometerTest.scala 155:29]
  wire  acc_queue_auto_out_out_valid; // @[SpectrometerTest.scala 155:29]
  wire [31:0] acc_queue_auto_out_out_bits_data; // @[SpectrometerTest.scala 155:29]
  wire  acc_queue_auto_out_out_bits_last; // @[SpectrometerTest.scala 155:29]
  wire  acc_queue_auto_in_in_ready; // @[SpectrometerTest.scala 155:29]
  wire  acc_queue_auto_in_in_valid; // @[SpectrometerTest.scala 155:29]
  wire [31:0] acc_queue_auto_in_in_bits_data; // @[SpectrometerTest.scala 155:29]
  wire  acc_queue_auto_in_in_bits_last; // @[SpectrometerTest.scala 155:29]
  wire  out_mux_clock; // @[SpectrometerTest.scala 157:29]
  wire  out_mux_reset; // @[SpectrometerTest.scala 157:29]
  wire  out_mux_auto_register_in_aw_ready; // @[SpectrometerTest.scala 157:29]
  wire  out_mux_auto_register_in_aw_valid; // @[SpectrometerTest.scala 157:29]
  wire  out_mux_auto_register_in_aw_bits_id; // @[SpectrometerTest.scala 157:29]
  wire [29:0] out_mux_auto_register_in_aw_bits_addr; // @[SpectrometerTest.scala 157:29]
  wire  out_mux_auto_register_in_w_ready; // @[SpectrometerTest.scala 157:29]
  wire  out_mux_auto_register_in_w_valid; // @[SpectrometerTest.scala 157:29]
  wire [31:0] out_mux_auto_register_in_w_bits_data; // @[SpectrometerTest.scala 157:29]
  wire [3:0] out_mux_auto_register_in_w_bits_strb; // @[SpectrometerTest.scala 157:29]
  wire  out_mux_auto_register_in_b_ready; // @[SpectrometerTest.scala 157:29]
  wire  out_mux_auto_register_in_b_valid; // @[SpectrometerTest.scala 157:29]
  wire  out_mux_auto_register_in_b_bits_id; // @[SpectrometerTest.scala 157:29]
  wire  out_mux_auto_register_in_ar_ready; // @[SpectrometerTest.scala 157:29]
  wire  out_mux_auto_register_in_ar_valid; // @[SpectrometerTest.scala 157:29]
  wire  out_mux_auto_register_in_ar_bits_id; // @[SpectrometerTest.scala 157:29]
  wire [29:0] out_mux_auto_register_in_ar_bits_addr; // @[SpectrometerTest.scala 157:29]
  wire [2:0] out_mux_auto_register_in_ar_bits_size; // @[SpectrometerTest.scala 157:29]
  wire  out_mux_auto_register_in_r_ready; // @[SpectrometerTest.scala 157:29]
  wire  out_mux_auto_register_in_r_valid; // @[SpectrometerTest.scala 157:29]
  wire  out_mux_auto_register_in_r_bits_id; // @[SpectrometerTest.scala 157:29]
  wire [31:0] out_mux_auto_register_in_r_bits_data; // @[SpectrometerTest.scala 157:29]
  wire  out_mux_auto_stream_in_6_ready; // @[SpectrometerTest.scala 157:29]
  wire  out_mux_auto_stream_in_6_valid; // @[SpectrometerTest.scala 157:29]
  wire [31:0] out_mux_auto_stream_in_6_bits_data; // @[SpectrometerTest.scala 157:29]
  wire  out_mux_auto_stream_in_6_bits_last; // @[SpectrometerTest.scala 157:29]
  wire  out_mux_auto_stream_in_5_ready; // @[SpectrometerTest.scala 157:29]
  wire  out_mux_auto_stream_in_5_valid; // @[SpectrometerTest.scala 157:29]
  wire [31:0] out_mux_auto_stream_in_5_bits_data; // @[SpectrometerTest.scala 157:29]
  wire  out_mux_auto_stream_in_5_bits_last; // @[SpectrometerTest.scala 157:29]
  wire  out_mux_auto_stream_in_4_ready; // @[SpectrometerTest.scala 157:29]
  wire  out_mux_auto_stream_in_4_valid; // @[SpectrometerTest.scala 157:29]
  wire [31:0] out_mux_auto_stream_in_4_bits_data; // @[SpectrometerTest.scala 157:29]
  wire  out_mux_auto_stream_in_4_bits_last; // @[SpectrometerTest.scala 157:29]
  wire  out_mux_auto_stream_in_3_ready; // @[SpectrometerTest.scala 157:29]
  wire  out_mux_auto_stream_in_3_valid; // @[SpectrometerTest.scala 157:29]
  wire [31:0] out_mux_auto_stream_in_3_bits_data; // @[SpectrometerTest.scala 157:29]
  wire  out_mux_auto_stream_in_3_bits_last; // @[SpectrometerTest.scala 157:29]
  wire  out_mux_auto_stream_in_2_ready; // @[SpectrometerTest.scala 157:29]
  wire  out_mux_auto_stream_in_2_valid; // @[SpectrometerTest.scala 157:29]
  wire [31:0] out_mux_auto_stream_in_2_bits_data; // @[SpectrometerTest.scala 157:29]
  wire  out_mux_auto_stream_in_2_bits_last; // @[SpectrometerTest.scala 157:29]
  wire  out_mux_auto_stream_in_1_ready; // @[SpectrometerTest.scala 157:29]
  wire  out_mux_auto_stream_in_1_valid; // @[SpectrometerTest.scala 157:29]
  wire [31:0] out_mux_auto_stream_in_1_bits_data; // @[SpectrometerTest.scala 157:29]
  wire  out_mux_auto_stream_in_1_bits_last; // @[SpectrometerTest.scala 157:29]
  wire  out_mux_auto_stream_in_0_ready; // @[SpectrometerTest.scala 157:29]
  wire  out_mux_auto_stream_in_0_valid; // @[SpectrometerTest.scala 157:29]
  wire [31:0] out_mux_auto_stream_in_0_bits_data; // @[SpectrometerTest.scala 157:29]
  wire  out_mux_auto_stream_in_0_bits_last; // @[SpectrometerTest.scala 157:29]
  wire  out_mux_auto_stream_out_1_ready; // @[SpectrometerTest.scala 157:29]
  wire  out_mux_auto_stream_out_1_valid; // @[SpectrometerTest.scala 157:29]
  wire [31:0] out_mux_auto_stream_out_1_bits_data; // @[SpectrometerTest.scala 157:29]
  wire  out_mux_auto_stream_out_1_bits_last; // @[SpectrometerTest.scala 157:29]
  wire  out_mux_auto_stream_out_0_ready; // @[SpectrometerTest.scala 157:29]
  wire  out_mux_auto_stream_out_0_valid; // @[SpectrometerTest.scala 157:29]
  wire [31:0] out_mux_auto_stream_out_0_bits_data; // @[SpectrometerTest.scala 157:29]
  wire  out_mux_auto_stream_out_0_bits_last; // @[SpectrometerTest.scala 157:29]
  wire  out_queue_clock; // @[SpectrometerTest.scala 158:29]
  wire  out_queue_reset; // @[SpectrometerTest.scala 158:29]
  wire  out_queue_auto_out_out_ready; // @[SpectrometerTest.scala 158:29]
  wire  out_queue_auto_out_out_valid; // @[SpectrometerTest.scala 158:29]
  wire [31:0] out_queue_auto_out_out_bits_data; // @[SpectrometerTest.scala 158:29]
  wire  out_queue_auto_out_out_bits_last; // @[SpectrometerTest.scala 158:29]
  wire  out_queue_auto_in_in_ready; // @[SpectrometerTest.scala 158:29]
  wire  out_queue_auto_in_in_valid; // @[SpectrometerTest.scala 158:29]
  wire [31:0] out_queue_auto_in_in_bits_data; // @[SpectrometerTest.scala 158:29]
  wire  out_queue_auto_in_in_bits_last; // @[SpectrometerTest.scala 158:29]
  wire  widthAdapter_2_clock; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_2_reset; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_2_auto_in_ready; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_2_auto_in_valid; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire [31:0] widthAdapter_2_auto_in_bits_data; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_2_auto_in_bits_last; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_2_auto_out_ready; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_2_auto_out_valid; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire [7:0] widthAdapter_2_auto_out_bits_data; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_2_auto_out_bits_last; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  uTx_queue_clock; // @[SpectrometerTest.scala 162:29]
  wire  uTx_queue_reset; // @[SpectrometerTest.scala 162:29]
  wire  uTx_queue_auto_out_out_ready; // @[SpectrometerTest.scala 162:29]
  wire  uTx_queue_auto_out_out_valid; // @[SpectrometerTest.scala 162:29]
  wire [31:0] uTx_queue_auto_out_out_bits_data; // @[SpectrometerTest.scala 162:29]
  wire  uTx_queue_auto_out_out_bits_last; // @[SpectrometerTest.scala 162:29]
  wire  uTx_queue_auto_in_in_ready; // @[SpectrometerTest.scala 162:29]
  wire  uTx_queue_auto_in_in_valid; // @[SpectrometerTest.scala 162:29]
  wire [31:0] uTx_queue_auto_in_in_bits_data; // @[SpectrometerTest.scala 162:29]
  wire  uTx_queue_auto_in_in_bits_last; // @[SpectrometerTest.scala 162:29]
  wire  widthAdapter_3_clock; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_3_reset; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_3_auto_in_ready; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_3_auto_in_valid; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire [31:0] widthAdapter_3_auto_in_bits_data; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_3_auto_in_bits_last; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_3_auto_out_ready; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_3_auto_out_valid; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire [7:0] widthAdapter_3_auto_out_bits_data; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_3_auto_out_bits_last; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_4_clock; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_4_reset; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_4_auto_in_ready; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_4_auto_in_valid; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire [7:0] widthAdapter_4_auto_in_bits_data; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_4_auto_in_bits_last; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_4_auto_out_ready; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_4_auto_out_valid; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire [31:0] widthAdapter_4_auto_out_bits_data; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_4_auto_out_bits_last; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  uRx_split_clock; // @[SpectrometerTest.scala 165:29]
  wire  uRx_split_reset; // @[SpectrometerTest.scala 165:29]
  wire  uRx_split_auto_mem_in_aw_ready; // @[SpectrometerTest.scala 165:29]
  wire  uRx_split_auto_mem_in_aw_valid; // @[SpectrometerTest.scala 165:29]
  wire  uRx_split_auto_mem_in_aw_bits_id; // @[SpectrometerTest.scala 165:29]
  wire [29:0] uRx_split_auto_mem_in_aw_bits_addr; // @[SpectrometerTest.scala 165:29]
  wire  uRx_split_auto_mem_in_w_ready; // @[SpectrometerTest.scala 165:29]
  wire  uRx_split_auto_mem_in_w_valid; // @[SpectrometerTest.scala 165:29]
  wire [31:0] uRx_split_auto_mem_in_w_bits_data; // @[SpectrometerTest.scala 165:29]
  wire [3:0] uRx_split_auto_mem_in_w_bits_strb; // @[SpectrometerTest.scala 165:29]
  wire  uRx_split_auto_mem_in_b_ready; // @[SpectrometerTest.scala 165:29]
  wire  uRx_split_auto_mem_in_b_valid; // @[SpectrometerTest.scala 165:29]
  wire  uRx_split_auto_mem_in_b_bits_id; // @[SpectrometerTest.scala 165:29]
  wire  uRx_split_auto_mem_in_ar_ready; // @[SpectrometerTest.scala 165:29]
  wire  uRx_split_auto_mem_in_ar_valid; // @[SpectrometerTest.scala 165:29]
  wire  uRx_split_auto_mem_in_ar_bits_id; // @[SpectrometerTest.scala 165:29]
  wire [29:0] uRx_split_auto_mem_in_ar_bits_addr; // @[SpectrometerTest.scala 165:29]
  wire [2:0] uRx_split_auto_mem_in_ar_bits_size; // @[SpectrometerTest.scala 165:29]
  wire  uRx_split_auto_mem_in_r_ready; // @[SpectrometerTest.scala 165:29]
  wire  uRx_split_auto_mem_in_r_valid; // @[SpectrometerTest.scala 165:29]
  wire  uRx_split_auto_mem_in_r_bits_id; // @[SpectrometerTest.scala 165:29]
  wire [31:0] uRx_split_auto_mem_in_r_bits_data; // @[SpectrometerTest.scala 165:29]
  wire  uRx_split_auto_stream_in_ready; // @[SpectrometerTest.scala 165:29]
  wire  uRx_split_auto_stream_in_valid; // @[SpectrometerTest.scala 165:29]
  wire [31:0] uRx_split_auto_stream_in_bits_data; // @[SpectrometerTest.scala 165:29]
  wire  uRx_split_auto_stream_in_bits_last; // @[SpectrometerTest.scala 165:29]
  wire  uRx_split_auto_stream_out_4_ready; // @[SpectrometerTest.scala 165:29]
  wire  uRx_split_auto_stream_out_4_valid; // @[SpectrometerTest.scala 165:29]
  wire [31:0] uRx_split_auto_stream_out_4_bits_data; // @[SpectrometerTest.scala 165:29]
  wire  uRx_split_auto_stream_out_4_bits_last; // @[SpectrometerTest.scala 165:29]
  wire  uRx_split_auto_stream_out_3_ready; // @[SpectrometerTest.scala 165:29]
  wire  uRx_split_auto_stream_out_3_valid; // @[SpectrometerTest.scala 165:29]
  wire [31:0] uRx_split_auto_stream_out_3_bits_data; // @[SpectrometerTest.scala 165:29]
  wire  uRx_split_auto_stream_out_3_bits_last; // @[SpectrometerTest.scala 165:29]
  wire  uRx_split_auto_stream_out_2_ready; // @[SpectrometerTest.scala 165:29]
  wire  uRx_split_auto_stream_out_2_valid; // @[SpectrometerTest.scala 165:29]
  wire [31:0] uRx_split_auto_stream_out_2_bits_data; // @[SpectrometerTest.scala 165:29]
  wire  uRx_split_auto_stream_out_2_bits_last; // @[SpectrometerTest.scala 165:29]
  wire  uRx_split_auto_stream_out_1_ready; // @[SpectrometerTest.scala 165:29]
  wire  uRx_split_auto_stream_out_1_valid; // @[SpectrometerTest.scala 165:29]
  wire [31:0] uRx_split_auto_stream_out_1_bits_data; // @[SpectrometerTest.scala 165:29]
  wire  uRx_split_auto_stream_out_1_bits_last; // @[SpectrometerTest.scala 165:29]
  wire  uRx_split_auto_stream_out_0_ready; // @[SpectrometerTest.scala 165:29]
  wire  uRx_split_auto_stream_out_0_valid; // @[SpectrometerTest.scala 165:29]
  wire [31:0] uRx_split_auto_stream_out_0_bits_data; // @[SpectrometerTest.scala 165:29]
  wire  uRx_split_auto_stream_out_0_bits_last; // @[SpectrometerTest.scala 165:29]
  wire  uart_clock; // @[SpectrometerTest.scala 166:29]
  wire  uart_reset; // @[SpectrometerTest.scala 166:29]
  wire  uart_auto_mem_in_aw_ready; // @[SpectrometerTest.scala 166:29]
  wire  uart_auto_mem_in_aw_valid; // @[SpectrometerTest.scala 166:29]
  wire  uart_auto_mem_in_aw_bits_id; // @[SpectrometerTest.scala 166:29]
  wire [29:0] uart_auto_mem_in_aw_bits_addr; // @[SpectrometerTest.scala 166:29]
  wire  uart_auto_mem_in_w_ready; // @[SpectrometerTest.scala 166:29]
  wire  uart_auto_mem_in_w_valid; // @[SpectrometerTest.scala 166:29]
  wire [31:0] uart_auto_mem_in_w_bits_data; // @[SpectrometerTest.scala 166:29]
  wire [3:0] uart_auto_mem_in_w_bits_strb; // @[SpectrometerTest.scala 166:29]
  wire  uart_auto_mem_in_b_ready; // @[SpectrometerTest.scala 166:29]
  wire  uart_auto_mem_in_b_valid; // @[SpectrometerTest.scala 166:29]
  wire  uart_auto_mem_in_b_bits_id; // @[SpectrometerTest.scala 166:29]
  wire  uart_auto_mem_in_ar_ready; // @[SpectrometerTest.scala 166:29]
  wire  uart_auto_mem_in_ar_valid; // @[SpectrometerTest.scala 166:29]
  wire  uart_auto_mem_in_ar_bits_id; // @[SpectrometerTest.scala 166:29]
  wire [29:0] uart_auto_mem_in_ar_bits_addr; // @[SpectrometerTest.scala 166:29]
  wire [2:0] uart_auto_mem_in_ar_bits_size; // @[SpectrometerTest.scala 166:29]
  wire  uart_auto_mem_in_r_ready; // @[SpectrometerTest.scala 166:29]
  wire  uart_auto_mem_in_r_valid; // @[SpectrometerTest.scala 166:29]
  wire  uart_auto_mem_in_r_bits_id; // @[SpectrometerTest.scala 166:29]
  wire [31:0] uart_auto_mem_in_r_bits_data; // @[SpectrometerTest.scala 166:29]
  wire  uart_auto_in_in_ready; // @[SpectrometerTest.scala 166:29]
  wire  uart_auto_in_in_valid; // @[SpectrometerTest.scala 166:29]
  wire [7:0] uart_auto_in_in_bits_data; // @[SpectrometerTest.scala 166:29]
  wire  uart_auto_out_out_ready; // @[SpectrometerTest.scala 166:29]
  wire  uart_auto_out_out_valid; // @[SpectrometerTest.scala 166:29]
  wire [7:0] uart_auto_out_out_bits_data; // @[SpectrometerTest.scala 166:29]
  wire  uart_int_0; // @[SpectrometerTest.scala 166:29]
  wire  uart_io_txd; // @[SpectrometerTest.scala 166:29]
  wire  uart_io_rxd; // @[SpectrometerTest.scala 166:29]
  wire  bus_clock; // @[SpectrometerTest.scala 180:23]
  wire  bus_reset; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_in_aw_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_in_aw_valid; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_in_aw_bits_id; // @[SpectrometerTest.scala 180:23]
  wire [29:0] bus_auto_in_aw_bits_addr; // @[SpectrometerTest.scala 180:23]
  wire [2:0] bus_auto_in_aw_bits_size; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_in_w_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_in_w_valid; // @[SpectrometerTest.scala 180:23]
  wire [31:0] bus_auto_in_w_bits_data; // @[SpectrometerTest.scala 180:23]
  wire [3:0] bus_auto_in_w_bits_strb; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_in_w_bits_last; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_in_b_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_in_b_valid; // @[SpectrometerTest.scala 180:23]
  wire [1:0] bus_auto_in_b_bits_resp; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_in_ar_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_in_ar_valid; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_in_ar_bits_id; // @[SpectrometerTest.scala 180:23]
  wire [29:0] bus_auto_in_ar_bits_addr; // @[SpectrometerTest.scala 180:23]
  wire [2:0] bus_auto_in_ar_bits_size; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_in_r_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_in_r_valid; // @[SpectrometerTest.scala 180:23]
  wire [31:0] bus_auto_in_r_bits_data; // @[SpectrometerTest.scala 180:23]
  wire [1:0] bus_auto_in_r_bits_resp; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_in_r_bits_last; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_20_aw_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_20_aw_valid; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_20_aw_bits_id; // @[SpectrometerTest.scala 180:23]
  wire [29:0] bus_auto_out_20_aw_bits_addr; // @[SpectrometerTest.scala 180:23]
  wire [2:0] bus_auto_out_20_aw_bits_size; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_20_w_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_20_w_valid; // @[SpectrometerTest.scala 180:23]
  wire [31:0] bus_auto_out_20_w_bits_data; // @[SpectrometerTest.scala 180:23]
  wire [3:0] bus_auto_out_20_w_bits_strb; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_20_w_bits_last; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_20_b_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_20_b_valid; // @[SpectrometerTest.scala 180:23]
  wire [1:0] bus_auto_out_20_b_bits_resp; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_20_ar_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_20_ar_valid; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_20_ar_bits_id; // @[SpectrometerTest.scala 180:23]
  wire [29:0] bus_auto_out_20_ar_bits_addr; // @[SpectrometerTest.scala 180:23]
  wire [2:0] bus_auto_out_20_ar_bits_size; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_20_r_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_20_r_valid; // @[SpectrometerTest.scala 180:23]
  wire [31:0] bus_auto_out_20_r_bits_data; // @[SpectrometerTest.scala 180:23]
  wire [1:0] bus_auto_out_20_r_bits_resp; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_20_r_bits_last; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_19_aw_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_19_aw_valid; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_19_aw_bits_id; // @[SpectrometerTest.scala 180:23]
  wire [29:0] bus_auto_out_19_aw_bits_addr; // @[SpectrometerTest.scala 180:23]
  wire [2:0] bus_auto_out_19_aw_bits_size; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_19_w_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_19_w_valid; // @[SpectrometerTest.scala 180:23]
  wire [31:0] bus_auto_out_19_w_bits_data; // @[SpectrometerTest.scala 180:23]
  wire [3:0] bus_auto_out_19_w_bits_strb; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_19_w_bits_last; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_19_b_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_19_b_valid; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_19_b_bits_id; // @[SpectrometerTest.scala 180:23]
  wire [1:0] bus_auto_out_19_b_bits_resp; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_19_ar_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_19_ar_valid; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_19_ar_bits_id; // @[SpectrometerTest.scala 180:23]
  wire [29:0] bus_auto_out_19_ar_bits_addr; // @[SpectrometerTest.scala 180:23]
  wire [2:0] bus_auto_out_19_ar_bits_size; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_19_r_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_19_r_valid; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_19_r_bits_id; // @[SpectrometerTest.scala 180:23]
  wire [31:0] bus_auto_out_19_r_bits_data; // @[SpectrometerTest.scala 180:23]
  wire [1:0] bus_auto_out_19_r_bits_resp; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_19_r_bits_last; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_18_aw_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_18_aw_valid; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_18_aw_bits_id; // @[SpectrometerTest.scala 180:23]
  wire [29:0] bus_auto_out_18_aw_bits_addr; // @[SpectrometerTest.scala 180:23]
  wire [2:0] bus_auto_out_18_aw_bits_size; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_18_w_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_18_w_valid; // @[SpectrometerTest.scala 180:23]
  wire [31:0] bus_auto_out_18_w_bits_data; // @[SpectrometerTest.scala 180:23]
  wire [3:0] bus_auto_out_18_w_bits_strb; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_18_w_bits_last; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_18_b_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_18_b_valid; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_18_b_bits_id; // @[SpectrometerTest.scala 180:23]
  wire [1:0] bus_auto_out_18_b_bits_resp; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_18_ar_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_18_ar_valid; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_18_ar_bits_id; // @[SpectrometerTest.scala 180:23]
  wire [29:0] bus_auto_out_18_ar_bits_addr; // @[SpectrometerTest.scala 180:23]
  wire [2:0] bus_auto_out_18_ar_bits_size; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_18_r_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_18_r_valid; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_18_r_bits_id; // @[SpectrometerTest.scala 180:23]
  wire [31:0] bus_auto_out_18_r_bits_data; // @[SpectrometerTest.scala 180:23]
  wire [1:0] bus_auto_out_18_r_bits_resp; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_18_r_bits_last; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_17_aw_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_17_aw_valid; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_17_aw_bits_id; // @[SpectrometerTest.scala 180:23]
  wire [29:0] bus_auto_out_17_aw_bits_addr; // @[SpectrometerTest.scala 180:23]
  wire [2:0] bus_auto_out_17_aw_bits_size; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_17_w_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_17_w_valid; // @[SpectrometerTest.scala 180:23]
  wire [31:0] bus_auto_out_17_w_bits_data; // @[SpectrometerTest.scala 180:23]
  wire [3:0] bus_auto_out_17_w_bits_strb; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_17_w_bits_last; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_17_b_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_17_b_valid; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_17_b_bits_id; // @[SpectrometerTest.scala 180:23]
  wire [1:0] bus_auto_out_17_b_bits_resp; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_17_ar_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_17_ar_valid; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_17_ar_bits_id; // @[SpectrometerTest.scala 180:23]
  wire [29:0] bus_auto_out_17_ar_bits_addr; // @[SpectrometerTest.scala 180:23]
  wire [2:0] bus_auto_out_17_ar_bits_size; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_17_r_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_17_r_valid; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_17_r_bits_id; // @[SpectrometerTest.scala 180:23]
  wire [31:0] bus_auto_out_17_r_bits_data; // @[SpectrometerTest.scala 180:23]
  wire [1:0] bus_auto_out_17_r_bits_resp; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_17_r_bits_last; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_16_aw_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_16_aw_valid; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_16_aw_bits_id; // @[SpectrometerTest.scala 180:23]
  wire [29:0] bus_auto_out_16_aw_bits_addr; // @[SpectrometerTest.scala 180:23]
  wire [2:0] bus_auto_out_16_aw_bits_size; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_16_w_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_16_w_valid; // @[SpectrometerTest.scala 180:23]
  wire [31:0] bus_auto_out_16_w_bits_data; // @[SpectrometerTest.scala 180:23]
  wire [3:0] bus_auto_out_16_w_bits_strb; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_16_w_bits_last; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_16_b_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_16_b_valid; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_16_b_bits_id; // @[SpectrometerTest.scala 180:23]
  wire [1:0] bus_auto_out_16_b_bits_resp; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_16_ar_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_16_ar_valid; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_16_ar_bits_id; // @[SpectrometerTest.scala 180:23]
  wire [29:0] bus_auto_out_16_ar_bits_addr; // @[SpectrometerTest.scala 180:23]
  wire [2:0] bus_auto_out_16_ar_bits_size; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_16_r_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_16_r_valid; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_16_r_bits_id; // @[SpectrometerTest.scala 180:23]
  wire [31:0] bus_auto_out_16_r_bits_data; // @[SpectrometerTest.scala 180:23]
  wire [1:0] bus_auto_out_16_r_bits_resp; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_16_r_bits_last; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_15_aw_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_15_aw_valid; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_15_aw_bits_id; // @[SpectrometerTest.scala 180:23]
  wire [29:0] bus_auto_out_15_aw_bits_addr; // @[SpectrometerTest.scala 180:23]
  wire [2:0] bus_auto_out_15_aw_bits_size; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_15_w_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_15_w_valid; // @[SpectrometerTest.scala 180:23]
  wire [31:0] bus_auto_out_15_w_bits_data; // @[SpectrometerTest.scala 180:23]
  wire [3:0] bus_auto_out_15_w_bits_strb; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_15_w_bits_last; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_15_b_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_15_b_valid; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_15_b_bits_id; // @[SpectrometerTest.scala 180:23]
  wire [1:0] bus_auto_out_15_b_bits_resp; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_15_ar_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_15_ar_valid; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_15_ar_bits_id; // @[SpectrometerTest.scala 180:23]
  wire [29:0] bus_auto_out_15_ar_bits_addr; // @[SpectrometerTest.scala 180:23]
  wire [2:0] bus_auto_out_15_ar_bits_size; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_15_r_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_15_r_valid; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_15_r_bits_id; // @[SpectrometerTest.scala 180:23]
  wire [31:0] bus_auto_out_15_r_bits_data; // @[SpectrometerTest.scala 180:23]
  wire [1:0] bus_auto_out_15_r_bits_resp; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_15_r_bits_last; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_14_aw_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_14_aw_valid; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_14_aw_bits_id; // @[SpectrometerTest.scala 180:23]
  wire [29:0] bus_auto_out_14_aw_bits_addr; // @[SpectrometerTest.scala 180:23]
  wire [2:0] bus_auto_out_14_aw_bits_size; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_14_w_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_14_w_valid; // @[SpectrometerTest.scala 180:23]
  wire [31:0] bus_auto_out_14_w_bits_data; // @[SpectrometerTest.scala 180:23]
  wire [3:0] bus_auto_out_14_w_bits_strb; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_14_w_bits_last; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_14_b_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_14_b_valid; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_14_b_bits_id; // @[SpectrometerTest.scala 180:23]
  wire [1:0] bus_auto_out_14_b_bits_resp; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_14_ar_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_14_ar_valid; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_14_ar_bits_id; // @[SpectrometerTest.scala 180:23]
  wire [29:0] bus_auto_out_14_ar_bits_addr; // @[SpectrometerTest.scala 180:23]
  wire [2:0] bus_auto_out_14_ar_bits_size; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_14_r_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_14_r_valid; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_14_r_bits_id; // @[SpectrometerTest.scala 180:23]
  wire [31:0] bus_auto_out_14_r_bits_data; // @[SpectrometerTest.scala 180:23]
  wire [1:0] bus_auto_out_14_r_bits_resp; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_14_r_bits_last; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_13_aw_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_13_aw_valid; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_13_aw_bits_id; // @[SpectrometerTest.scala 180:23]
  wire [29:0] bus_auto_out_13_aw_bits_addr; // @[SpectrometerTest.scala 180:23]
  wire [2:0] bus_auto_out_13_aw_bits_size; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_13_w_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_13_w_valid; // @[SpectrometerTest.scala 180:23]
  wire [31:0] bus_auto_out_13_w_bits_data; // @[SpectrometerTest.scala 180:23]
  wire [3:0] bus_auto_out_13_w_bits_strb; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_13_w_bits_last; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_13_b_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_13_b_valid; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_13_b_bits_id; // @[SpectrometerTest.scala 180:23]
  wire [1:0] bus_auto_out_13_b_bits_resp; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_13_ar_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_13_ar_valid; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_13_ar_bits_id; // @[SpectrometerTest.scala 180:23]
  wire [29:0] bus_auto_out_13_ar_bits_addr; // @[SpectrometerTest.scala 180:23]
  wire [2:0] bus_auto_out_13_ar_bits_size; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_13_r_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_13_r_valid; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_13_r_bits_id; // @[SpectrometerTest.scala 180:23]
  wire [31:0] bus_auto_out_13_r_bits_data; // @[SpectrometerTest.scala 180:23]
  wire [1:0] bus_auto_out_13_r_bits_resp; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_13_r_bits_last; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_12_aw_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_12_aw_valid; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_12_aw_bits_id; // @[SpectrometerTest.scala 180:23]
  wire [29:0] bus_auto_out_12_aw_bits_addr; // @[SpectrometerTest.scala 180:23]
  wire [2:0] bus_auto_out_12_aw_bits_size; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_12_w_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_12_w_valid; // @[SpectrometerTest.scala 180:23]
  wire [31:0] bus_auto_out_12_w_bits_data; // @[SpectrometerTest.scala 180:23]
  wire [3:0] bus_auto_out_12_w_bits_strb; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_12_w_bits_last; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_12_b_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_12_b_valid; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_12_b_bits_id; // @[SpectrometerTest.scala 180:23]
  wire [1:0] bus_auto_out_12_b_bits_resp; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_12_ar_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_12_ar_valid; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_12_ar_bits_id; // @[SpectrometerTest.scala 180:23]
  wire [29:0] bus_auto_out_12_ar_bits_addr; // @[SpectrometerTest.scala 180:23]
  wire [2:0] bus_auto_out_12_ar_bits_size; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_12_r_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_12_r_valid; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_12_r_bits_id; // @[SpectrometerTest.scala 180:23]
  wire [31:0] bus_auto_out_12_r_bits_data; // @[SpectrometerTest.scala 180:23]
  wire [1:0] bus_auto_out_12_r_bits_resp; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_12_r_bits_last; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_11_aw_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_11_aw_valid; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_11_aw_bits_id; // @[SpectrometerTest.scala 180:23]
  wire [29:0] bus_auto_out_11_aw_bits_addr; // @[SpectrometerTest.scala 180:23]
  wire [2:0] bus_auto_out_11_aw_bits_size; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_11_w_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_11_w_valid; // @[SpectrometerTest.scala 180:23]
  wire [31:0] bus_auto_out_11_w_bits_data; // @[SpectrometerTest.scala 180:23]
  wire [3:0] bus_auto_out_11_w_bits_strb; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_11_w_bits_last; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_11_b_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_11_b_valid; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_11_b_bits_id; // @[SpectrometerTest.scala 180:23]
  wire [1:0] bus_auto_out_11_b_bits_resp; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_11_ar_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_11_ar_valid; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_11_ar_bits_id; // @[SpectrometerTest.scala 180:23]
  wire [29:0] bus_auto_out_11_ar_bits_addr; // @[SpectrometerTest.scala 180:23]
  wire [2:0] bus_auto_out_11_ar_bits_size; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_11_r_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_11_r_valid; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_11_r_bits_id; // @[SpectrometerTest.scala 180:23]
  wire [31:0] bus_auto_out_11_r_bits_data; // @[SpectrometerTest.scala 180:23]
  wire [1:0] bus_auto_out_11_r_bits_resp; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_11_r_bits_last; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_10_aw_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_10_aw_valid; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_10_aw_bits_id; // @[SpectrometerTest.scala 180:23]
  wire [29:0] bus_auto_out_10_aw_bits_addr; // @[SpectrometerTest.scala 180:23]
  wire [2:0] bus_auto_out_10_aw_bits_size; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_10_w_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_10_w_valid; // @[SpectrometerTest.scala 180:23]
  wire [31:0] bus_auto_out_10_w_bits_data; // @[SpectrometerTest.scala 180:23]
  wire [3:0] bus_auto_out_10_w_bits_strb; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_10_w_bits_last; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_10_b_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_10_b_valid; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_10_b_bits_id; // @[SpectrometerTest.scala 180:23]
  wire [1:0] bus_auto_out_10_b_bits_resp; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_10_ar_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_10_ar_valid; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_10_ar_bits_id; // @[SpectrometerTest.scala 180:23]
  wire [29:0] bus_auto_out_10_ar_bits_addr; // @[SpectrometerTest.scala 180:23]
  wire [2:0] bus_auto_out_10_ar_bits_size; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_10_r_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_10_r_valid; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_10_r_bits_id; // @[SpectrometerTest.scala 180:23]
  wire [31:0] bus_auto_out_10_r_bits_data; // @[SpectrometerTest.scala 180:23]
  wire [1:0] bus_auto_out_10_r_bits_resp; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_10_r_bits_last; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_9_aw_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_9_aw_valid; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_9_aw_bits_id; // @[SpectrometerTest.scala 180:23]
  wire [29:0] bus_auto_out_9_aw_bits_addr; // @[SpectrometerTest.scala 180:23]
  wire [2:0] bus_auto_out_9_aw_bits_size; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_9_w_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_9_w_valid; // @[SpectrometerTest.scala 180:23]
  wire [31:0] bus_auto_out_9_w_bits_data; // @[SpectrometerTest.scala 180:23]
  wire [3:0] bus_auto_out_9_w_bits_strb; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_9_w_bits_last; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_9_b_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_9_b_valid; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_9_b_bits_id; // @[SpectrometerTest.scala 180:23]
  wire [1:0] bus_auto_out_9_b_bits_resp; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_9_ar_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_9_ar_valid; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_9_ar_bits_id; // @[SpectrometerTest.scala 180:23]
  wire [29:0] bus_auto_out_9_ar_bits_addr; // @[SpectrometerTest.scala 180:23]
  wire [2:0] bus_auto_out_9_ar_bits_size; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_9_r_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_9_r_valid; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_9_r_bits_id; // @[SpectrometerTest.scala 180:23]
  wire [31:0] bus_auto_out_9_r_bits_data; // @[SpectrometerTest.scala 180:23]
  wire [1:0] bus_auto_out_9_r_bits_resp; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_9_r_bits_last; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_8_aw_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_8_aw_valid; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_8_aw_bits_id; // @[SpectrometerTest.scala 180:23]
  wire [29:0] bus_auto_out_8_aw_bits_addr; // @[SpectrometerTest.scala 180:23]
  wire [2:0] bus_auto_out_8_aw_bits_size; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_8_w_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_8_w_valid; // @[SpectrometerTest.scala 180:23]
  wire [31:0] bus_auto_out_8_w_bits_data; // @[SpectrometerTest.scala 180:23]
  wire [3:0] bus_auto_out_8_w_bits_strb; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_8_w_bits_last; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_8_b_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_8_b_valid; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_8_b_bits_id; // @[SpectrometerTest.scala 180:23]
  wire [1:0] bus_auto_out_8_b_bits_resp; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_8_ar_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_8_ar_valid; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_8_ar_bits_id; // @[SpectrometerTest.scala 180:23]
  wire [29:0] bus_auto_out_8_ar_bits_addr; // @[SpectrometerTest.scala 180:23]
  wire [2:0] bus_auto_out_8_ar_bits_size; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_8_r_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_8_r_valid; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_8_r_bits_id; // @[SpectrometerTest.scala 180:23]
  wire [31:0] bus_auto_out_8_r_bits_data; // @[SpectrometerTest.scala 180:23]
  wire [1:0] bus_auto_out_8_r_bits_resp; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_8_r_bits_last; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_7_aw_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_7_aw_valid; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_7_aw_bits_id; // @[SpectrometerTest.scala 180:23]
  wire [29:0] bus_auto_out_7_aw_bits_addr; // @[SpectrometerTest.scala 180:23]
  wire [2:0] bus_auto_out_7_aw_bits_size; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_7_w_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_7_w_valid; // @[SpectrometerTest.scala 180:23]
  wire [31:0] bus_auto_out_7_w_bits_data; // @[SpectrometerTest.scala 180:23]
  wire [3:0] bus_auto_out_7_w_bits_strb; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_7_w_bits_last; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_7_b_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_7_b_valid; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_7_b_bits_id; // @[SpectrometerTest.scala 180:23]
  wire [1:0] bus_auto_out_7_b_bits_resp; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_7_ar_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_7_ar_valid; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_7_ar_bits_id; // @[SpectrometerTest.scala 180:23]
  wire [29:0] bus_auto_out_7_ar_bits_addr; // @[SpectrometerTest.scala 180:23]
  wire [2:0] bus_auto_out_7_ar_bits_size; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_7_r_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_7_r_valid; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_7_r_bits_id; // @[SpectrometerTest.scala 180:23]
  wire [31:0] bus_auto_out_7_r_bits_data; // @[SpectrometerTest.scala 180:23]
  wire [1:0] bus_auto_out_7_r_bits_resp; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_7_r_bits_last; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_6_aw_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_6_aw_valid; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_6_aw_bits_id; // @[SpectrometerTest.scala 180:23]
  wire [29:0] bus_auto_out_6_aw_bits_addr; // @[SpectrometerTest.scala 180:23]
  wire [2:0] bus_auto_out_6_aw_bits_size; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_6_w_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_6_w_valid; // @[SpectrometerTest.scala 180:23]
  wire [31:0] bus_auto_out_6_w_bits_data; // @[SpectrometerTest.scala 180:23]
  wire [3:0] bus_auto_out_6_w_bits_strb; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_6_w_bits_last; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_6_b_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_6_b_valid; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_6_b_bits_id; // @[SpectrometerTest.scala 180:23]
  wire [1:0] bus_auto_out_6_b_bits_resp; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_6_ar_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_6_ar_valid; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_6_ar_bits_id; // @[SpectrometerTest.scala 180:23]
  wire [29:0] bus_auto_out_6_ar_bits_addr; // @[SpectrometerTest.scala 180:23]
  wire [2:0] bus_auto_out_6_ar_bits_size; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_6_r_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_6_r_valid; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_6_r_bits_id; // @[SpectrometerTest.scala 180:23]
  wire [31:0] bus_auto_out_6_r_bits_data; // @[SpectrometerTest.scala 180:23]
  wire [1:0] bus_auto_out_6_r_bits_resp; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_6_r_bits_last; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_5_aw_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_5_aw_valid; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_5_aw_bits_id; // @[SpectrometerTest.scala 180:23]
  wire [29:0] bus_auto_out_5_aw_bits_addr; // @[SpectrometerTest.scala 180:23]
  wire [2:0] bus_auto_out_5_aw_bits_size; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_5_w_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_5_w_valid; // @[SpectrometerTest.scala 180:23]
  wire [31:0] bus_auto_out_5_w_bits_data; // @[SpectrometerTest.scala 180:23]
  wire [3:0] bus_auto_out_5_w_bits_strb; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_5_w_bits_last; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_5_b_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_5_b_valid; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_5_b_bits_id; // @[SpectrometerTest.scala 180:23]
  wire [1:0] bus_auto_out_5_b_bits_resp; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_5_ar_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_5_ar_valid; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_5_ar_bits_id; // @[SpectrometerTest.scala 180:23]
  wire [29:0] bus_auto_out_5_ar_bits_addr; // @[SpectrometerTest.scala 180:23]
  wire [2:0] bus_auto_out_5_ar_bits_size; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_5_r_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_5_r_valid; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_5_r_bits_id; // @[SpectrometerTest.scala 180:23]
  wire [31:0] bus_auto_out_5_r_bits_data; // @[SpectrometerTest.scala 180:23]
  wire [1:0] bus_auto_out_5_r_bits_resp; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_5_r_bits_last; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_4_aw_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_4_aw_valid; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_4_aw_bits_id; // @[SpectrometerTest.scala 180:23]
  wire [29:0] bus_auto_out_4_aw_bits_addr; // @[SpectrometerTest.scala 180:23]
  wire [2:0] bus_auto_out_4_aw_bits_size; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_4_w_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_4_w_valid; // @[SpectrometerTest.scala 180:23]
  wire [31:0] bus_auto_out_4_w_bits_data; // @[SpectrometerTest.scala 180:23]
  wire [3:0] bus_auto_out_4_w_bits_strb; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_4_w_bits_last; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_4_b_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_4_b_valid; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_4_b_bits_id; // @[SpectrometerTest.scala 180:23]
  wire [1:0] bus_auto_out_4_b_bits_resp; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_4_ar_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_4_ar_valid; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_4_ar_bits_id; // @[SpectrometerTest.scala 180:23]
  wire [29:0] bus_auto_out_4_ar_bits_addr; // @[SpectrometerTest.scala 180:23]
  wire [2:0] bus_auto_out_4_ar_bits_size; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_4_r_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_4_r_valid; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_4_r_bits_id; // @[SpectrometerTest.scala 180:23]
  wire [31:0] bus_auto_out_4_r_bits_data; // @[SpectrometerTest.scala 180:23]
  wire [1:0] bus_auto_out_4_r_bits_resp; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_4_r_bits_last; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_3_aw_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_3_aw_valid; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_3_aw_bits_id; // @[SpectrometerTest.scala 180:23]
  wire [29:0] bus_auto_out_3_aw_bits_addr; // @[SpectrometerTest.scala 180:23]
  wire [2:0] bus_auto_out_3_aw_bits_size; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_3_w_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_3_w_valid; // @[SpectrometerTest.scala 180:23]
  wire [31:0] bus_auto_out_3_w_bits_data; // @[SpectrometerTest.scala 180:23]
  wire [3:0] bus_auto_out_3_w_bits_strb; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_3_w_bits_last; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_3_b_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_3_b_valid; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_3_b_bits_id; // @[SpectrometerTest.scala 180:23]
  wire [1:0] bus_auto_out_3_b_bits_resp; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_3_ar_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_3_ar_valid; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_3_ar_bits_id; // @[SpectrometerTest.scala 180:23]
  wire [29:0] bus_auto_out_3_ar_bits_addr; // @[SpectrometerTest.scala 180:23]
  wire [2:0] bus_auto_out_3_ar_bits_size; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_3_r_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_3_r_valid; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_3_r_bits_id; // @[SpectrometerTest.scala 180:23]
  wire [31:0] bus_auto_out_3_r_bits_data; // @[SpectrometerTest.scala 180:23]
  wire [1:0] bus_auto_out_3_r_bits_resp; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_3_r_bits_last; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_2_aw_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_2_aw_valid; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_2_aw_bits_id; // @[SpectrometerTest.scala 180:23]
  wire [29:0] bus_auto_out_2_aw_bits_addr; // @[SpectrometerTest.scala 180:23]
  wire [2:0] bus_auto_out_2_aw_bits_size; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_2_w_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_2_w_valid; // @[SpectrometerTest.scala 180:23]
  wire [31:0] bus_auto_out_2_w_bits_data; // @[SpectrometerTest.scala 180:23]
  wire [3:0] bus_auto_out_2_w_bits_strb; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_2_w_bits_last; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_2_b_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_2_b_valid; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_2_b_bits_id; // @[SpectrometerTest.scala 180:23]
  wire [1:0] bus_auto_out_2_b_bits_resp; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_2_ar_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_2_ar_valid; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_2_ar_bits_id; // @[SpectrometerTest.scala 180:23]
  wire [29:0] bus_auto_out_2_ar_bits_addr; // @[SpectrometerTest.scala 180:23]
  wire [2:0] bus_auto_out_2_ar_bits_size; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_2_r_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_2_r_valid; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_2_r_bits_id; // @[SpectrometerTest.scala 180:23]
  wire [31:0] bus_auto_out_2_r_bits_data; // @[SpectrometerTest.scala 180:23]
  wire [1:0] bus_auto_out_2_r_bits_resp; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_2_r_bits_last; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_1_aw_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_1_aw_valid; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_1_aw_bits_id; // @[SpectrometerTest.scala 180:23]
  wire [29:0] bus_auto_out_1_aw_bits_addr; // @[SpectrometerTest.scala 180:23]
  wire [2:0] bus_auto_out_1_aw_bits_size; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_1_w_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_1_w_valid; // @[SpectrometerTest.scala 180:23]
  wire [31:0] bus_auto_out_1_w_bits_data; // @[SpectrometerTest.scala 180:23]
  wire [3:0] bus_auto_out_1_w_bits_strb; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_1_w_bits_last; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_1_b_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_1_b_valid; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_1_b_bits_id; // @[SpectrometerTest.scala 180:23]
  wire [1:0] bus_auto_out_1_b_bits_resp; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_1_ar_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_1_ar_valid; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_1_ar_bits_id; // @[SpectrometerTest.scala 180:23]
  wire [29:0] bus_auto_out_1_ar_bits_addr; // @[SpectrometerTest.scala 180:23]
  wire [2:0] bus_auto_out_1_ar_bits_size; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_1_r_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_1_r_valid; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_1_r_bits_id; // @[SpectrometerTest.scala 180:23]
  wire [31:0] bus_auto_out_1_r_bits_data; // @[SpectrometerTest.scala 180:23]
  wire [1:0] bus_auto_out_1_r_bits_resp; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_1_r_bits_last; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_0_aw_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_0_aw_valid; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_0_aw_bits_id; // @[SpectrometerTest.scala 180:23]
  wire [29:0] bus_auto_out_0_aw_bits_addr; // @[SpectrometerTest.scala 180:23]
  wire [2:0] bus_auto_out_0_aw_bits_size; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_0_w_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_0_w_valid; // @[SpectrometerTest.scala 180:23]
  wire [31:0] bus_auto_out_0_w_bits_data; // @[SpectrometerTest.scala 180:23]
  wire [3:0] bus_auto_out_0_w_bits_strb; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_0_w_bits_last; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_0_b_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_0_b_valid; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_0_b_bits_id; // @[SpectrometerTest.scala 180:23]
  wire [1:0] bus_auto_out_0_b_bits_resp; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_0_ar_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_0_ar_valid; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_0_ar_bits_id; // @[SpectrometerTest.scala 180:23]
  wire [29:0] bus_auto_out_0_ar_bits_addr; // @[SpectrometerTest.scala 180:23]
  wire [2:0] bus_auto_out_0_ar_bits_size; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_0_r_ready; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_0_r_valid; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_0_r_bits_id; // @[SpectrometerTest.scala 180:23]
  wire [31:0] bus_auto_out_0_r_bits_data; // @[SpectrometerTest.scala 180:23]
  wire [1:0] bus_auto_out_0_r_bits_resp; // @[SpectrometerTest.scala 180:23]
  wire  bus_auto_out_0_r_bits_last; // @[SpectrometerTest.scala 180:23]
  wire  axi4buf_clock; // @[Buffer.scala 58:29]
  wire  axi4buf_reset; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_in_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_in_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_in_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_auto_in_aw_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_auto_in_aw_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_in_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_in_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_auto_in_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_auto_in_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_in_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_in_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_in_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_in_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_auto_in_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_in_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_in_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_in_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_auto_in_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_auto_in_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_in_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_in_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_in_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_auto_in_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_auto_in_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_in_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_out_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_out_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_out_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_auto_out_aw_bits_addr; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_out_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_out_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_auto_out_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_auto_out_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_out_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_out_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_out_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_out_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_auto_out_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_out_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_out_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_out_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_auto_out_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_auto_out_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_out_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_out_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_out_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_auto_out_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_auto_out_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_out_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_1_clock; // @[Buffer.scala 58:29]
  wire  axi4buf_1_reset; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_in_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_in_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_in_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_1_auto_in_aw_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_1_auto_in_aw_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_in_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_in_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_1_auto_in_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_1_auto_in_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_in_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_in_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_in_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_in_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_1_auto_in_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_in_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_in_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_in_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_1_auto_in_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_1_auto_in_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_in_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_in_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_in_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_1_auto_in_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_1_auto_in_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_in_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_out_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_out_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_out_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_1_auto_out_aw_bits_addr; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_out_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_out_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_1_auto_out_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_1_auto_out_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_out_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_out_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_out_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_out_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_1_auto_out_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_out_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_out_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_out_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_1_auto_out_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_1_auto_out_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_out_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_out_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_out_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_1_auto_out_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_1_auto_out_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_out_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_2_clock; // @[Buffer.scala 58:29]
  wire  axi4buf_2_reset; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_in_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_in_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_in_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_2_auto_in_aw_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_2_auto_in_aw_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_in_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_in_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_2_auto_in_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_2_auto_in_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_in_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_in_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_in_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_in_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_2_auto_in_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_in_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_in_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_in_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_2_auto_in_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_2_auto_in_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_in_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_in_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_in_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_2_auto_in_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_2_auto_in_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_in_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_out_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_out_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_out_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_2_auto_out_aw_bits_addr; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_out_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_out_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_2_auto_out_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_2_auto_out_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_out_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_out_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_out_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_out_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_2_auto_out_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_out_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_out_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_out_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_2_auto_out_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_2_auto_out_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_out_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_out_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_out_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_2_auto_out_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_2_auto_out_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_out_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_3_clock; // @[Buffer.scala 58:29]
  wire  axi4buf_3_reset; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_in_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_in_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_in_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_3_auto_in_aw_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_3_auto_in_aw_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_in_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_in_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_3_auto_in_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_3_auto_in_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_in_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_in_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_in_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_in_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_3_auto_in_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_in_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_in_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_in_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_3_auto_in_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_3_auto_in_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_in_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_in_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_in_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_3_auto_in_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_3_auto_in_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_in_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_out_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_out_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_out_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_3_auto_out_aw_bits_addr; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_out_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_out_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_3_auto_out_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_3_auto_out_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_out_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_out_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_out_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_out_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_3_auto_out_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_out_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_out_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_out_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_3_auto_out_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_3_auto_out_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_out_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_out_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_out_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_3_auto_out_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_3_auto_out_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_out_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_4_clock; // @[Buffer.scala 58:29]
  wire  axi4buf_4_reset; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_in_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_in_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_in_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_4_auto_in_aw_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_4_auto_in_aw_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_in_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_in_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_4_auto_in_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_4_auto_in_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_in_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_in_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_in_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_in_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_4_auto_in_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_in_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_in_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_in_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_4_auto_in_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_4_auto_in_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_in_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_in_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_in_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_4_auto_in_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_4_auto_in_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_in_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_out_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_out_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_out_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_4_auto_out_aw_bits_addr; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_out_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_out_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_4_auto_out_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_4_auto_out_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_out_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_out_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_out_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_out_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_4_auto_out_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_out_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_out_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_out_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_4_auto_out_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_4_auto_out_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_out_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_out_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_out_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_4_auto_out_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_4_auto_out_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_out_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_5_clock; // @[Buffer.scala 58:29]
  wire  axi4buf_5_reset; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_in_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_in_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_in_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_5_auto_in_aw_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_5_auto_in_aw_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_in_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_in_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_5_auto_in_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_5_auto_in_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_in_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_in_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_in_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_in_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_5_auto_in_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_in_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_in_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_in_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_5_auto_in_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_5_auto_in_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_in_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_in_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_in_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_5_auto_in_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_5_auto_in_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_in_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_out_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_out_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_out_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_5_auto_out_aw_bits_addr; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_out_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_out_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_5_auto_out_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_5_auto_out_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_out_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_out_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_out_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_out_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_5_auto_out_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_out_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_out_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_out_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_5_auto_out_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_5_auto_out_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_out_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_out_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_out_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_5_auto_out_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_5_auto_out_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_out_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_6_clock; // @[Buffer.scala 58:29]
  wire  axi4buf_6_reset; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_in_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_in_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_in_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_6_auto_in_aw_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_6_auto_in_aw_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_in_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_in_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_6_auto_in_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_6_auto_in_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_in_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_in_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_in_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_in_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_6_auto_in_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_in_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_in_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_in_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_6_auto_in_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_6_auto_in_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_in_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_in_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_in_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_6_auto_in_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_6_auto_in_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_in_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_out_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_out_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_out_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_6_auto_out_aw_bits_addr; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_out_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_out_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_6_auto_out_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_6_auto_out_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_out_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_out_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_out_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_out_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_6_auto_out_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_out_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_out_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_out_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_6_auto_out_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_6_auto_out_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_out_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_out_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_out_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_6_auto_out_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_6_auto_out_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_out_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_7_clock; // @[Buffer.scala 58:29]
  wire  axi4buf_7_reset; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_in_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_in_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_in_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_7_auto_in_aw_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_7_auto_in_aw_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_in_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_in_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_7_auto_in_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_7_auto_in_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_in_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_in_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_in_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_in_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_7_auto_in_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_in_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_in_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_in_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_7_auto_in_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_7_auto_in_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_in_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_in_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_in_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_7_auto_in_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_7_auto_in_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_in_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_out_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_out_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_out_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_7_auto_out_aw_bits_addr; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_out_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_out_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_7_auto_out_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_7_auto_out_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_out_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_out_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_out_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_out_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_7_auto_out_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_out_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_out_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_out_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_7_auto_out_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_7_auto_out_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_out_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_out_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_out_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_7_auto_out_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_7_auto_out_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_out_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_8_clock; // @[Buffer.scala 58:29]
  wire  axi4buf_8_reset; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_in_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_in_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_in_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_8_auto_in_aw_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_8_auto_in_aw_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_in_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_in_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_8_auto_in_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_8_auto_in_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_in_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_in_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_in_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_in_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_8_auto_in_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_in_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_in_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_in_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_8_auto_in_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_8_auto_in_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_in_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_in_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_in_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_8_auto_in_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_8_auto_in_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_in_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_out_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_out_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_out_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_8_auto_out_aw_bits_addr; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_out_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_out_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_8_auto_out_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_8_auto_out_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_out_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_out_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_out_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_out_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_8_auto_out_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_out_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_out_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_out_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_8_auto_out_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_8_auto_out_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_out_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_out_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_out_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_8_auto_out_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_8_auto_out_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_out_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_9_clock; // @[Buffer.scala 58:29]
  wire  axi4buf_9_reset; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_in_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_in_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_in_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_9_auto_in_aw_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_9_auto_in_aw_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_in_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_in_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_9_auto_in_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_9_auto_in_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_in_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_in_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_in_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_in_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_9_auto_in_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_in_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_in_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_in_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_9_auto_in_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_9_auto_in_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_in_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_in_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_in_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_9_auto_in_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_9_auto_in_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_in_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_out_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_out_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_out_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_9_auto_out_aw_bits_addr; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_out_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_out_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_9_auto_out_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_9_auto_out_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_out_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_out_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_out_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_out_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_9_auto_out_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_out_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_out_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_out_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_9_auto_out_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_9_auto_out_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_out_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_out_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_out_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_9_auto_out_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_9_auto_out_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_out_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_10_clock; // @[Buffer.scala 58:29]
  wire  axi4buf_10_reset; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_in_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_in_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_in_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_10_auto_in_aw_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_10_auto_in_aw_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_in_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_in_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_10_auto_in_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_10_auto_in_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_in_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_in_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_in_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_in_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_10_auto_in_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_in_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_in_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_in_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_10_auto_in_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_10_auto_in_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_in_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_in_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_in_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_10_auto_in_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_10_auto_in_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_in_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_out_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_out_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_out_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_10_auto_out_aw_bits_addr; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_out_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_out_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_10_auto_out_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_10_auto_out_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_out_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_out_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_out_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_out_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_10_auto_out_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_out_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_out_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_out_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_10_auto_out_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_10_auto_out_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_out_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_out_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_out_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_10_auto_out_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_10_auto_out_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_out_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_11_clock; // @[Buffer.scala 58:29]
  wire  axi4buf_11_reset; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_in_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_in_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_in_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_11_auto_in_aw_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_11_auto_in_aw_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_in_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_in_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_11_auto_in_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_11_auto_in_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_in_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_in_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_in_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_in_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_11_auto_in_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_in_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_in_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_in_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_11_auto_in_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_11_auto_in_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_in_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_in_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_in_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_11_auto_in_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_11_auto_in_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_in_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_out_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_out_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_out_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_11_auto_out_aw_bits_addr; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_out_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_out_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_11_auto_out_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_11_auto_out_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_out_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_out_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_out_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_out_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_11_auto_out_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_out_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_out_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_out_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_11_auto_out_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_11_auto_out_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_out_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_out_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_out_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_11_auto_out_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_11_auto_out_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_out_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_12_clock; // @[Buffer.scala 58:29]
  wire  axi4buf_12_reset; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_in_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_in_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_in_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_12_auto_in_aw_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_12_auto_in_aw_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_in_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_in_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_12_auto_in_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_12_auto_in_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_in_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_in_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_in_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_in_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_12_auto_in_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_in_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_in_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_in_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_12_auto_in_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_12_auto_in_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_in_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_in_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_in_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_12_auto_in_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_12_auto_in_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_in_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_out_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_out_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_out_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_12_auto_out_aw_bits_addr; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_out_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_out_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_12_auto_out_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_12_auto_out_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_out_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_out_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_out_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_out_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_12_auto_out_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_out_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_out_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_out_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_12_auto_out_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_12_auto_out_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_out_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_out_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_out_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_12_auto_out_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_12_auto_out_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_out_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_13_clock; // @[Buffer.scala 58:29]
  wire  axi4buf_13_reset; // @[Buffer.scala 58:29]
  wire  axi4buf_13_auto_in_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_13_auto_in_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_13_auto_in_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_13_auto_in_aw_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_13_auto_in_aw_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_13_auto_in_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_13_auto_in_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_13_auto_in_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_13_auto_in_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_13_auto_in_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_13_auto_in_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_13_auto_in_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_13_auto_in_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_13_auto_in_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_13_auto_in_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_13_auto_in_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_13_auto_in_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_13_auto_in_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_13_auto_in_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_13_auto_in_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_13_auto_in_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_13_auto_in_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_13_auto_in_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_13_auto_in_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_13_auto_in_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_13_auto_out_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_13_auto_out_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_13_auto_out_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_13_auto_out_aw_bits_addr; // @[Buffer.scala 58:29]
  wire  axi4buf_13_auto_out_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_13_auto_out_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_13_auto_out_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_13_auto_out_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_13_auto_out_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_13_auto_out_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_13_auto_out_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_13_auto_out_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_13_auto_out_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_13_auto_out_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_13_auto_out_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_13_auto_out_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_13_auto_out_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_13_auto_out_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_13_auto_out_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_13_auto_out_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_13_auto_out_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_13_auto_out_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_13_auto_out_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_13_auto_out_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_14_clock; // @[Buffer.scala 58:29]
  wire  axi4buf_14_reset; // @[Buffer.scala 58:29]
  wire  axi4buf_14_auto_in_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_14_auto_in_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_14_auto_in_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_14_auto_in_aw_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_14_auto_in_aw_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_14_auto_in_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_14_auto_in_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_14_auto_in_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_14_auto_in_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_14_auto_in_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_14_auto_in_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_14_auto_in_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_14_auto_in_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_14_auto_in_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_14_auto_in_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_14_auto_in_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_14_auto_in_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_14_auto_in_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_14_auto_in_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_14_auto_in_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_14_auto_in_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_14_auto_in_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_14_auto_in_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_14_auto_in_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_14_auto_in_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_14_auto_out_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_14_auto_out_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_14_auto_out_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_14_auto_out_aw_bits_addr; // @[Buffer.scala 58:29]
  wire  axi4buf_14_auto_out_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_14_auto_out_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_14_auto_out_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_14_auto_out_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_14_auto_out_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_14_auto_out_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_14_auto_out_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_14_auto_out_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_14_auto_out_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_14_auto_out_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_14_auto_out_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_14_auto_out_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_14_auto_out_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_14_auto_out_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_14_auto_out_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_14_auto_out_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_14_auto_out_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_14_auto_out_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_14_auto_out_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_14_auto_out_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_15_clock; // @[Buffer.scala 58:29]
  wire  axi4buf_15_reset; // @[Buffer.scala 58:29]
  wire  axi4buf_15_auto_in_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_15_auto_in_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_15_auto_in_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_15_auto_in_aw_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_15_auto_in_aw_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_15_auto_in_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_15_auto_in_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_15_auto_in_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_15_auto_in_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_15_auto_in_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_15_auto_in_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_15_auto_in_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_15_auto_in_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_15_auto_in_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_15_auto_in_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_15_auto_in_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_15_auto_in_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_15_auto_in_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_15_auto_in_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_15_auto_in_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_15_auto_in_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_15_auto_in_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_15_auto_in_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_15_auto_in_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_15_auto_in_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_15_auto_out_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_15_auto_out_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_15_auto_out_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_15_auto_out_aw_bits_addr; // @[Buffer.scala 58:29]
  wire  axi4buf_15_auto_out_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_15_auto_out_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_15_auto_out_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_15_auto_out_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_15_auto_out_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_15_auto_out_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_15_auto_out_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_15_auto_out_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_15_auto_out_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_15_auto_out_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_15_auto_out_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_15_auto_out_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_15_auto_out_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_15_auto_out_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_15_auto_out_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_15_auto_out_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_15_auto_out_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_15_auto_out_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_15_auto_out_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_15_auto_out_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_16_clock; // @[Buffer.scala 58:29]
  wire  axi4buf_16_reset; // @[Buffer.scala 58:29]
  wire  axi4buf_16_auto_in_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_16_auto_in_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_16_auto_in_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_16_auto_in_aw_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_16_auto_in_aw_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_16_auto_in_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_16_auto_in_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_16_auto_in_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_16_auto_in_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_16_auto_in_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_16_auto_in_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_16_auto_in_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_16_auto_in_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_16_auto_in_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_16_auto_in_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_16_auto_in_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_16_auto_in_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_16_auto_in_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_16_auto_in_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_16_auto_in_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_16_auto_in_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_16_auto_in_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_16_auto_in_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_16_auto_in_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_16_auto_in_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_16_auto_out_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_16_auto_out_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_16_auto_out_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_16_auto_out_aw_bits_addr; // @[Buffer.scala 58:29]
  wire  axi4buf_16_auto_out_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_16_auto_out_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_16_auto_out_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_16_auto_out_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_16_auto_out_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_16_auto_out_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_16_auto_out_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_16_auto_out_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_16_auto_out_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_16_auto_out_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_16_auto_out_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_16_auto_out_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_16_auto_out_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_16_auto_out_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_16_auto_out_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_16_auto_out_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_16_auto_out_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_16_auto_out_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_16_auto_out_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_16_auto_out_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_17_clock; // @[Buffer.scala 58:29]
  wire  axi4buf_17_reset; // @[Buffer.scala 58:29]
  wire  axi4buf_17_auto_in_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_17_auto_in_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_17_auto_in_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_17_auto_in_aw_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_17_auto_in_aw_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_17_auto_in_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_17_auto_in_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_17_auto_in_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_17_auto_in_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_17_auto_in_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_17_auto_in_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_17_auto_in_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_17_auto_in_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_17_auto_in_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_17_auto_in_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_17_auto_in_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_17_auto_in_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_17_auto_in_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_17_auto_in_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_17_auto_in_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_17_auto_in_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_17_auto_in_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_17_auto_in_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_17_auto_in_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_17_auto_in_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_17_auto_out_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_17_auto_out_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_17_auto_out_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_17_auto_out_aw_bits_addr; // @[Buffer.scala 58:29]
  wire  axi4buf_17_auto_out_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_17_auto_out_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_17_auto_out_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_17_auto_out_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_17_auto_out_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_17_auto_out_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_17_auto_out_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_17_auto_out_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_17_auto_out_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_17_auto_out_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_17_auto_out_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_17_auto_out_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_17_auto_out_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_17_auto_out_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_17_auto_out_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_17_auto_out_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_17_auto_out_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_17_auto_out_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_17_auto_out_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_17_auto_out_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_18_clock; // @[Buffer.scala 58:29]
  wire  axi4buf_18_reset; // @[Buffer.scala 58:29]
  wire  axi4buf_18_auto_in_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_18_auto_in_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_18_auto_in_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_18_auto_in_aw_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_18_auto_in_aw_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_18_auto_in_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_18_auto_in_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_18_auto_in_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_18_auto_in_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_18_auto_in_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_18_auto_in_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_18_auto_in_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_18_auto_in_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_18_auto_in_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_18_auto_in_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_18_auto_in_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_18_auto_in_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_18_auto_in_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_18_auto_in_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_18_auto_in_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_18_auto_in_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_18_auto_in_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_18_auto_in_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_18_auto_in_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_18_auto_in_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_18_auto_out_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_18_auto_out_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_18_auto_out_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_18_auto_out_aw_bits_addr; // @[Buffer.scala 58:29]
  wire  axi4buf_18_auto_out_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_18_auto_out_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_18_auto_out_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_18_auto_out_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_18_auto_out_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_18_auto_out_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_18_auto_out_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_18_auto_out_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_18_auto_out_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_18_auto_out_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_18_auto_out_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_18_auto_out_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_18_auto_out_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_18_auto_out_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_18_auto_out_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_18_auto_out_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_18_auto_out_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_18_auto_out_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_18_auto_out_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_18_auto_out_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_19_clock; // @[Buffer.scala 58:29]
  wire  axi4buf_19_reset; // @[Buffer.scala 58:29]
  wire  axi4buf_19_auto_in_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_19_auto_in_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_19_auto_in_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_19_auto_in_aw_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_19_auto_in_aw_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_19_auto_in_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_19_auto_in_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_19_auto_in_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_19_auto_in_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_19_auto_in_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_19_auto_in_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_19_auto_in_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_19_auto_in_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_19_auto_in_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_19_auto_in_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_19_auto_in_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_19_auto_in_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_19_auto_in_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_19_auto_in_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_19_auto_in_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_19_auto_in_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_19_auto_in_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_19_auto_in_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_19_auto_in_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_19_auto_in_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_19_auto_out_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_19_auto_out_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_19_auto_out_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_19_auto_out_aw_bits_addr; // @[Buffer.scala 58:29]
  wire  axi4buf_19_auto_out_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_19_auto_out_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_19_auto_out_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_19_auto_out_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_19_auto_out_w_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_19_auto_out_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_19_auto_out_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_19_auto_out_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_19_auto_out_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_19_auto_out_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_19_auto_out_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_19_auto_out_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_19_auto_out_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_19_auto_out_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_19_auto_out_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_19_auto_out_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_19_auto_out_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_19_auto_out_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_19_auto_out_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_19_auto_out_r_bits_last; // @[Buffer.scala 58:29]
  wire  buffer_clock; // @[Buffer.scala 29:28]
  wire  buffer_reset; // @[Buffer.scala 29:28]
  wire  buffer_auto_in_ready; // @[Buffer.scala 29:28]
  wire  buffer_auto_in_valid; // @[Buffer.scala 29:28]
  wire [31:0] buffer_auto_in_bits_data; // @[Buffer.scala 29:28]
  wire  buffer_auto_in_bits_last; // @[Buffer.scala 29:28]
  wire  buffer_auto_out_ready; // @[Buffer.scala 29:28]
  wire  buffer_auto_out_valid; // @[Buffer.scala 29:28]
  wire [31:0] buffer_auto_out_bits_data; // @[Buffer.scala 29:28]
  wire  buffer_auto_out_bits_last; // @[Buffer.scala 29:28]
  wire  buffer_1_clock; // @[Buffer.scala 29:28]
  wire  buffer_1_reset; // @[Buffer.scala 29:28]
  wire  buffer_1_auto_in_ready; // @[Buffer.scala 29:28]
  wire  buffer_1_auto_in_valid; // @[Buffer.scala 29:28]
  wire [31:0] buffer_1_auto_in_bits_data; // @[Buffer.scala 29:28]
  wire  buffer_1_auto_in_bits_last; // @[Buffer.scala 29:28]
  wire  buffer_1_auto_out_ready; // @[Buffer.scala 29:28]
  wire  buffer_1_auto_out_valid; // @[Buffer.scala 29:28]
  wire [31:0] buffer_1_auto_out_bits_data; // @[Buffer.scala 29:28]
  wire  buffer_1_auto_out_bits_last; // @[Buffer.scala 29:28]
  wire  buffer_2_clock; // @[Buffer.scala 29:28]
  wire  buffer_2_reset; // @[Buffer.scala 29:28]
  wire  buffer_2_auto_in_ready; // @[Buffer.scala 29:28]
  wire  buffer_2_auto_in_valid; // @[Buffer.scala 29:28]
  wire [31:0] buffer_2_auto_in_bits_data; // @[Buffer.scala 29:28]
  wire  buffer_2_auto_in_bits_last; // @[Buffer.scala 29:28]
  wire  buffer_2_auto_out_ready; // @[Buffer.scala 29:28]
  wire  buffer_2_auto_out_valid; // @[Buffer.scala 29:28]
  wire [31:0] buffer_2_auto_out_bits_data; // @[Buffer.scala 29:28]
  wire  buffer_2_auto_out_bits_last; // @[Buffer.scala 29:28]
  wire  buffer_3_clock; // @[Buffer.scala 29:28]
  wire  buffer_3_reset; // @[Buffer.scala 29:28]
  wire  buffer_3_auto_in_ready; // @[Buffer.scala 29:28]
  wire  buffer_3_auto_in_valid; // @[Buffer.scala 29:28]
  wire [31:0] buffer_3_auto_in_bits_data; // @[Buffer.scala 29:28]
  wire  buffer_3_auto_in_bits_last; // @[Buffer.scala 29:28]
  wire  buffer_3_auto_out_ready; // @[Buffer.scala 29:28]
  wire  buffer_3_auto_out_valid; // @[Buffer.scala 29:28]
  wire [31:0] buffer_3_auto_out_bits_data; // @[Buffer.scala 29:28]
  wire  buffer_3_auto_out_bits_last; // @[Buffer.scala 29:28]
  wire  buffer_4_clock; // @[Buffer.scala 29:28]
  wire  buffer_4_reset; // @[Buffer.scala 29:28]
  wire  buffer_4_auto_in_ready; // @[Buffer.scala 29:28]
  wire  buffer_4_auto_in_valid; // @[Buffer.scala 29:28]
  wire [31:0] buffer_4_auto_in_bits_data; // @[Buffer.scala 29:28]
  wire  buffer_4_auto_in_bits_last; // @[Buffer.scala 29:28]
  wire  buffer_4_auto_out_ready; // @[Buffer.scala 29:28]
  wire  buffer_4_auto_out_valid; // @[Buffer.scala 29:28]
  wire [31:0] buffer_4_auto_out_bits_data; // @[Buffer.scala 29:28]
  wire  buffer_4_auto_out_bits_last; // @[Buffer.scala 29:28]
  wire  buffer_5_clock; // @[Buffer.scala 29:28]
  wire  buffer_5_reset; // @[Buffer.scala 29:28]
  wire  buffer_5_auto_in_ready; // @[Buffer.scala 29:28]
  wire  buffer_5_auto_in_valid; // @[Buffer.scala 29:28]
  wire [31:0] buffer_5_auto_in_bits_data; // @[Buffer.scala 29:28]
  wire  buffer_5_auto_in_bits_last; // @[Buffer.scala 29:28]
  wire  buffer_5_auto_out_ready; // @[Buffer.scala 29:28]
  wire  buffer_5_auto_out_valid; // @[Buffer.scala 29:28]
  wire [31:0] buffer_5_auto_out_bits_data; // @[Buffer.scala 29:28]
  wire  buffer_5_auto_out_bits_last; // @[Buffer.scala 29:28]
  wire  buffer_6_clock; // @[Buffer.scala 29:28]
  wire  buffer_6_reset; // @[Buffer.scala 29:28]
  wire  buffer_6_auto_in_ready; // @[Buffer.scala 29:28]
  wire  buffer_6_auto_in_valid; // @[Buffer.scala 29:28]
  wire [31:0] buffer_6_auto_in_bits_data; // @[Buffer.scala 29:28]
  wire  buffer_6_auto_in_bits_last; // @[Buffer.scala 29:28]
  wire  buffer_6_auto_out_ready; // @[Buffer.scala 29:28]
  wire  buffer_6_auto_out_valid; // @[Buffer.scala 29:28]
  wire [31:0] buffer_6_auto_out_bits_data; // @[Buffer.scala 29:28]
  wire  buffer_6_auto_out_bits_last; // @[Buffer.scala 29:28]
  wire  buffer_7_clock; // @[Buffer.scala 29:28]
  wire  buffer_7_reset; // @[Buffer.scala 29:28]
  wire  buffer_7_auto_in_ready; // @[Buffer.scala 29:28]
  wire  buffer_7_auto_in_valid; // @[Buffer.scala 29:28]
  wire [31:0] buffer_7_auto_in_bits_data; // @[Buffer.scala 29:28]
  wire  buffer_7_auto_in_bits_last; // @[Buffer.scala 29:28]
  wire  buffer_7_auto_out_ready; // @[Buffer.scala 29:28]
  wire  buffer_7_auto_out_valid; // @[Buffer.scala 29:28]
  wire [31:0] buffer_7_auto_out_bits_data; // @[Buffer.scala 29:28]
  wire  buffer_7_auto_out_bits_last; // @[Buffer.scala 29:28]
  wire  buffer_8_clock; // @[Buffer.scala 29:28]
  wire  buffer_8_reset; // @[Buffer.scala 29:28]
  wire  buffer_8_auto_in_ready; // @[Buffer.scala 29:28]
  wire  buffer_8_auto_in_valid; // @[Buffer.scala 29:28]
  wire [31:0] buffer_8_auto_in_bits_data; // @[Buffer.scala 29:28]
  wire  buffer_8_auto_in_bits_last; // @[Buffer.scala 29:28]
  wire  buffer_8_auto_out_ready; // @[Buffer.scala 29:28]
  wire  buffer_8_auto_out_valid; // @[Buffer.scala 29:28]
  wire [31:0] buffer_8_auto_out_bits_data; // @[Buffer.scala 29:28]
  wire  buffer_8_auto_out_bits_last; // @[Buffer.scala 29:28]
  wire  buffer_9_clock; // @[Buffer.scala 29:28]
  wire  buffer_9_reset; // @[Buffer.scala 29:28]
  wire  buffer_9_auto_in_ready; // @[Buffer.scala 29:28]
  wire  buffer_9_auto_in_valid; // @[Buffer.scala 29:28]
  wire [31:0] buffer_9_auto_in_bits_data; // @[Buffer.scala 29:28]
  wire  buffer_9_auto_in_bits_last; // @[Buffer.scala 29:28]
  wire  buffer_9_auto_out_ready; // @[Buffer.scala 29:28]
  wire  buffer_9_auto_out_valid; // @[Buffer.scala 29:28]
  wire [31:0] buffer_9_auto_out_bits_data; // @[Buffer.scala 29:28]
  wire  buffer_9_auto_out_bits_last; // @[Buffer.scala 29:28]
  wire  converter_auto_in_aw_ready; // @[Node.scala 65:31]
  wire  converter_auto_in_aw_valid; // @[Node.scala 65:31]
  wire  converter_auto_in_aw_bits_id; // @[Node.scala 65:31]
  wire [31:0] converter_auto_in_aw_bits_addr; // @[Node.scala 65:31]
  wire [2:0] converter_auto_in_aw_bits_size; // @[Node.scala 65:31]
  wire  converter_auto_in_w_ready; // @[Node.scala 65:31]
  wire  converter_auto_in_w_valid; // @[Node.scala 65:31]
  wire [31:0] converter_auto_in_w_bits_data; // @[Node.scala 65:31]
  wire [3:0] converter_auto_in_w_bits_strb; // @[Node.scala 65:31]
  wire  converter_auto_in_w_bits_last; // @[Node.scala 65:31]
  wire  converter_auto_in_b_ready; // @[Node.scala 65:31]
  wire  converter_auto_in_b_valid; // @[Node.scala 65:31]
  wire [1:0] converter_auto_in_b_bits_resp; // @[Node.scala 65:31]
  wire  converter_auto_in_ar_ready; // @[Node.scala 65:31]
  wire  converter_auto_in_ar_valid; // @[Node.scala 65:31]
  wire  converter_auto_in_ar_bits_id; // @[Node.scala 65:31]
  wire [31:0] converter_auto_in_ar_bits_addr; // @[Node.scala 65:31]
  wire [2:0] converter_auto_in_ar_bits_size; // @[Node.scala 65:31]
  wire  converter_auto_in_r_ready; // @[Node.scala 65:31]
  wire  converter_auto_in_r_valid; // @[Node.scala 65:31]
  wire [31:0] converter_auto_in_r_bits_data; // @[Node.scala 65:31]
  wire [1:0] converter_auto_in_r_bits_resp; // @[Node.scala 65:31]
  wire  converter_auto_in_r_bits_last; // @[Node.scala 65:31]
  wire  converter_auto_out_aw_ready; // @[Node.scala 65:31]
  wire  converter_auto_out_aw_valid; // @[Node.scala 65:31]
  wire  converter_auto_out_aw_bits_id; // @[Node.scala 65:31]
  wire [29:0] converter_auto_out_aw_bits_addr; // @[Node.scala 65:31]
  wire [2:0] converter_auto_out_aw_bits_size; // @[Node.scala 65:31]
  wire  converter_auto_out_w_ready; // @[Node.scala 65:31]
  wire  converter_auto_out_w_valid; // @[Node.scala 65:31]
  wire [31:0] converter_auto_out_w_bits_data; // @[Node.scala 65:31]
  wire [3:0] converter_auto_out_w_bits_strb; // @[Node.scala 65:31]
  wire  converter_auto_out_w_bits_last; // @[Node.scala 65:31]
  wire  converter_auto_out_b_ready; // @[Node.scala 65:31]
  wire  converter_auto_out_b_valid; // @[Node.scala 65:31]
  wire [1:0] converter_auto_out_b_bits_resp; // @[Node.scala 65:31]
  wire  converter_auto_out_ar_ready; // @[Node.scala 65:31]
  wire  converter_auto_out_ar_valid; // @[Node.scala 65:31]
  wire  converter_auto_out_ar_bits_id; // @[Node.scala 65:31]
  wire [29:0] converter_auto_out_ar_bits_addr; // @[Node.scala 65:31]
  wire [2:0] converter_auto_out_ar_bits_size; // @[Node.scala 65:31]
  wire  converter_auto_out_r_ready; // @[Node.scala 65:31]
  wire  converter_auto_out_r_valid; // @[Node.scala 65:31]
  wire [31:0] converter_auto_out_r_bits_data; // @[Node.scala 65:31]
  wire [1:0] converter_auto_out_r_bits_resp; // @[Node.scala 65:31]
  wire  converter_auto_out_r_bits_last; // @[Node.scala 65:31]
  wire  converter_1_auto_in_ready; // @[Nodes.scala 165:31]
  wire  converter_1_auto_in_valid; // @[Nodes.scala 165:31]
  wire [7:0] converter_1_auto_in_bits_data; // @[Nodes.scala 165:31]
  wire  converter_1_auto_in_bits_last; // @[Nodes.scala 165:31]
  wire  converter_1_auto_out_ready; // @[Nodes.scala 165:31]
  wire  converter_1_auto_out_valid; // @[Nodes.scala 165:31]
  wire [7:0] converter_1_auto_out_bits_data; // @[Nodes.scala 165:31]
  wire  converter_1_auto_out_bits_last; // @[Nodes.scala 165:31]
  wire  converter_2_auto_in_ready; // @[Nodes.scala 201:31]
  wire  converter_2_auto_in_valid; // @[Nodes.scala 201:31]
  wire [7:0] converter_2_auto_in_bits_data; // @[Nodes.scala 201:31]
  wire  converter_2_auto_in_bits_last; // @[Nodes.scala 201:31]
  wire  converter_2_auto_out_ready; // @[Nodes.scala 201:31]
  wire  converter_2_auto_out_valid; // @[Nodes.scala 201:31]
  wire [7:0] converter_2_auto_out_bits_data; // @[Nodes.scala 201:31]
  wire  converter_2_auto_out_bits_last; // @[Nodes.scala 201:31]
  AXI4StreamWidthAdapater_4_to_1 widthAdapter ( // @[AXI4StreamWidthAdapter.scala 82:34]
    .clock(widthAdapter_clock),
    .reset(widthAdapter_reset),
    .auto_in_ready(widthAdapter_auto_in_ready),
    .auto_in_valid(widthAdapter_auto_in_valid),
    .auto_in_bits_data(widthAdapter_auto_in_bits_data),
    .auto_in_bits_last(widthAdapter_auto_in_bits_last),
    .auto_out_ready(widthAdapter_auto_out_ready),
    .auto_out_valid(widthAdapter_auto_out_valid),
    .auto_out_bits_data(widthAdapter_auto_out_bits_data),
    .auto_out_bits_last(widthAdapter_auto_out_bits_last)
  );
  AXI4Splitter in_split ( // @[SpectrometerTest.scala 114:29]
    .clock(in_split_clock),
    .reset(in_split_reset),
    .auto_mem_in_aw_ready(in_split_auto_mem_in_aw_ready),
    .auto_mem_in_aw_valid(in_split_auto_mem_in_aw_valid),
    .auto_mem_in_aw_bits_id(in_split_auto_mem_in_aw_bits_id),
    .auto_mem_in_aw_bits_addr(in_split_auto_mem_in_aw_bits_addr),
    .auto_mem_in_w_ready(in_split_auto_mem_in_w_ready),
    .auto_mem_in_w_valid(in_split_auto_mem_in_w_valid),
    .auto_mem_in_w_bits_data(in_split_auto_mem_in_w_bits_data),
    .auto_mem_in_w_bits_strb(in_split_auto_mem_in_w_bits_strb),
    .auto_mem_in_b_ready(in_split_auto_mem_in_b_ready),
    .auto_mem_in_b_valid(in_split_auto_mem_in_b_valid),
    .auto_mem_in_b_bits_id(in_split_auto_mem_in_b_bits_id),
    .auto_mem_in_ar_ready(in_split_auto_mem_in_ar_ready),
    .auto_mem_in_ar_valid(in_split_auto_mem_in_ar_valid),
    .auto_mem_in_ar_bits_id(in_split_auto_mem_in_ar_bits_id),
    .auto_mem_in_ar_bits_addr(in_split_auto_mem_in_ar_bits_addr),
    .auto_mem_in_ar_bits_size(in_split_auto_mem_in_ar_bits_size),
    .auto_mem_in_r_ready(in_split_auto_mem_in_r_ready),
    .auto_mem_in_r_valid(in_split_auto_mem_in_r_valid),
    .auto_mem_in_r_bits_id(in_split_auto_mem_in_r_bits_id),
    .auto_mem_in_r_bits_data(in_split_auto_mem_in_r_bits_data),
    .auto_stream_in_ready(in_split_auto_stream_in_ready),
    .auto_stream_in_valid(in_split_auto_stream_in_valid),
    .auto_stream_in_bits_data(in_split_auto_stream_in_bits_data),
    .auto_stream_in_bits_last(in_split_auto_stream_in_bits_last),
    .auto_stream_out_4_ready(in_split_auto_stream_out_4_ready),
    .auto_stream_out_4_valid(in_split_auto_stream_out_4_valid),
    .auto_stream_out_4_bits_data(in_split_auto_stream_out_4_bits_data),
    .auto_stream_out_4_bits_last(in_split_auto_stream_out_4_bits_last),
    .auto_stream_out_3_ready(in_split_auto_stream_out_3_ready),
    .auto_stream_out_3_valid(in_split_auto_stream_out_3_valid),
    .auto_stream_out_3_bits_data(in_split_auto_stream_out_3_bits_data),
    .auto_stream_out_3_bits_last(in_split_auto_stream_out_3_bits_last),
    .auto_stream_out_2_ready(in_split_auto_stream_out_2_ready),
    .auto_stream_out_2_valid(in_split_auto_stream_out_2_valid),
    .auto_stream_out_2_bits_data(in_split_auto_stream_out_2_bits_data),
    .auto_stream_out_2_bits_last(in_split_auto_stream_out_2_bits_last),
    .auto_stream_out_1_ready(in_split_auto_stream_out_1_ready),
    .auto_stream_out_1_valid(in_split_auto_stream_out_1_valid),
    .auto_stream_out_1_bits_data(in_split_auto_stream_out_1_bits_data),
    .auto_stream_out_1_bits_last(in_split_auto_stream_out_1_bits_last),
    .auto_stream_out_0_ready(in_split_auto_stream_out_0_ready),
    .auto_stream_out_0_valid(in_split_auto_stream_out_0_valid),
    .auto_stream_out_0_bits_data(in_split_auto_stream_out_0_bits_data),
    .auto_stream_out_0_bits_last(in_split_auto_stream_out_0_bits_last)
  );
  StreamBuffer in_queue ( // @[SpectrometerTest.scala 115:29]
    .clock(in_queue_clock),
    .reset(in_queue_reset),
    .auto_out_out_ready(in_queue_auto_out_out_ready),
    .auto_out_out_valid(in_queue_auto_out_out_valid),
    .auto_out_out_bits_data(in_queue_auto_out_out_bits_data),
    .auto_out_out_bits_last(in_queue_auto_out_out_bits_last),
    .auto_in_in_ready(in_queue_auto_in_in_ready),
    .auto_in_in_valid(in_queue_auto_in_in_valid),
    .auto_in_in_bits_data(in_queue_auto_in_in_bits_data),
    .auto_in_in_bits_last(in_queue_auto_in_in_bits_last)
  );
  PLFGDspBlockMem plfg ( // @[SpectrometerTest.scala 117:30]
    .clock(plfg_clock),
    .reset(plfg_reset),
    .auto_mem_in_aw_ready(plfg_auto_mem_in_aw_ready),
    .auto_mem_in_aw_valid(plfg_auto_mem_in_aw_valid),
    .auto_mem_in_aw_bits_id(plfg_auto_mem_in_aw_bits_id),
    .auto_mem_in_aw_bits_addr(plfg_auto_mem_in_aw_bits_addr),
    .auto_mem_in_w_ready(plfg_auto_mem_in_w_ready),
    .auto_mem_in_w_valid(plfg_auto_mem_in_w_valid),
    .auto_mem_in_w_bits_data(plfg_auto_mem_in_w_bits_data),
    .auto_mem_in_w_bits_strb(plfg_auto_mem_in_w_bits_strb),
    .auto_mem_in_w_bits_last(plfg_auto_mem_in_w_bits_last),
    .auto_mem_in_b_ready(plfg_auto_mem_in_b_ready),
    .auto_mem_in_b_valid(plfg_auto_mem_in_b_valid),
    .auto_mem_in_b_bits_resp(plfg_auto_mem_in_b_bits_resp),
    .auto_mem_in_ar_ready(plfg_auto_mem_in_ar_ready),
    .auto_mem_in_ar_valid(plfg_auto_mem_in_ar_valid),
    .auto_mem_in_ar_bits_id(plfg_auto_mem_in_ar_bits_id),
    .auto_mem_in_ar_bits_addr(plfg_auto_mem_in_ar_bits_addr),
    .auto_mem_in_ar_bits_size(plfg_auto_mem_in_ar_bits_size),
    .auto_mem_in_r_ready(plfg_auto_mem_in_r_ready),
    .auto_mem_in_r_valid(plfg_auto_mem_in_r_valid),
    .auto_mem_in_r_bits_data(plfg_auto_mem_in_r_bits_data),
    .auto_mem_in_r_bits_resp(plfg_auto_mem_in_r_bits_resp),
    .auto_mem_in_r_bits_last(plfg_auto_mem_in_r_bits_last),
    .auto_stream_out_ready(plfg_auto_stream_out_ready),
    .auto_stream_out_valid(plfg_auto_stream_out_valid),
    .auto_stream_out_bits_data(plfg_auto_stream_out_bits_data),
    .auto_stream_out_bits_last(plfg_auto_stream_out_bits_last)
  );
  AXI4Splitter_1 plfg_split ( // @[SpectrometerTest.scala 118:30]
    .clock(plfg_split_clock),
    .reset(plfg_split_reset),
    .auto_mem_in_aw_ready(plfg_split_auto_mem_in_aw_ready),
    .auto_mem_in_aw_valid(plfg_split_auto_mem_in_aw_valid),
    .auto_mem_in_aw_bits_id(plfg_split_auto_mem_in_aw_bits_id),
    .auto_mem_in_aw_bits_addr(plfg_split_auto_mem_in_aw_bits_addr),
    .auto_mem_in_w_ready(plfg_split_auto_mem_in_w_ready),
    .auto_mem_in_w_valid(plfg_split_auto_mem_in_w_valid),
    .auto_mem_in_w_bits_data(plfg_split_auto_mem_in_w_bits_data),
    .auto_mem_in_w_bits_strb(plfg_split_auto_mem_in_w_bits_strb),
    .auto_mem_in_b_ready(plfg_split_auto_mem_in_b_ready),
    .auto_mem_in_b_valid(plfg_split_auto_mem_in_b_valid),
    .auto_mem_in_b_bits_id(plfg_split_auto_mem_in_b_bits_id),
    .auto_mem_in_ar_ready(plfg_split_auto_mem_in_ar_ready),
    .auto_mem_in_ar_valid(plfg_split_auto_mem_in_ar_valid),
    .auto_mem_in_ar_bits_id(plfg_split_auto_mem_in_ar_bits_id),
    .auto_mem_in_ar_bits_addr(plfg_split_auto_mem_in_ar_bits_addr),
    .auto_mem_in_ar_bits_size(plfg_split_auto_mem_in_ar_bits_size),
    .auto_mem_in_r_ready(plfg_split_auto_mem_in_r_ready),
    .auto_mem_in_r_valid(plfg_split_auto_mem_in_r_valid),
    .auto_mem_in_r_bits_id(plfg_split_auto_mem_in_r_bits_id),
    .auto_mem_in_r_bits_data(plfg_split_auto_mem_in_r_bits_data),
    .auto_stream_in_ready(plfg_split_auto_stream_in_ready),
    .auto_stream_in_valid(plfg_split_auto_stream_in_valid),
    .auto_stream_in_bits_data(plfg_split_auto_stream_in_bits_data),
    .auto_stream_in_bits_last(plfg_split_auto_stream_in_bits_last),
    .auto_stream_out_1_ready(plfg_split_auto_stream_out_1_ready),
    .auto_stream_out_1_valid(plfg_split_auto_stream_out_1_valid),
    .auto_stream_out_1_bits_data(plfg_split_auto_stream_out_1_bits_data),
    .auto_stream_out_1_bits_last(plfg_split_auto_stream_out_1_bits_last),
    .auto_stream_out_0_ready(plfg_split_auto_stream_out_0_ready),
    .auto_stream_out_0_valid(plfg_split_auto_stream_out_0_valid),
    .auto_stream_out_0_bits_data(plfg_split_auto_stream_out_0_bits_data),
    .auto_stream_out_0_bits_last(plfg_split_auto_stream_out_0_bits_last)
  );
  AXI4StreamMux plfg_mux_0 ( // @[SpectrometerTest.scala 119:30]
    .clock(plfg_mux_0_clock),
    .reset(plfg_mux_0_reset),
    .auto_register_in_aw_ready(plfg_mux_0_auto_register_in_aw_ready),
    .auto_register_in_aw_valid(plfg_mux_0_auto_register_in_aw_valid),
    .auto_register_in_aw_bits_id(plfg_mux_0_auto_register_in_aw_bits_id),
    .auto_register_in_aw_bits_addr(plfg_mux_0_auto_register_in_aw_bits_addr),
    .auto_register_in_w_ready(plfg_mux_0_auto_register_in_w_ready),
    .auto_register_in_w_valid(plfg_mux_0_auto_register_in_w_valid),
    .auto_register_in_w_bits_data(plfg_mux_0_auto_register_in_w_bits_data),
    .auto_register_in_w_bits_strb(plfg_mux_0_auto_register_in_w_bits_strb),
    .auto_register_in_b_ready(plfg_mux_0_auto_register_in_b_ready),
    .auto_register_in_b_valid(plfg_mux_0_auto_register_in_b_valid),
    .auto_register_in_b_bits_id(plfg_mux_0_auto_register_in_b_bits_id),
    .auto_register_in_ar_ready(plfg_mux_0_auto_register_in_ar_ready),
    .auto_register_in_ar_valid(plfg_mux_0_auto_register_in_ar_valid),
    .auto_register_in_ar_bits_id(plfg_mux_0_auto_register_in_ar_bits_id),
    .auto_register_in_ar_bits_addr(plfg_mux_0_auto_register_in_ar_bits_addr),
    .auto_register_in_ar_bits_size(plfg_mux_0_auto_register_in_ar_bits_size),
    .auto_register_in_r_ready(plfg_mux_0_auto_register_in_r_ready),
    .auto_register_in_r_valid(plfg_mux_0_auto_register_in_r_valid),
    .auto_register_in_r_bits_id(plfg_mux_0_auto_register_in_r_bits_id),
    .auto_register_in_r_bits_data(plfg_mux_0_auto_register_in_r_bits_data),
    .auto_stream_in_2_ready(plfg_mux_0_auto_stream_in_2_ready),
    .auto_stream_in_2_valid(plfg_mux_0_auto_stream_in_2_valid),
    .auto_stream_in_2_bits_data(plfg_mux_0_auto_stream_in_2_bits_data),
    .auto_stream_in_2_bits_last(plfg_mux_0_auto_stream_in_2_bits_last),
    .auto_stream_in_1_ready(plfg_mux_0_auto_stream_in_1_ready),
    .auto_stream_in_1_valid(plfg_mux_0_auto_stream_in_1_valid),
    .auto_stream_in_1_bits_data(plfg_mux_0_auto_stream_in_1_bits_data),
    .auto_stream_in_1_bits_last(plfg_mux_0_auto_stream_in_1_bits_last),
    .auto_stream_in_0_ready(plfg_mux_0_auto_stream_in_0_ready),
    .auto_stream_in_0_valid(plfg_mux_0_auto_stream_in_0_valid),
    .auto_stream_in_0_bits_data(plfg_mux_0_auto_stream_in_0_bits_data),
    .auto_stream_in_0_bits_last(plfg_mux_0_auto_stream_in_0_bits_last),
    .auto_stream_out_0_ready(plfg_mux_0_auto_stream_out_0_ready),
    .auto_stream_out_0_valid(plfg_mux_0_auto_stream_out_0_valid),
    .auto_stream_out_0_bits_data(plfg_mux_0_auto_stream_out_0_bits_data),
    .auto_stream_out_0_bits_last(plfg_mux_0_auto_stream_out_0_bits_last)
  );
  AXI4StreamMux_1 plfg_mux_1 ( // @[SpectrometerTest.scala 120:30]
    .clock(plfg_mux_1_clock),
    .reset(plfg_mux_1_reset),
    .auto_register_in_aw_ready(plfg_mux_1_auto_register_in_aw_ready),
    .auto_register_in_aw_valid(plfg_mux_1_auto_register_in_aw_valid),
    .auto_register_in_aw_bits_id(plfg_mux_1_auto_register_in_aw_bits_id),
    .auto_register_in_aw_bits_addr(plfg_mux_1_auto_register_in_aw_bits_addr),
    .auto_register_in_w_ready(plfg_mux_1_auto_register_in_w_ready),
    .auto_register_in_w_valid(plfg_mux_1_auto_register_in_w_valid),
    .auto_register_in_w_bits_data(plfg_mux_1_auto_register_in_w_bits_data),
    .auto_register_in_w_bits_strb(plfg_mux_1_auto_register_in_w_bits_strb),
    .auto_register_in_b_ready(plfg_mux_1_auto_register_in_b_ready),
    .auto_register_in_b_valid(plfg_mux_1_auto_register_in_b_valid),
    .auto_register_in_b_bits_id(plfg_mux_1_auto_register_in_b_bits_id),
    .auto_register_in_ar_ready(plfg_mux_1_auto_register_in_ar_ready),
    .auto_register_in_ar_valid(plfg_mux_1_auto_register_in_ar_valid),
    .auto_register_in_ar_bits_id(plfg_mux_1_auto_register_in_ar_bits_id),
    .auto_register_in_ar_bits_addr(plfg_mux_1_auto_register_in_ar_bits_addr),
    .auto_register_in_ar_bits_size(plfg_mux_1_auto_register_in_ar_bits_size),
    .auto_register_in_r_ready(plfg_mux_1_auto_register_in_r_ready),
    .auto_register_in_r_valid(plfg_mux_1_auto_register_in_r_valid),
    .auto_register_in_r_bits_id(plfg_mux_1_auto_register_in_r_bits_id),
    .auto_register_in_r_bits_data(plfg_mux_1_auto_register_in_r_bits_data),
    .auto_stream_in_ready(plfg_mux_1_auto_stream_in_ready),
    .auto_stream_in_valid(plfg_mux_1_auto_stream_in_valid),
    .auto_stream_in_bits_data(plfg_mux_1_auto_stream_in_bits_data),
    .auto_stream_in_bits_last(plfg_mux_1_auto_stream_in_bits_last),
    .auto_stream_out_1_ready(plfg_mux_1_auto_stream_out_1_ready),
    .auto_stream_out_1_valid(plfg_mux_1_auto_stream_out_1_valid),
    .auto_stream_out_1_bits_data(plfg_mux_1_auto_stream_out_1_bits_data),
    .auto_stream_out_1_bits_last(plfg_mux_1_auto_stream_out_1_bits_last)
  );
  AXI4NCOLazyModuleBlock nco ( // @[SpectrometerTest.scala 126:29]
    .clock(nco_clock),
    .reset(nco_reset),
    .auto_stream_out_ready(nco_auto_stream_out_ready),
    .auto_stream_out_valid(nco_auto_stream_out_valid),
    .auto_stream_out_bits_data(nco_auto_stream_out_bits_data),
    .auto_stream_out_bits_last(nco_auto_stream_out_bits_last),
    .auto_freq_in_ready(nco_auto_freq_in_ready),
    .auto_freq_in_valid(nco_auto_freq_in_valid),
    .auto_freq_in_bits_data(nco_auto_freq_in_bits_data),
    .auto_freq_in_bits_last(nco_auto_freq_in_bits_last)
  );
  AXI4Splitter_2 nco_split ( // @[SpectrometerTest.scala 127:29]
    .clock(nco_split_clock),
    .reset(nco_split_reset),
    .auto_mem_in_aw_ready(nco_split_auto_mem_in_aw_ready),
    .auto_mem_in_aw_valid(nco_split_auto_mem_in_aw_valid),
    .auto_mem_in_aw_bits_id(nco_split_auto_mem_in_aw_bits_id),
    .auto_mem_in_aw_bits_addr(nco_split_auto_mem_in_aw_bits_addr),
    .auto_mem_in_w_ready(nco_split_auto_mem_in_w_ready),
    .auto_mem_in_w_valid(nco_split_auto_mem_in_w_valid),
    .auto_mem_in_w_bits_data(nco_split_auto_mem_in_w_bits_data),
    .auto_mem_in_w_bits_strb(nco_split_auto_mem_in_w_bits_strb),
    .auto_mem_in_b_ready(nco_split_auto_mem_in_b_ready),
    .auto_mem_in_b_valid(nco_split_auto_mem_in_b_valid),
    .auto_mem_in_b_bits_id(nco_split_auto_mem_in_b_bits_id),
    .auto_mem_in_ar_ready(nco_split_auto_mem_in_ar_ready),
    .auto_mem_in_ar_valid(nco_split_auto_mem_in_ar_valid),
    .auto_mem_in_ar_bits_id(nco_split_auto_mem_in_ar_bits_id),
    .auto_mem_in_ar_bits_addr(nco_split_auto_mem_in_ar_bits_addr),
    .auto_mem_in_ar_bits_size(nco_split_auto_mem_in_ar_bits_size),
    .auto_mem_in_r_ready(nco_split_auto_mem_in_r_ready),
    .auto_mem_in_r_valid(nco_split_auto_mem_in_r_valid),
    .auto_mem_in_r_bits_id(nco_split_auto_mem_in_r_bits_id),
    .auto_mem_in_r_bits_data(nco_split_auto_mem_in_r_bits_data),
    .auto_stream_in_ready(nco_split_auto_stream_in_ready),
    .auto_stream_in_valid(nco_split_auto_stream_in_valid),
    .auto_stream_in_bits_data(nco_split_auto_stream_in_bits_data),
    .auto_stream_in_bits_last(nco_split_auto_stream_in_bits_last),
    .auto_stream_out_1_ready(nco_split_auto_stream_out_1_ready),
    .auto_stream_out_1_valid(nco_split_auto_stream_out_1_valid),
    .auto_stream_out_1_bits_data(nco_split_auto_stream_out_1_bits_data),
    .auto_stream_out_1_bits_last(nco_split_auto_stream_out_1_bits_last),
    .auto_stream_out_0_ready(nco_split_auto_stream_out_0_ready),
    .auto_stream_out_0_valid(nco_split_auto_stream_out_0_valid),
    .auto_stream_out_0_bits_data(nco_split_auto_stream_out_0_bits_data),
    .auto_stream_out_0_bits_last(nco_split_auto_stream_out_0_bits_last)
  );
  AXI4StreamMux_2 nco_mux_0 ( // @[SpectrometerTest.scala 128:29]
    .clock(nco_mux_0_clock),
    .reset(nco_mux_0_reset),
    .auto_register_in_aw_ready(nco_mux_0_auto_register_in_aw_ready),
    .auto_register_in_aw_valid(nco_mux_0_auto_register_in_aw_valid),
    .auto_register_in_aw_bits_id(nco_mux_0_auto_register_in_aw_bits_id),
    .auto_register_in_aw_bits_addr(nco_mux_0_auto_register_in_aw_bits_addr),
    .auto_register_in_w_ready(nco_mux_0_auto_register_in_w_ready),
    .auto_register_in_w_valid(nco_mux_0_auto_register_in_w_valid),
    .auto_register_in_w_bits_data(nco_mux_0_auto_register_in_w_bits_data),
    .auto_register_in_w_bits_strb(nco_mux_0_auto_register_in_w_bits_strb),
    .auto_register_in_b_ready(nco_mux_0_auto_register_in_b_ready),
    .auto_register_in_b_valid(nco_mux_0_auto_register_in_b_valid),
    .auto_register_in_b_bits_id(nco_mux_0_auto_register_in_b_bits_id),
    .auto_register_in_ar_ready(nco_mux_0_auto_register_in_ar_ready),
    .auto_register_in_ar_valid(nco_mux_0_auto_register_in_ar_valid),
    .auto_register_in_ar_bits_id(nco_mux_0_auto_register_in_ar_bits_id),
    .auto_register_in_ar_bits_addr(nco_mux_0_auto_register_in_ar_bits_addr),
    .auto_register_in_ar_bits_size(nco_mux_0_auto_register_in_ar_bits_size),
    .auto_register_in_r_ready(nco_mux_0_auto_register_in_r_ready),
    .auto_register_in_r_valid(nco_mux_0_auto_register_in_r_valid),
    .auto_register_in_r_bits_id(nco_mux_0_auto_register_in_r_bits_id),
    .auto_register_in_r_bits_data(nco_mux_0_auto_register_in_r_bits_data),
    .auto_stream_in_2_ready(nco_mux_0_auto_stream_in_2_ready),
    .auto_stream_in_2_valid(nco_mux_0_auto_stream_in_2_valid),
    .auto_stream_in_2_bits_data(nco_mux_0_auto_stream_in_2_bits_data),
    .auto_stream_in_2_bits_last(nco_mux_0_auto_stream_in_2_bits_last),
    .auto_stream_in_1_ready(nco_mux_0_auto_stream_in_1_ready),
    .auto_stream_in_1_valid(nco_mux_0_auto_stream_in_1_valid),
    .auto_stream_in_1_bits_data(nco_mux_0_auto_stream_in_1_bits_data),
    .auto_stream_in_1_bits_last(nco_mux_0_auto_stream_in_1_bits_last),
    .auto_stream_in_0_ready(nco_mux_0_auto_stream_in_0_ready),
    .auto_stream_in_0_valid(nco_mux_0_auto_stream_in_0_valid),
    .auto_stream_in_0_bits_data(nco_mux_0_auto_stream_in_0_bits_data),
    .auto_stream_in_0_bits_last(nco_mux_0_auto_stream_in_0_bits_last),
    .auto_stream_out_0_ready(nco_mux_0_auto_stream_out_0_ready),
    .auto_stream_out_0_valid(nco_mux_0_auto_stream_out_0_valid),
    .auto_stream_out_0_bits_data(nco_mux_0_auto_stream_out_0_bits_data),
    .auto_stream_out_0_bits_last(nco_mux_0_auto_stream_out_0_bits_last)
  );
  AXI4StreamMux_1 nco_mux_1 ( // @[SpectrometerTest.scala 129:29]
    .clock(nco_mux_1_clock),
    .reset(nco_mux_1_reset),
    .auto_register_in_aw_ready(nco_mux_1_auto_register_in_aw_ready),
    .auto_register_in_aw_valid(nco_mux_1_auto_register_in_aw_valid),
    .auto_register_in_aw_bits_id(nco_mux_1_auto_register_in_aw_bits_id),
    .auto_register_in_aw_bits_addr(nco_mux_1_auto_register_in_aw_bits_addr),
    .auto_register_in_w_ready(nco_mux_1_auto_register_in_w_ready),
    .auto_register_in_w_valid(nco_mux_1_auto_register_in_w_valid),
    .auto_register_in_w_bits_data(nco_mux_1_auto_register_in_w_bits_data),
    .auto_register_in_w_bits_strb(nco_mux_1_auto_register_in_w_bits_strb),
    .auto_register_in_b_ready(nco_mux_1_auto_register_in_b_ready),
    .auto_register_in_b_valid(nco_mux_1_auto_register_in_b_valid),
    .auto_register_in_b_bits_id(nco_mux_1_auto_register_in_b_bits_id),
    .auto_register_in_ar_ready(nco_mux_1_auto_register_in_ar_ready),
    .auto_register_in_ar_valid(nco_mux_1_auto_register_in_ar_valid),
    .auto_register_in_ar_bits_id(nco_mux_1_auto_register_in_ar_bits_id),
    .auto_register_in_ar_bits_addr(nco_mux_1_auto_register_in_ar_bits_addr),
    .auto_register_in_ar_bits_size(nco_mux_1_auto_register_in_ar_bits_size),
    .auto_register_in_r_ready(nco_mux_1_auto_register_in_r_ready),
    .auto_register_in_r_valid(nco_mux_1_auto_register_in_r_valid),
    .auto_register_in_r_bits_id(nco_mux_1_auto_register_in_r_bits_id),
    .auto_register_in_r_bits_data(nco_mux_1_auto_register_in_r_bits_data),
    .auto_stream_in_ready(nco_mux_1_auto_stream_in_ready),
    .auto_stream_in_valid(nco_mux_1_auto_stream_in_valid),
    .auto_stream_in_bits_data(nco_mux_1_auto_stream_in_bits_data),
    .auto_stream_in_bits_last(nco_mux_1_auto_stream_in_bits_last),
    .auto_stream_out_1_ready(nco_mux_1_auto_stream_out_1_ready),
    .auto_stream_out_1_valid(nco_mux_1_auto_stream_out_1_valid),
    .auto_stream_out_1_bits_data(nco_mux_1_auto_stream_out_1_bits_data),
    .auto_stream_out_1_bits_last(nco_mux_1_auto_stream_out_1_bits_last)
  );
  AXI4FFTBlock fft ( // @[SpectrometerTest.scala 135:29]
    .clock(fft_clock),
    .reset(fft_reset),
    .auto_mem_in_aw_ready(fft_auto_mem_in_aw_ready),
    .auto_mem_in_aw_valid(fft_auto_mem_in_aw_valid),
    .auto_mem_in_aw_bits_id(fft_auto_mem_in_aw_bits_id),
    .auto_mem_in_aw_bits_addr(fft_auto_mem_in_aw_bits_addr),
    .auto_mem_in_w_ready(fft_auto_mem_in_w_ready),
    .auto_mem_in_w_valid(fft_auto_mem_in_w_valid),
    .auto_mem_in_w_bits_data(fft_auto_mem_in_w_bits_data),
    .auto_mem_in_w_bits_strb(fft_auto_mem_in_w_bits_strb),
    .auto_mem_in_b_ready(fft_auto_mem_in_b_ready),
    .auto_mem_in_b_valid(fft_auto_mem_in_b_valid),
    .auto_mem_in_b_bits_id(fft_auto_mem_in_b_bits_id),
    .auto_mem_in_ar_ready(fft_auto_mem_in_ar_ready),
    .auto_mem_in_ar_valid(fft_auto_mem_in_ar_valid),
    .auto_mem_in_ar_bits_id(fft_auto_mem_in_ar_bits_id),
    .auto_mem_in_ar_bits_addr(fft_auto_mem_in_ar_bits_addr),
    .auto_mem_in_ar_bits_size(fft_auto_mem_in_ar_bits_size),
    .auto_mem_in_r_ready(fft_auto_mem_in_r_ready),
    .auto_mem_in_r_valid(fft_auto_mem_in_r_valid),
    .auto_mem_in_r_bits_id(fft_auto_mem_in_r_bits_id),
    .auto_mem_in_r_bits_data(fft_auto_mem_in_r_bits_data),
    .auto_stream_in_ready(fft_auto_stream_in_ready),
    .auto_stream_in_valid(fft_auto_stream_in_valid),
    .auto_stream_in_bits_data(fft_auto_stream_in_bits_data),
    .auto_stream_in_bits_last(fft_auto_stream_in_bits_last),
    .auto_stream_out_ready(fft_auto_stream_out_ready),
    .auto_stream_out_valid(fft_auto_stream_out_valid),
    .auto_stream_out_bits_data(fft_auto_stream_out_bits_data),
    .auto_stream_out_bits_last(fft_auto_stream_out_bits_last)
  );
  AXI4Splitter_3 fft_split ( // @[SpectrometerTest.scala 136:29]
    .clock(fft_split_clock),
    .reset(fft_split_reset),
    .auto_mem_in_aw_ready(fft_split_auto_mem_in_aw_ready),
    .auto_mem_in_aw_valid(fft_split_auto_mem_in_aw_valid),
    .auto_mem_in_aw_bits_id(fft_split_auto_mem_in_aw_bits_id),
    .auto_mem_in_aw_bits_addr(fft_split_auto_mem_in_aw_bits_addr),
    .auto_mem_in_w_ready(fft_split_auto_mem_in_w_ready),
    .auto_mem_in_w_valid(fft_split_auto_mem_in_w_valid),
    .auto_mem_in_w_bits_data(fft_split_auto_mem_in_w_bits_data),
    .auto_mem_in_w_bits_strb(fft_split_auto_mem_in_w_bits_strb),
    .auto_mem_in_b_ready(fft_split_auto_mem_in_b_ready),
    .auto_mem_in_b_valid(fft_split_auto_mem_in_b_valid),
    .auto_mem_in_b_bits_id(fft_split_auto_mem_in_b_bits_id),
    .auto_mem_in_ar_ready(fft_split_auto_mem_in_ar_ready),
    .auto_mem_in_ar_valid(fft_split_auto_mem_in_ar_valid),
    .auto_mem_in_ar_bits_id(fft_split_auto_mem_in_ar_bits_id),
    .auto_mem_in_ar_bits_addr(fft_split_auto_mem_in_ar_bits_addr),
    .auto_mem_in_ar_bits_size(fft_split_auto_mem_in_ar_bits_size),
    .auto_mem_in_r_ready(fft_split_auto_mem_in_r_ready),
    .auto_mem_in_r_valid(fft_split_auto_mem_in_r_valid),
    .auto_mem_in_r_bits_id(fft_split_auto_mem_in_r_bits_id),
    .auto_mem_in_r_bits_data(fft_split_auto_mem_in_r_bits_data),
    .auto_stream_in_ready(fft_split_auto_stream_in_ready),
    .auto_stream_in_valid(fft_split_auto_stream_in_valid),
    .auto_stream_in_bits_data(fft_split_auto_stream_in_bits_data),
    .auto_stream_in_bits_last(fft_split_auto_stream_in_bits_last),
    .auto_stream_out_1_ready(fft_split_auto_stream_out_1_ready),
    .auto_stream_out_1_valid(fft_split_auto_stream_out_1_valid),
    .auto_stream_out_1_bits_data(fft_split_auto_stream_out_1_bits_data),
    .auto_stream_out_1_bits_last(fft_split_auto_stream_out_1_bits_last),
    .auto_stream_out_0_ready(fft_split_auto_stream_out_0_ready),
    .auto_stream_out_0_valid(fft_split_auto_stream_out_0_valid),
    .auto_stream_out_0_bits_data(fft_split_auto_stream_out_0_bits_data),
    .auto_stream_out_0_bits_last(fft_split_auto_stream_out_0_bits_last)
  );
  AXI4StreamMux_4 fft_mux_0 ( // @[SpectrometerTest.scala 137:29]
    .clock(fft_mux_0_clock),
    .reset(fft_mux_0_reset),
    .auto_register_in_aw_ready(fft_mux_0_auto_register_in_aw_ready),
    .auto_register_in_aw_valid(fft_mux_0_auto_register_in_aw_valid),
    .auto_register_in_aw_bits_id(fft_mux_0_auto_register_in_aw_bits_id),
    .auto_register_in_aw_bits_addr(fft_mux_0_auto_register_in_aw_bits_addr),
    .auto_register_in_w_ready(fft_mux_0_auto_register_in_w_ready),
    .auto_register_in_w_valid(fft_mux_0_auto_register_in_w_valid),
    .auto_register_in_w_bits_data(fft_mux_0_auto_register_in_w_bits_data),
    .auto_register_in_w_bits_strb(fft_mux_0_auto_register_in_w_bits_strb),
    .auto_register_in_b_ready(fft_mux_0_auto_register_in_b_ready),
    .auto_register_in_b_valid(fft_mux_0_auto_register_in_b_valid),
    .auto_register_in_b_bits_id(fft_mux_0_auto_register_in_b_bits_id),
    .auto_register_in_ar_ready(fft_mux_0_auto_register_in_ar_ready),
    .auto_register_in_ar_valid(fft_mux_0_auto_register_in_ar_valid),
    .auto_register_in_ar_bits_id(fft_mux_0_auto_register_in_ar_bits_id),
    .auto_register_in_ar_bits_addr(fft_mux_0_auto_register_in_ar_bits_addr),
    .auto_register_in_ar_bits_size(fft_mux_0_auto_register_in_ar_bits_size),
    .auto_register_in_r_ready(fft_mux_0_auto_register_in_r_ready),
    .auto_register_in_r_valid(fft_mux_0_auto_register_in_r_valid),
    .auto_register_in_r_bits_id(fft_mux_0_auto_register_in_r_bits_id),
    .auto_register_in_r_bits_data(fft_mux_0_auto_register_in_r_bits_data),
    .auto_stream_in_2_ready(fft_mux_0_auto_stream_in_2_ready),
    .auto_stream_in_2_valid(fft_mux_0_auto_stream_in_2_valid),
    .auto_stream_in_2_bits_data(fft_mux_0_auto_stream_in_2_bits_data),
    .auto_stream_in_2_bits_last(fft_mux_0_auto_stream_in_2_bits_last),
    .auto_stream_in_1_ready(fft_mux_0_auto_stream_in_1_ready),
    .auto_stream_in_1_valid(fft_mux_0_auto_stream_in_1_valid),
    .auto_stream_in_1_bits_data(fft_mux_0_auto_stream_in_1_bits_data),
    .auto_stream_in_1_bits_last(fft_mux_0_auto_stream_in_1_bits_last),
    .auto_stream_in_0_ready(fft_mux_0_auto_stream_in_0_ready),
    .auto_stream_in_0_valid(fft_mux_0_auto_stream_in_0_valid),
    .auto_stream_in_0_bits_data(fft_mux_0_auto_stream_in_0_bits_data),
    .auto_stream_in_0_bits_last(fft_mux_0_auto_stream_in_0_bits_last),
    .auto_stream_out_0_ready(fft_mux_0_auto_stream_out_0_ready),
    .auto_stream_out_0_valid(fft_mux_0_auto_stream_out_0_valid),
    .auto_stream_out_0_bits_data(fft_mux_0_auto_stream_out_0_bits_data),
    .auto_stream_out_0_bits_last(fft_mux_0_auto_stream_out_0_bits_last)
  );
  AXI4StreamMux_5 fft_mux_1 ( // @[SpectrometerTest.scala 138:29]
    .clock(fft_mux_1_clock),
    .reset(fft_mux_1_reset),
    .auto_register_in_aw_ready(fft_mux_1_auto_register_in_aw_ready),
    .auto_register_in_aw_valid(fft_mux_1_auto_register_in_aw_valid),
    .auto_register_in_aw_bits_id(fft_mux_1_auto_register_in_aw_bits_id),
    .auto_register_in_aw_bits_addr(fft_mux_1_auto_register_in_aw_bits_addr),
    .auto_register_in_w_ready(fft_mux_1_auto_register_in_w_ready),
    .auto_register_in_w_valid(fft_mux_1_auto_register_in_w_valid),
    .auto_register_in_w_bits_data(fft_mux_1_auto_register_in_w_bits_data),
    .auto_register_in_w_bits_strb(fft_mux_1_auto_register_in_w_bits_strb),
    .auto_register_in_b_ready(fft_mux_1_auto_register_in_b_ready),
    .auto_register_in_b_valid(fft_mux_1_auto_register_in_b_valid),
    .auto_register_in_b_bits_id(fft_mux_1_auto_register_in_b_bits_id),
    .auto_register_in_ar_ready(fft_mux_1_auto_register_in_ar_ready),
    .auto_register_in_ar_valid(fft_mux_1_auto_register_in_ar_valid),
    .auto_register_in_ar_bits_id(fft_mux_1_auto_register_in_ar_bits_id),
    .auto_register_in_ar_bits_addr(fft_mux_1_auto_register_in_ar_bits_addr),
    .auto_register_in_ar_bits_size(fft_mux_1_auto_register_in_ar_bits_size),
    .auto_register_in_r_ready(fft_mux_1_auto_register_in_r_ready),
    .auto_register_in_r_valid(fft_mux_1_auto_register_in_r_valid),
    .auto_register_in_r_bits_id(fft_mux_1_auto_register_in_r_bits_id),
    .auto_register_in_r_bits_data(fft_mux_1_auto_register_in_r_bits_data),
    .auto_stream_in_ready(fft_mux_1_auto_stream_in_ready),
    .auto_stream_in_valid(fft_mux_1_auto_stream_in_valid),
    .auto_stream_in_bits_data(fft_mux_1_auto_stream_in_bits_data),
    .auto_stream_in_bits_last(fft_mux_1_auto_stream_in_bits_last),
    .auto_stream_out_1_ready(fft_mux_1_auto_stream_out_1_ready),
    .auto_stream_out_1_valid(fft_mux_1_auto_stream_out_1_valid),
    .auto_stream_out_1_bits_data(fft_mux_1_auto_stream_out_1_bits_data),
    .auto_stream_out_1_bits_last(fft_mux_1_auto_stream_out_1_bits_last)
  );
  AXI4LogMagMuxBlock mag ( // @[SpectrometerTest.scala 144:29]
    .clock(mag_clock),
    .reset(mag_reset),
    .auto_mem_in_aw_ready(mag_auto_mem_in_aw_ready),
    .auto_mem_in_aw_valid(mag_auto_mem_in_aw_valid),
    .auto_mem_in_aw_bits_id(mag_auto_mem_in_aw_bits_id),
    .auto_mem_in_aw_bits_addr(mag_auto_mem_in_aw_bits_addr),
    .auto_mem_in_w_ready(mag_auto_mem_in_w_ready),
    .auto_mem_in_w_valid(mag_auto_mem_in_w_valid),
    .auto_mem_in_w_bits_data(mag_auto_mem_in_w_bits_data),
    .auto_mem_in_w_bits_strb(mag_auto_mem_in_w_bits_strb),
    .auto_mem_in_b_ready(mag_auto_mem_in_b_ready),
    .auto_mem_in_b_valid(mag_auto_mem_in_b_valid),
    .auto_mem_in_b_bits_id(mag_auto_mem_in_b_bits_id),
    .auto_mem_in_ar_ready(mag_auto_mem_in_ar_ready),
    .auto_mem_in_ar_valid(mag_auto_mem_in_ar_valid),
    .auto_mem_in_ar_bits_id(mag_auto_mem_in_ar_bits_id),
    .auto_mem_in_ar_bits_addr(mag_auto_mem_in_ar_bits_addr),
    .auto_mem_in_ar_bits_size(mag_auto_mem_in_ar_bits_size),
    .auto_mem_in_r_ready(mag_auto_mem_in_r_ready),
    .auto_mem_in_r_valid(mag_auto_mem_in_r_valid),
    .auto_mem_in_r_bits_id(mag_auto_mem_in_r_bits_id),
    .auto_mem_in_r_bits_data(mag_auto_mem_in_r_bits_data),
    .auto_stream_in_ready(mag_auto_stream_in_ready),
    .auto_stream_in_valid(mag_auto_stream_in_valid),
    .auto_stream_in_bits_data(mag_auto_stream_in_bits_data),
    .auto_stream_in_bits_last(mag_auto_stream_in_bits_last),
    .auto_stream_out_ready(mag_auto_stream_out_ready),
    .auto_stream_out_valid(mag_auto_stream_out_valid),
    .auto_stream_out_bits_data(mag_auto_stream_out_bits_data),
    .auto_stream_out_bits_last(mag_auto_stream_out_bits_last)
  );
  AXI4Splitter_4 mag_split ( // @[SpectrometerTest.scala 145:29]
    .clock(mag_split_clock),
    .reset(mag_split_reset),
    .auto_mem_in_aw_ready(mag_split_auto_mem_in_aw_ready),
    .auto_mem_in_aw_valid(mag_split_auto_mem_in_aw_valid),
    .auto_mem_in_aw_bits_id(mag_split_auto_mem_in_aw_bits_id),
    .auto_mem_in_aw_bits_addr(mag_split_auto_mem_in_aw_bits_addr),
    .auto_mem_in_w_ready(mag_split_auto_mem_in_w_ready),
    .auto_mem_in_w_valid(mag_split_auto_mem_in_w_valid),
    .auto_mem_in_w_bits_data(mag_split_auto_mem_in_w_bits_data),
    .auto_mem_in_w_bits_strb(mag_split_auto_mem_in_w_bits_strb),
    .auto_mem_in_b_ready(mag_split_auto_mem_in_b_ready),
    .auto_mem_in_b_valid(mag_split_auto_mem_in_b_valid),
    .auto_mem_in_b_bits_id(mag_split_auto_mem_in_b_bits_id),
    .auto_mem_in_ar_ready(mag_split_auto_mem_in_ar_ready),
    .auto_mem_in_ar_valid(mag_split_auto_mem_in_ar_valid),
    .auto_mem_in_ar_bits_id(mag_split_auto_mem_in_ar_bits_id),
    .auto_mem_in_ar_bits_addr(mag_split_auto_mem_in_ar_bits_addr),
    .auto_mem_in_ar_bits_size(mag_split_auto_mem_in_ar_bits_size),
    .auto_mem_in_r_ready(mag_split_auto_mem_in_r_ready),
    .auto_mem_in_r_valid(mag_split_auto_mem_in_r_valid),
    .auto_mem_in_r_bits_id(mag_split_auto_mem_in_r_bits_id),
    .auto_mem_in_r_bits_data(mag_split_auto_mem_in_r_bits_data),
    .auto_stream_in_ready(mag_split_auto_stream_in_ready),
    .auto_stream_in_valid(mag_split_auto_stream_in_valid),
    .auto_stream_in_bits_data(mag_split_auto_stream_in_bits_data),
    .auto_stream_in_bits_last(mag_split_auto_stream_in_bits_last),
    .auto_stream_out_1_ready(mag_split_auto_stream_out_1_ready),
    .auto_stream_out_1_valid(mag_split_auto_stream_out_1_valid),
    .auto_stream_out_1_bits_data(mag_split_auto_stream_out_1_bits_data),
    .auto_stream_out_1_bits_last(mag_split_auto_stream_out_1_bits_last),
    .auto_stream_out_0_ready(mag_split_auto_stream_out_0_ready),
    .auto_stream_out_0_valid(mag_split_auto_stream_out_0_valid),
    .auto_stream_out_0_bits_data(mag_split_auto_stream_out_0_bits_data),
    .auto_stream_out_0_bits_last(mag_split_auto_stream_out_0_bits_last)
  );
  AXI4StreamMux_6 mag_mux_0 ( // @[SpectrometerTest.scala 146:29]
    .clock(mag_mux_0_clock),
    .reset(mag_mux_0_reset),
    .auto_register_in_aw_ready(mag_mux_0_auto_register_in_aw_ready),
    .auto_register_in_aw_valid(mag_mux_0_auto_register_in_aw_valid),
    .auto_register_in_aw_bits_id(mag_mux_0_auto_register_in_aw_bits_id),
    .auto_register_in_aw_bits_addr(mag_mux_0_auto_register_in_aw_bits_addr),
    .auto_register_in_w_ready(mag_mux_0_auto_register_in_w_ready),
    .auto_register_in_w_valid(mag_mux_0_auto_register_in_w_valid),
    .auto_register_in_w_bits_data(mag_mux_0_auto_register_in_w_bits_data),
    .auto_register_in_w_bits_strb(mag_mux_0_auto_register_in_w_bits_strb),
    .auto_register_in_b_ready(mag_mux_0_auto_register_in_b_ready),
    .auto_register_in_b_valid(mag_mux_0_auto_register_in_b_valid),
    .auto_register_in_b_bits_id(mag_mux_0_auto_register_in_b_bits_id),
    .auto_register_in_ar_ready(mag_mux_0_auto_register_in_ar_ready),
    .auto_register_in_ar_valid(mag_mux_0_auto_register_in_ar_valid),
    .auto_register_in_ar_bits_id(mag_mux_0_auto_register_in_ar_bits_id),
    .auto_register_in_ar_bits_addr(mag_mux_0_auto_register_in_ar_bits_addr),
    .auto_register_in_ar_bits_size(mag_mux_0_auto_register_in_ar_bits_size),
    .auto_register_in_r_ready(mag_mux_0_auto_register_in_r_ready),
    .auto_register_in_r_valid(mag_mux_0_auto_register_in_r_valid),
    .auto_register_in_r_bits_id(mag_mux_0_auto_register_in_r_bits_id),
    .auto_register_in_r_bits_data(mag_mux_0_auto_register_in_r_bits_data),
    .auto_stream_in_2_ready(mag_mux_0_auto_stream_in_2_ready),
    .auto_stream_in_2_valid(mag_mux_0_auto_stream_in_2_valid),
    .auto_stream_in_2_bits_data(mag_mux_0_auto_stream_in_2_bits_data),
    .auto_stream_in_2_bits_last(mag_mux_0_auto_stream_in_2_bits_last),
    .auto_stream_in_1_ready(mag_mux_0_auto_stream_in_1_ready),
    .auto_stream_in_1_valid(mag_mux_0_auto_stream_in_1_valid),
    .auto_stream_in_1_bits_data(mag_mux_0_auto_stream_in_1_bits_data),
    .auto_stream_in_1_bits_last(mag_mux_0_auto_stream_in_1_bits_last),
    .auto_stream_in_0_ready(mag_mux_0_auto_stream_in_0_ready),
    .auto_stream_in_0_valid(mag_mux_0_auto_stream_in_0_valid),
    .auto_stream_in_0_bits_data(mag_mux_0_auto_stream_in_0_bits_data),
    .auto_stream_in_0_bits_last(mag_mux_0_auto_stream_in_0_bits_last),
    .auto_stream_out_0_ready(mag_mux_0_auto_stream_out_0_ready),
    .auto_stream_out_0_valid(mag_mux_0_auto_stream_out_0_valid),
    .auto_stream_out_0_bits_data(mag_mux_0_auto_stream_out_0_bits_data),
    .auto_stream_out_0_bits_last(mag_mux_0_auto_stream_out_0_bits_last)
  );
  AXI4StreamMux_7 mag_mux_1 ( // @[SpectrometerTest.scala 147:29]
    .clock(mag_mux_1_clock),
    .reset(mag_mux_1_reset),
    .auto_register_in_aw_ready(mag_mux_1_auto_register_in_aw_ready),
    .auto_register_in_aw_valid(mag_mux_1_auto_register_in_aw_valid),
    .auto_register_in_aw_bits_id(mag_mux_1_auto_register_in_aw_bits_id),
    .auto_register_in_aw_bits_addr(mag_mux_1_auto_register_in_aw_bits_addr),
    .auto_register_in_w_ready(mag_mux_1_auto_register_in_w_ready),
    .auto_register_in_w_valid(mag_mux_1_auto_register_in_w_valid),
    .auto_register_in_w_bits_data(mag_mux_1_auto_register_in_w_bits_data),
    .auto_register_in_w_bits_strb(mag_mux_1_auto_register_in_w_bits_strb),
    .auto_register_in_b_ready(mag_mux_1_auto_register_in_b_ready),
    .auto_register_in_b_valid(mag_mux_1_auto_register_in_b_valid),
    .auto_register_in_b_bits_id(mag_mux_1_auto_register_in_b_bits_id),
    .auto_register_in_ar_ready(mag_mux_1_auto_register_in_ar_ready),
    .auto_register_in_ar_valid(mag_mux_1_auto_register_in_ar_valid),
    .auto_register_in_ar_bits_id(mag_mux_1_auto_register_in_ar_bits_id),
    .auto_register_in_ar_bits_addr(mag_mux_1_auto_register_in_ar_bits_addr),
    .auto_register_in_ar_bits_size(mag_mux_1_auto_register_in_ar_bits_size),
    .auto_register_in_r_ready(mag_mux_1_auto_register_in_r_ready),
    .auto_register_in_r_valid(mag_mux_1_auto_register_in_r_valid),
    .auto_register_in_r_bits_id(mag_mux_1_auto_register_in_r_bits_id),
    .auto_register_in_r_bits_data(mag_mux_1_auto_register_in_r_bits_data),
    .auto_stream_in_ready(mag_mux_1_auto_stream_in_ready),
    .auto_stream_in_valid(mag_mux_1_auto_stream_in_valid),
    .auto_stream_in_bits_data(mag_mux_1_auto_stream_in_bits_data),
    .auto_stream_in_bits_last(mag_mux_1_auto_stream_in_bits_last),
    .auto_stream_out_1_ready(mag_mux_1_auto_stream_out_1_ready),
    .auto_stream_out_1_valid(mag_mux_1_auto_stream_out_1_valid),
    .auto_stream_out_1_bits_data(mag_mux_1_auto_stream_out_1_bits_data),
    .auto_stream_out_1_bits_last(mag_mux_1_auto_stream_out_1_bits_last)
  );
  AccumulatorChain acc ( // @[SpectrometerTest.scala 153:29]
    .clock(acc_clock),
    .reset(acc_reset),
    .auto_bus_in_aw_ready(acc_auto_bus_in_aw_ready),
    .auto_bus_in_aw_valid(acc_auto_bus_in_aw_valid),
    .auto_bus_in_aw_bits_id(acc_auto_bus_in_aw_bits_id),
    .auto_bus_in_aw_bits_addr(acc_auto_bus_in_aw_bits_addr),
    .auto_bus_in_aw_bits_size(acc_auto_bus_in_aw_bits_size),
    .auto_bus_in_w_ready(acc_auto_bus_in_w_ready),
    .auto_bus_in_w_valid(acc_auto_bus_in_w_valid),
    .auto_bus_in_w_bits_data(acc_auto_bus_in_w_bits_data),
    .auto_bus_in_w_bits_strb(acc_auto_bus_in_w_bits_strb),
    .auto_bus_in_w_bits_last(acc_auto_bus_in_w_bits_last),
    .auto_bus_in_b_ready(acc_auto_bus_in_b_ready),
    .auto_bus_in_b_valid(acc_auto_bus_in_b_valid),
    .auto_bus_in_b_bits_resp(acc_auto_bus_in_b_bits_resp),
    .auto_bus_in_ar_ready(acc_auto_bus_in_ar_ready),
    .auto_bus_in_ar_valid(acc_auto_bus_in_ar_valid),
    .auto_bus_in_ar_bits_id(acc_auto_bus_in_ar_bits_id),
    .auto_bus_in_ar_bits_addr(acc_auto_bus_in_ar_bits_addr),
    .auto_bus_in_ar_bits_size(acc_auto_bus_in_ar_bits_size),
    .auto_bus_in_r_ready(acc_auto_bus_in_r_ready),
    .auto_bus_in_r_valid(acc_auto_bus_in_r_valid),
    .auto_bus_in_r_bits_data(acc_auto_bus_in_r_bits_data),
    .auto_bus_in_r_bits_resp(acc_auto_bus_in_r_bits_resp),
    .auto_bus_in_r_bits_last(acc_auto_bus_in_r_bits_last),
    .auto_dspQueue_stream_out_ready(acc_auto_dspQueue_stream_out_ready),
    .auto_dspQueue_stream_out_valid(acc_auto_dspQueue_stream_out_valid),
    .auto_dspQueue_stream_out_bits_data(acc_auto_dspQueue_stream_out_bits_data),
    .auto_dspQueue_stream_out_bits_last(acc_auto_dspQueue_stream_out_bits_last),
    .auto_accumulator_slave_in_ready(acc_auto_accumulator_slave_in_ready),
    .auto_accumulator_slave_in_valid(acc_auto_accumulator_slave_in_valid),
    .auto_accumulator_slave_in_bits_data(acc_auto_accumulator_slave_in_bits_data),
    .auto_accumulator_slave_in_bits_last(acc_auto_accumulator_slave_in_bits_last)
  );
  AXI4StreamWidthAdapater_2_to_1 widthAdapter_1 ( // @[AXI4StreamWidthAdapter.scala 82:34]
    .clock(widthAdapter_1_clock),
    .reset(widthAdapter_1_reset),
    .auto_in_ready(widthAdapter_1_auto_in_ready),
    .auto_in_valid(widthAdapter_1_auto_in_valid),
    .auto_in_bits_data(widthAdapter_1_auto_in_bits_data),
    .auto_in_bits_last(widthAdapter_1_auto_in_bits_last),
    .auto_out_ready(widthAdapter_1_auto_out_ready),
    .auto_out_valid(widthAdapter_1_auto_out_valid),
    .auto_out_bits_data(widthAdapter_1_auto_out_bits_data),
    .auto_out_bits_last(widthAdapter_1_auto_out_bits_last)
  );
  StreamBuffer_1 acc_queue ( // @[SpectrometerTest.scala 155:29]
    .clock(acc_queue_clock),
    .reset(acc_queue_reset),
    .auto_out_out_ready(acc_queue_auto_out_out_ready),
    .auto_out_out_valid(acc_queue_auto_out_out_valid),
    .auto_out_out_bits_data(acc_queue_auto_out_out_bits_data),
    .auto_out_out_bits_last(acc_queue_auto_out_out_bits_last),
    .auto_in_in_ready(acc_queue_auto_in_in_ready),
    .auto_in_in_valid(acc_queue_auto_in_in_valid),
    .auto_in_in_bits_data(acc_queue_auto_in_in_bits_data),
    .auto_in_in_bits_last(acc_queue_auto_in_in_bits_last)
  );
  AXI4StreamMux_8 out_mux ( // @[SpectrometerTest.scala 157:29]
    .clock(out_mux_clock),
    .reset(out_mux_reset),
    .auto_register_in_aw_ready(out_mux_auto_register_in_aw_ready),
    .auto_register_in_aw_valid(out_mux_auto_register_in_aw_valid),
    .auto_register_in_aw_bits_id(out_mux_auto_register_in_aw_bits_id),
    .auto_register_in_aw_bits_addr(out_mux_auto_register_in_aw_bits_addr),
    .auto_register_in_w_ready(out_mux_auto_register_in_w_ready),
    .auto_register_in_w_valid(out_mux_auto_register_in_w_valid),
    .auto_register_in_w_bits_data(out_mux_auto_register_in_w_bits_data),
    .auto_register_in_w_bits_strb(out_mux_auto_register_in_w_bits_strb),
    .auto_register_in_b_ready(out_mux_auto_register_in_b_ready),
    .auto_register_in_b_valid(out_mux_auto_register_in_b_valid),
    .auto_register_in_b_bits_id(out_mux_auto_register_in_b_bits_id),
    .auto_register_in_ar_ready(out_mux_auto_register_in_ar_ready),
    .auto_register_in_ar_valid(out_mux_auto_register_in_ar_valid),
    .auto_register_in_ar_bits_id(out_mux_auto_register_in_ar_bits_id),
    .auto_register_in_ar_bits_addr(out_mux_auto_register_in_ar_bits_addr),
    .auto_register_in_ar_bits_size(out_mux_auto_register_in_ar_bits_size),
    .auto_register_in_r_ready(out_mux_auto_register_in_r_ready),
    .auto_register_in_r_valid(out_mux_auto_register_in_r_valid),
    .auto_register_in_r_bits_id(out_mux_auto_register_in_r_bits_id),
    .auto_register_in_r_bits_data(out_mux_auto_register_in_r_bits_data),
    .auto_stream_in_6_ready(out_mux_auto_stream_in_6_ready),
    .auto_stream_in_6_valid(out_mux_auto_stream_in_6_valid),
    .auto_stream_in_6_bits_data(out_mux_auto_stream_in_6_bits_data),
    .auto_stream_in_6_bits_last(out_mux_auto_stream_in_6_bits_last),
    .auto_stream_in_5_ready(out_mux_auto_stream_in_5_ready),
    .auto_stream_in_5_valid(out_mux_auto_stream_in_5_valid),
    .auto_stream_in_5_bits_data(out_mux_auto_stream_in_5_bits_data),
    .auto_stream_in_5_bits_last(out_mux_auto_stream_in_5_bits_last),
    .auto_stream_in_4_ready(out_mux_auto_stream_in_4_ready),
    .auto_stream_in_4_valid(out_mux_auto_stream_in_4_valid),
    .auto_stream_in_4_bits_data(out_mux_auto_stream_in_4_bits_data),
    .auto_stream_in_4_bits_last(out_mux_auto_stream_in_4_bits_last),
    .auto_stream_in_3_ready(out_mux_auto_stream_in_3_ready),
    .auto_stream_in_3_valid(out_mux_auto_stream_in_3_valid),
    .auto_stream_in_3_bits_data(out_mux_auto_stream_in_3_bits_data),
    .auto_stream_in_3_bits_last(out_mux_auto_stream_in_3_bits_last),
    .auto_stream_in_2_ready(out_mux_auto_stream_in_2_ready),
    .auto_stream_in_2_valid(out_mux_auto_stream_in_2_valid),
    .auto_stream_in_2_bits_data(out_mux_auto_stream_in_2_bits_data),
    .auto_stream_in_2_bits_last(out_mux_auto_stream_in_2_bits_last),
    .auto_stream_in_1_ready(out_mux_auto_stream_in_1_ready),
    .auto_stream_in_1_valid(out_mux_auto_stream_in_1_valid),
    .auto_stream_in_1_bits_data(out_mux_auto_stream_in_1_bits_data),
    .auto_stream_in_1_bits_last(out_mux_auto_stream_in_1_bits_last),
    .auto_stream_in_0_ready(out_mux_auto_stream_in_0_ready),
    .auto_stream_in_0_valid(out_mux_auto_stream_in_0_valid),
    .auto_stream_in_0_bits_data(out_mux_auto_stream_in_0_bits_data),
    .auto_stream_in_0_bits_last(out_mux_auto_stream_in_0_bits_last),
    .auto_stream_out_1_ready(out_mux_auto_stream_out_1_ready),
    .auto_stream_out_1_valid(out_mux_auto_stream_out_1_valid),
    .auto_stream_out_1_bits_data(out_mux_auto_stream_out_1_bits_data),
    .auto_stream_out_1_bits_last(out_mux_auto_stream_out_1_bits_last),
    .auto_stream_out_0_ready(out_mux_auto_stream_out_0_ready),
    .auto_stream_out_0_valid(out_mux_auto_stream_out_0_valid),
    .auto_stream_out_0_bits_data(out_mux_auto_stream_out_0_bits_data),
    .auto_stream_out_0_bits_last(out_mux_auto_stream_out_0_bits_last)
  );
  StreamBuffer_2 out_queue ( // @[SpectrometerTest.scala 158:29]
    .clock(out_queue_clock),
    .reset(out_queue_reset),
    .auto_out_out_ready(out_queue_auto_out_out_ready),
    .auto_out_out_valid(out_queue_auto_out_out_valid),
    .auto_out_out_bits_data(out_queue_auto_out_out_bits_data),
    .auto_out_out_bits_last(out_queue_auto_out_out_bits_last),
    .auto_in_in_ready(out_queue_auto_in_in_ready),
    .auto_in_in_valid(out_queue_auto_in_in_valid),
    .auto_in_in_bits_data(out_queue_auto_in_in_bits_data),
    .auto_in_in_bits_last(out_queue_auto_in_in_bits_last)
  );
  AXI4StreamWidthAdapater_1_to_4 widthAdapter_2 ( // @[AXI4StreamWidthAdapter.scala 82:34]
    .clock(widthAdapter_2_clock),
    .reset(widthAdapter_2_reset),
    .auto_in_ready(widthAdapter_2_auto_in_ready),
    .auto_in_valid(widthAdapter_2_auto_in_valid),
    .auto_in_bits_data(widthAdapter_2_auto_in_bits_data),
    .auto_in_bits_last(widthAdapter_2_auto_in_bits_last),
    .auto_out_ready(widthAdapter_2_auto_out_ready),
    .auto_out_valid(widthAdapter_2_auto_out_valid),
    .auto_out_bits_data(widthAdapter_2_auto_out_bits_data),
    .auto_out_bits_last(widthAdapter_2_auto_out_bits_last)
  );
  StreamBuffer_3 uTx_queue ( // @[SpectrometerTest.scala 162:29]
    .clock(uTx_queue_clock),
    .reset(uTx_queue_reset),
    .auto_out_out_ready(uTx_queue_auto_out_out_ready),
    .auto_out_out_valid(uTx_queue_auto_out_out_valid),
    .auto_out_out_bits_data(uTx_queue_auto_out_out_bits_data),
    .auto_out_out_bits_last(uTx_queue_auto_out_out_bits_last),
    .auto_in_in_ready(uTx_queue_auto_in_in_ready),
    .auto_in_in_valid(uTx_queue_auto_in_in_valid),
    .auto_in_in_bits_data(uTx_queue_auto_in_in_bits_data),
    .auto_in_in_bits_last(uTx_queue_auto_in_in_bits_last)
  );
  AXI4StreamWidthAdapater_1_to_4 widthAdapter_3 ( // @[AXI4StreamWidthAdapter.scala 82:34]
    .clock(widthAdapter_3_clock),
    .reset(widthAdapter_3_reset),
    .auto_in_ready(widthAdapter_3_auto_in_ready),
    .auto_in_valid(widthAdapter_3_auto_in_valid),
    .auto_in_bits_data(widthAdapter_3_auto_in_bits_data),
    .auto_in_bits_last(widthAdapter_3_auto_in_bits_last),
    .auto_out_ready(widthAdapter_3_auto_out_ready),
    .auto_out_valid(widthAdapter_3_auto_out_valid),
    .auto_out_bits_data(widthAdapter_3_auto_out_bits_data),
    .auto_out_bits_last(widthAdapter_3_auto_out_bits_last)
  );
  AXI4StreamWidthAdapater_4_to_1 widthAdapter_4 ( // @[AXI4StreamWidthAdapter.scala 82:34]
    .clock(widthAdapter_4_clock),
    .reset(widthAdapter_4_reset),
    .auto_in_ready(widthAdapter_4_auto_in_ready),
    .auto_in_valid(widthAdapter_4_auto_in_valid),
    .auto_in_bits_data(widthAdapter_4_auto_in_bits_data),
    .auto_in_bits_last(widthAdapter_4_auto_in_bits_last),
    .auto_out_ready(widthAdapter_4_auto_out_ready),
    .auto_out_valid(widthAdapter_4_auto_out_valid),
    .auto_out_bits_data(widthAdapter_4_auto_out_bits_data),
    .auto_out_bits_last(widthAdapter_4_auto_out_bits_last)
  );
  AXI4Splitter uRx_split ( // @[SpectrometerTest.scala 165:29]
    .clock(uRx_split_clock),
    .reset(uRx_split_reset),
    .auto_mem_in_aw_ready(uRx_split_auto_mem_in_aw_ready),
    .auto_mem_in_aw_valid(uRx_split_auto_mem_in_aw_valid),
    .auto_mem_in_aw_bits_id(uRx_split_auto_mem_in_aw_bits_id),
    .auto_mem_in_aw_bits_addr(uRx_split_auto_mem_in_aw_bits_addr),
    .auto_mem_in_w_ready(uRx_split_auto_mem_in_w_ready),
    .auto_mem_in_w_valid(uRx_split_auto_mem_in_w_valid),
    .auto_mem_in_w_bits_data(uRx_split_auto_mem_in_w_bits_data),
    .auto_mem_in_w_bits_strb(uRx_split_auto_mem_in_w_bits_strb),
    .auto_mem_in_b_ready(uRx_split_auto_mem_in_b_ready),
    .auto_mem_in_b_valid(uRx_split_auto_mem_in_b_valid),
    .auto_mem_in_b_bits_id(uRx_split_auto_mem_in_b_bits_id),
    .auto_mem_in_ar_ready(uRx_split_auto_mem_in_ar_ready),
    .auto_mem_in_ar_valid(uRx_split_auto_mem_in_ar_valid),
    .auto_mem_in_ar_bits_id(uRx_split_auto_mem_in_ar_bits_id),
    .auto_mem_in_ar_bits_addr(uRx_split_auto_mem_in_ar_bits_addr),
    .auto_mem_in_ar_bits_size(uRx_split_auto_mem_in_ar_bits_size),
    .auto_mem_in_r_ready(uRx_split_auto_mem_in_r_ready),
    .auto_mem_in_r_valid(uRx_split_auto_mem_in_r_valid),
    .auto_mem_in_r_bits_id(uRx_split_auto_mem_in_r_bits_id),
    .auto_mem_in_r_bits_data(uRx_split_auto_mem_in_r_bits_data),
    .auto_stream_in_ready(uRx_split_auto_stream_in_ready),
    .auto_stream_in_valid(uRx_split_auto_stream_in_valid),
    .auto_stream_in_bits_data(uRx_split_auto_stream_in_bits_data),
    .auto_stream_in_bits_last(uRx_split_auto_stream_in_bits_last),
    .auto_stream_out_4_ready(uRx_split_auto_stream_out_4_ready),
    .auto_stream_out_4_valid(uRx_split_auto_stream_out_4_valid),
    .auto_stream_out_4_bits_data(uRx_split_auto_stream_out_4_bits_data),
    .auto_stream_out_4_bits_last(uRx_split_auto_stream_out_4_bits_last),
    .auto_stream_out_3_ready(uRx_split_auto_stream_out_3_ready),
    .auto_stream_out_3_valid(uRx_split_auto_stream_out_3_valid),
    .auto_stream_out_3_bits_data(uRx_split_auto_stream_out_3_bits_data),
    .auto_stream_out_3_bits_last(uRx_split_auto_stream_out_3_bits_last),
    .auto_stream_out_2_ready(uRx_split_auto_stream_out_2_ready),
    .auto_stream_out_2_valid(uRx_split_auto_stream_out_2_valid),
    .auto_stream_out_2_bits_data(uRx_split_auto_stream_out_2_bits_data),
    .auto_stream_out_2_bits_last(uRx_split_auto_stream_out_2_bits_last),
    .auto_stream_out_1_ready(uRx_split_auto_stream_out_1_ready),
    .auto_stream_out_1_valid(uRx_split_auto_stream_out_1_valid),
    .auto_stream_out_1_bits_data(uRx_split_auto_stream_out_1_bits_data),
    .auto_stream_out_1_bits_last(uRx_split_auto_stream_out_1_bits_last),
    .auto_stream_out_0_ready(uRx_split_auto_stream_out_0_ready),
    .auto_stream_out_0_valid(uRx_split_auto_stream_out_0_valid),
    .auto_stream_out_0_bits_data(uRx_split_auto_stream_out_0_bits_data),
    .auto_stream_out_0_bits_last(uRx_split_auto_stream_out_0_bits_last)
  );
  AXI4UARTBlock uart ( // @[SpectrometerTest.scala 166:29]
    .clock(uart_clock),
    .reset(uart_reset),
    .auto_mem_in_aw_ready(uart_auto_mem_in_aw_ready),
    .auto_mem_in_aw_valid(uart_auto_mem_in_aw_valid),
    .auto_mem_in_aw_bits_id(uart_auto_mem_in_aw_bits_id),
    .auto_mem_in_aw_bits_addr(uart_auto_mem_in_aw_bits_addr),
    .auto_mem_in_w_ready(uart_auto_mem_in_w_ready),
    .auto_mem_in_w_valid(uart_auto_mem_in_w_valid),
    .auto_mem_in_w_bits_data(uart_auto_mem_in_w_bits_data),
    .auto_mem_in_w_bits_strb(uart_auto_mem_in_w_bits_strb),
    .auto_mem_in_b_ready(uart_auto_mem_in_b_ready),
    .auto_mem_in_b_valid(uart_auto_mem_in_b_valid),
    .auto_mem_in_b_bits_id(uart_auto_mem_in_b_bits_id),
    .auto_mem_in_ar_ready(uart_auto_mem_in_ar_ready),
    .auto_mem_in_ar_valid(uart_auto_mem_in_ar_valid),
    .auto_mem_in_ar_bits_id(uart_auto_mem_in_ar_bits_id),
    .auto_mem_in_ar_bits_addr(uart_auto_mem_in_ar_bits_addr),
    .auto_mem_in_ar_bits_size(uart_auto_mem_in_ar_bits_size),
    .auto_mem_in_r_ready(uart_auto_mem_in_r_ready),
    .auto_mem_in_r_valid(uart_auto_mem_in_r_valid),
    .auto_mem_in_r_bits_id(uart_auto_mem_in_r_bits_id),
    .auto_mem_in_r_bits_data(uart_auto_mem_in_r_bits_data),
    .auto_in_in_ready(uart_auto_in_in_ready),
    .auto_in_in_valid(uart_auto_in_in_valid),
    .auto_in_in_bits_data(uart_auto_in_in_bits_data),
    .auto_out_out_ready(uart_auto_out_out_ready),
    .auto_out_out_valid(uart_auto_out_out_valid),
    .auto_out_out_bits_data(uart_auto_out_out_bits_data),
    .int_0(uart_int_0),
    .io_txd(uart_io_txd),
    .io_rxd(uart_io_rxd)
  );
  AXI4Xbar_2 bus ( // @[SpectrometerTest.scala 180:23]
    .clock(bus_clock),
    .reset(bus_reset),
    .auto_in_aw_ready(bus_auto_in_aw_ready),
    .auto_in_aw_valid(bus_auto_in_aw_valid),
    .auto_in_aw_bits_id(bus_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(bus_auto_in_aw_bits_addr),
    .auto_in_aw_bits_size(bus_auto_in_aw_bits_size),
    .auto_in_w_ready(bus_auto_in_w_ready),
    .auto_in_w_valid(bus_auto_in_w_valid),
    .auto_in_w_bits_data(bus_auto_in_w_bits_data),
    .auto_in_w_bits_strb(bus_auto_in_w_bits_strb),
    .auto_in_w_bits_last(bus_auto_in_w_bits_last),
    .auto_in_b_ready(bus_auto_in_b_ready),
    .auto_in_b_valid(bus_auto_in_b_valid),
    .auto_in_b_bits_resp(bus_auto_in_b_bits_resp),
    .auto_in_ar_ready(bus_auto_in_ar_ready),
    .auto_in_ar_valid(bus_auto_in_ar_valid),
    .auto_in_ar_bits_id(bus_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(bus_auto_in_ar_bits_addr),
    .auto_in_ar_bits_size(bus_auto_in_ar_bits_size),
    .auto_in_r_ready(bus_auto_in_r_ready),
    .auto_in_r_valid(bus_auto_in_r_valid),
    .auto_in_r_bits_data(bus_auto_in_r_bits_data),
    .auto_in_r_bits_resp(bus_auto_in_r_bits_resp),
    .auto_in_r_bits_last(bus_auto_in_r_bits_last),
    .auto_out_20_aw_ready(bus_auto_out_20_aw_ready),
    .auto_out_20_aw_valid(bus_auto_out_20_aw_valid),
    .auto_out_20_aw_bits_id(bus_auto_out_20_aw_bits_id),
    .auto_out_20_aw_bits_addr(bus_auto_out_20_aw_bits_addr),
    .auto_out_20_aw_bits_size(bus_auto_out_20_aw_bits_size),
    .auto_out_20_w_ready(bus_auto_out_20_w_ready),
    .auto_out_20_w_valid(bus_auto_out_20_w_valid),
    .auto_out_20_w_bits_data(bus_auto_out_20_w_bits_data),
    .auto_out_20_w_bits_strb(bus_auto_out_20_w_bits_strb),
    .auto_out_20_w_bits_last(bus_auto_out_20_w_bits_last),
    .auto_out_20_b_ready(bus_auto_out_20_b_ready),
    .auto_out_20_b_valid(bus_auto_out_20_b_valid),
    .auto_out_20_b_bits_resp(bus_auto_out_20_b_bits_resp),
    .auto_out_20_ar_ready(bus_auto_out_20_ar_ready),
    .auto_out_20_ar_valid(bus_auto_out_20_ar_valid),
    .auto_out_20_ar_bits_id(bus_auto_out_20_ar_bits_id),
    .auto_out_20_ar_bits_addr(bus_auto_out_20_ar_bits_addr),
    .auto_out_20_ar_bits_size(bus_auto_out_20_ar_bits_size),
    .auto_out_20_r_ready(bus_auto_out_20_r_ready),
    .auto_out_20_r_valid(bus_auto_out_20_r_valid),
    .auto_out_20_r_bits_data(bus_auto_out_20_r_bits_data),
    .auto_out_20_r_bits_resp(bus_auto_out_20_r_bits_resp),
    .auto_out_20_r_bits_last(bus_auto_out_20_r_bits_last),
    .auto_out_19_aw_ready(bus_auto_out_19_aw_ready),
    .auto_out_19_aw_valid(bus_auto_out_19_aw_valid),
    .auto_out_19_aw_bits_id(bus_auto_out_19_aw_bits_id),
    .auto_out_19_aw_bits_addr(bus_auto_out_19_aw_bits_addr),
    .auto_out_19_aw_bits_size(bus_auto_out_19_aw_bits_size),
    .auto_out_19_w_ready(bus_auto_out_19_w_ready),
    .auto_out_19_w_valid(bus_auto_out_19_w_valid),
    .auto_out_19_w_bits_data(bus_auto_out_19_w_bits_data),
    .auto_out_19_w_bits_strb(bus_auto_out_19_w_bits_strb),
    .auto_out_19_w_bits_last(bus_auto_out_19_w_bits_last),
    .auto_out_19_b_ready(bus_auto_out_19_b_ready),
    .auto_out_19_b_valid(bus_auto_out_19_b_valid),
    .auto_out_19_b_bits_id(bus_auto_out_19_b_bits_id),
    .auto_out_19_b_bits_resp(bus_auto_out_19_b_bits_resp),
    .auto_out_19_ar_ready(bus_auto_out_19_ar_ready),
    .auto_out_19_ar_valid(bus_auto_out_19_ar_valid),
    .auto_out_19_ar_bits_id(bus_auto_out_19_ar_bits_id),
    .auto_out_19_ar_bits_addr(bus_auto_out_19_ar_bits_addr),
    .auto_out_19_ar_bits_size(bus_auto_out_19_ar_bits_size),
    .auto_out_19_r_ready(bus_auto_out_19_r_ready),
    .auto_out_19_r_valid(bus_auto_out_19_r_valid),
    .auto_out_19_r_bits_id(bus_auto_out_19_r_bits_id),
    .auto_out_19_r_bits_data(bus_auto_out_19_r_bits_data),
    .auto_out_19_r_bits_resp(bus_auto_out_19_r_bits_resp),
    .auto_out_19_r_bits_last(bus_auto_out_19_r_bits_last),
    .auto_out_18_aw_ready(bus_auto_out_18_aw_ready),
    .auto_out_18_aw_valid(bus_auto_out_18_aw_valid),
    .auto_out_18_aw_bits_id(bus_auto_out_18_aw_bits_id),
    .auto_out_18_aw_bits_addr(bus_auto_out_18_aw_bits_addr),
    .auto_out_18_aw_bits_size(bus_auto_out_18_aw_bits_size),
    .auto_out_18_w_ready(bus_auto_out_18_w_ready),
    .auto_out_18_w_valid(bus_auto_out_18_w_valid),
    .auto_out_18_w_bits_data(bus_auto_out_18_w_bits_data),
    .auto_out_18_w_bits_strb(bus_auto_out_18_w_bits_strb),
    .auto_out_18_w_bits_last(bus_auto_out_18_w_bits_last),
    .auto_out_18_b_ready(bus_auto_out_18_b_ready),
    .auto_out_18_b_valid(bus_auto_out_18_b_valid),
    .auto_out_18_b_bits_id(bus_auto_out_18_b_bits_id),
    .auto_out_18_b_bits_resp(bus_auto_out_18_b_bits_resp),
    .auto_out_18_ar_ready(bus_auto_out_18_ar_ready),
    .auto_out_18_ar_valid(bus_auto_out_18_ar_valid),
    .auto_out_18_ar_bits_id(bus_auto_out_18_ar_bits_id),
    .auto_out_18_ar_bits_addr(bus_auto_out_18_ar_bits_addr),
    .auto_out_18_ar_bits_size(bus_auto_out_18_ar_bits_size),
    .auto_out_18_r_ready(bus_auto_out_18_r_ready),
    .auto_out_18_r_valid(bus_auto_out_18_r_valid),
    .auto_out_18_r_bits_id(bus_auto_out_18_r_bits_id),
    .auto_out_18_r_bits_data(bus_auto_out_18_r_bits_data),
    .auto_out_18_r_bits_resp(bus_auto_out_18_r_bits_resp),
    .auto_out_18_r_bits_last(bus_auto_out_18_r_bits_last),
    .auto_out_17_aw_ready(bus_auto_out_17_aw_ready),
    .auto_out_17_aw_valid(bus_auto_out_17_aw_valid),
    .auto_out_17_aw_bits_id(bus_auto_out_17_aw_bits_id),
    .auto_out_17_aw_bits_addr(bus_auto_out_17_aw_bits_addr),
    .auto_out_17_aw_bits_size(bus_auto_out_17_aw_bits_size),
    .auto_out_17_w_ready(bus_auto_out_17_w_ready),
    .auto_out_17_w_valid(bus_auto_out_17_w_valid),
    .auto_out_17_w_bits_data(bus_auto_out_17_w_bits_data),
    .auto_out_17_w_bits_strb(bus_auto_out_17_w_bits_strb),
    .auto_out_17_w_bits_last(bus_auto_out_17_w_bits_last),
    .auto_out_17_b_ready(bus_auto_out_17_b_ready),
    .auto_out_17_b_valid(bus_auto_out_17_b_valid),
    .auto_out_17_b_bits_id(bus_auto_out_17_b_bits_id),
    .auto_out_17_b_bits_resp(bus_auto_out_17_b_bits_resp),
    .auto_out_17_ar_ready(bus_auto_out_17_ar_ready),
    .auto_out_17_ar_valid(bus_auto_out_17_ar_valid),
    .auto_out_17_ar_bits_id(bus_auto_out_17_ar_bits_id),
    .auto_out_17_ar_bits_addr(bus_auto_out_17_ar_bits_addr),
    .auto_out_17_ar_bits_size(bus_auto_out_17_ar_bits_size),
    .auto_out_17_r_ready(bus_auto_out_17_r_ready),
    .auto_out_17_r_valid(bus_auto_out_17_r_valid),
    .auto_out_17_r_bits_id(bus_auto_out_17_r_bits_id),
    .auto_out_17_r_bits_data(bus_auto_out_17_r_bits_data),
    .auto_out_17_r_bits_resp(bus_auto_out_17_r_bits_resp),
    .auto_out_17_r_bits_last(bus_auto_out_17_r_bits_last),
    .auto_out_16_aw_ready(bus_auto_out_16_aw_ready),
    .auto_out_16_aw_valid(bus_auto_out_16_aw_valid),
    .auto_out_16_aw_bits_id(bus_auto_out_16_aw_bits_id),
    .auto_out_16_aw_bits_addr(bus_auto_out_16_aw_bits_addr),
    .auto_out_16_aw_bits_size(bus_auto_out_16_aw_bits_size),
    .auto_out_16_w_ready(bus_auto_out_16_w_ready),
    .auto_out_16_w_valid(bus_auto_out_16_w_valid),
    .auto_out_16_w_bits_data(bus_auto_out_16_w_bits_data),
    .auto_out_16_w_bits_strb(bus_auto_out_16_w_bits_strb),
    .auto_out_16_w_bits_last(bus_auto_out_16_w_bits_last),
    .auto_out_16_b_ready(bus_auto_out_16_b_ready),
    .auto_out_16_b_valid(bus_auto_out_16_b_valid),
    .auto_out_16_b_bits_id(bus_auto_out_16_b_bits_id),
    .auto_out_16_b_bits_resp(bus_auto_out_16_b_bits_resp),
    .auto_out_16_ar_ready(bus_auto_out_16_ar_ready),
    .auto_out_16_ar_valid(bus_auto_out_16_ar_valid),
    .auto_out_16_ar_bits_id(bus_auto_out_16_ar_bits_id),
    .auto_out_16_ar_bits_addr(bus_auto_out_16_ar_bits_addr),
    .auto_out_16_ar_bits_size(bus_auto_out_16_ar_bits_size),
    .auto_out_16_r_ready(bus_auto_out_16_r_ready),
    .auto_out_16_r_valid(bus_auto_out_16_r_valid),
    .auto_out_16_r_bits_id(bus_auto_out_16_r_bits_id),
    .auto_out_16_r_bits_data(bus_auto_out_16_r_bits_data),
    .auto_out_16_r_bits_resp(bus_auto_out_16_r_bits_resp),
    .auto_out_16_r_bits_last(bus_auto_out_16_r_bits_last),
    .auto_out_15_aw_ready(bus_auto_out_15_aw_ready),
    .auto_out_15_aw_valid(bus_auto_out_15_aw_valid),
    .auto_out_15_aw_bits_id(bus_auto_out_15_aw_bits_id),
    .auto_out_15_aw_bits_addr(bus_auto_out_15_aw_bits_addr),
    .auto_out_15_aw_bits_size(bus_auto_out_15_aw_bits_size),
    .auto_out_15_w_ready(bus_auto_out_15_w_ready),
    .auto_out_15_w_valid(bus_auto_out_15_w_valid),
    .auto_out_15_w_bits_data(bus_auto_out_15_w_bits_data),
    .auto_out_15_w_bits_strb(bus_auto_out_15_w_bits_strb),
    .auto_out_15_w_bits_last(bus_auto_out_15_w_bits_last),
    .auto_out_15_b_ready(bus_auto_out_15_b_ready),
    .auto_out_15_b_valid(bus_auto_out_15_b_valid),
    .auto_out_15_b_bits_id(bus_auto_out_15_b_bits_id),
    .auto_out_15_b_bits_resp(bus_auto_out_15_b_bits_resp),
    .auto_out_15_ar_ready(bus_auto_out_15_ar_ready),
    .auto_out_15_ar_valid(bus_auto_out_15_ar_valid),
    .auto_out_15_ar_bits_id(bus_auto_out_15_ar_bits_id),
    .auto_out_15_ar_bits_addr(bus_auto_out_15_ar_bits_addr),
    .auto_out_15_ar_bits_size(bus_auto_out_15_ar_bits_size),
    .auto_out_15_r_ready(bus_auto_out_15_r_ready),
    .auto_out_15_r_valid(bus_auto_out_15_r_valid),
    .auto_out_15_r_bits_id(bus_auto_out_15_r_bits_id),
    .auto_out_15_r_bits_data(bus_auto_out_15_r_bits_data),
    .auto_out_15_r_bits_resp(bus_auto_out_15_r_bits_resp),
    .auto_out_15_r_bits_last(bus_auto_out_15_r_bits_last),
    .auto_out_14_aw_ready(bus_auto_out_14_aw_ready),
    .auto_out_14_aw_valid(bus_auto_out_14_aw_valid),
    .auto_out_14_aw_bits_id(bus_auto_out_14_aw_bits_id),
    .auto_out_14_aw_bits_addr(bus_auto_out_14_aw_bits_addr),
    .auto_out_14_aw_bits_size(bus_auto_out_14_aw_bits_size),
    .auto_out_14_w_ready(bus_auto_out_14_w_ready),
    .auto_out_14_w_valid(bus_auto_out_14_w_valid),
    .auto_out_14_w_bits_data(bus_auto_out_14_w_bits_data),
    .auto_out_14_w_bits_strb(bus_auto_out_14_w_bits_strb),
    .auto_out_14_w_bits_last(bus_auto_out_14_w_bits_last),
    .auto_out_14_b_ready(bus_auto_out_14_b_ready),
    .auto_out_14_b_valid(bus_auto_out_14_b_valid),
    .auto_out_14_b_bits_id(bus_auto_out_14_b_bits_id),
    .auto_out_14_b_bits_resp(bus_auto_out_14_b_bits_resp),
    .auto_out_14_ar_ready(bus_auto_out_14_ar_ready),
    .auto_out_14_ar_valid(bus_auto_out_14_ar_valid),
    .auto_out_14_ar_bits_id(bus_auto_out_14_ar_bits_id),
    .auto_out_14_ar_bits_addr(bus_auto_out_14_ar_bits_addr),
    .auto_out_14_ar_bits_size(bus_auto_out_14_ar_bits_size),
    .auto_out_14_r_ready(bus_auto_out_14_r_ready),
    .auto_out_14_r_valid(bus_auto_out_14_r_valid),
    .auto_out_14_r_bits_id(bus_auto_out_14_r_bits_id),
    .auto_out_14_r_bits_data(bus_auto_out_14_r_bits_data),
    .auto_out_14_r_bits_resp(bus_auto_out_14_r_bits_resp),
    .auto_out_14_r_bits_last(bus_auto_out_14_r_bits_last),
    .auto_out_13_aw_ready(bus_auto_out_13_aw_ready),
    .auto_out_13_aw_valid(bus_auto_out_13_aw_valid),
    .auto_out_13_aw_bits_id(bus_auto_out_13_aw_bits_id),
    .auto_out_13_aw_bits_addr(bus_auto_out_13_aw_bits_addr),
    .auto_out_13_aw_bits_size(bus_auto_out_13_aw_bits_size),
    .auto_out_13_w_ready(bus_auto_out_13_w_ready),
    .auto_out_13_w_valid(bus_auto_out_13_w_valid),
    .auto_out_13_w_bits_data(bus_auto_out_13_w_bits_data),
    .auto_out_13_w_bits_strb(bus_auto_out_13_w_bits_strb),
    .auto_out_13_w_bits_last(bus_auto_out_13_w_bits_last),
    .auto_out_13_b_ready(bus_auto_out_13_b_ready),
    .auto_out_13_b_valid(bus_auto_out_13_b_valid),
    .auto_out_13_b_bits_id(bus_auto_out_13_b_bits_id),
    .auto_out_13_b_bits_resp(bus_auto_out_13_b_bits_resp),
    .auto_out_13_ar_ready(bus_auto_out_13_ar_ready),
    .auto_out_13_ar_valid(bus_auto_out_13_ar_valid),
    .auto_out_13_ar_bits_id(bus_auto_out_13_ar_bits_id),
    .auto_out_13_ar_bits_addr(bus_auto_out_13_ar_bits_addr),
    .auto_out_13_ar_bits_size(bus_auto_out_13_ar_bits_size),
    .auto_out_13_r_ready(bus_auto_out_13_r_ready),
    .auto_out_13_r_valid(bus_auto_out_13_r_valid),
    .auto_out_13_r_bits_id(bus_auto_out_13_r_bits_id),
    .auto_out_13_r_bits_data(bus_auto_out_13_r_bits_data),
    .auto_out_13_r_bits_resp(bus_auto_out_13_r_bits_resp),
    .auto_out_13_r_bits_last(bus_auto_out_13_r_bits_last),
    .auto_out_12_aw_ready(bus_auto_out_12_aw_ready),
    .auto_out_12_aw_valid(bus_auto_out_12_aw_valid),
    .auto_out_12_aw_bits_id(bus_auto_out_12_aw_bits_id),
    .auto_out_12_aw_bits_addr(bus_auto_out_12_aw_bits_addr),
    .auto_out_12_aw_bits_size(bus_auto_out_12_aw_bits_size),
    .auto_out_12_w_ready(bus_auto_out_12_w_ready),
    .auto_out_12_w_valid(bus_auto_out_12_w_valid),
    .auto_out_12_w_bits_data(bus_auto_out_12_w_bits_data),
    .auto_out_12_w_bits_strb(bus_auto_out_12_w_bits_strb),
    .auto_out_12_w_bits_last(bus_auto_out_12_w_bits_last),
    .auto_out_12_b_ready(bus_auto_out_12_b_ready),
    .auto_out_12_b_valid(bus_auto_out_12_b_valid),
    .auto_out_12_b_bits_id(bus_auto_out_12_b_bits_id),
    .auto_out_12_b_bits_resp(bus_auto_out_12_b_bits_resp),
    .auto_out_12_ar_ready(bus_auto_out_12_ar_ready),
    .auto_out_12_ar_valid(bus_auto_out_12_ar_valid),
    .auto_out_12_ar_bits_id(bus_auto_out_12_ar_bits_id),
    .auto_out_12_ar_bits_addr(bus_auto_out_12_ar_bits_addr),
    .auto_out_12_ar_bits_size(bus_auto_out_12_ar_bits_size),
    .auto_out_12_r_ready(bus_auto_out_12_r_ready),
    .auto_out_12_r_valid(bus_auto_out_12_r_valid),
    .auto_out_12_r_bits_id(bus_auto_out_12_r_bits_id),
    .auto_out_12_r_bits_data(bus_auto_out_12_r_bits_data),
    .auto_out_12_r_bits_resp(bus_auto_out_12_r_bits_resp),
    .auto_out_12_r_bits_last(bus_auto_out_12_r_bits_last),
    .auto_out_11_aw_ready(bus_auto_out_11_aw_ready),
    .auto_out_11_aw_valid(bus_auto_out_11_aw_valid),
    .auto_out_11_aw_bits_id(bus_auto_out_11_aw_bits_id),
    .auto_out_11_aw_bits_addr(bus_auto_out_11_aw_bits_addr),
    .auto_out_11_aw_bits_size(bus_auto_out_11_aw_bits_size),
    .auto_out_11_w_ready(bus_auto_out_11_w_ready),
    .auto_out_11_w_valid(bus_auto_out_11_w_valid),
    .auto_out_11_w_bits_data(bus_auto_out_11_w_bits_data),
    .auto_out_11_w_bits_strb(bus_auto_out_11_w_bits_strb),
    .auto_out_11_w_bits_last(bus_auto_out_11_w_bits_last),
    .auto_out_11_b_ready(bus_auto_out_11_b_ready),
    .auto_out_11_b_valid(bus_auto_out_11_b_valid),
    .auto_out_11_b_bits_id(bus_auto_out_11_b_bits_id),
    .auto_out_11_b_bits_resp(bus_auto_out_11_b_bits_resp),
    .auto_out_11_ar_ready(bus_auto_out_11_ar_ready),
    .auto_out_11_ar_valid(bus_auto_out_11_ar_valid),
    .auto_out_11_ar_bits_id(bus_auto_out_11_ar_bits_id),
    .auto_out_11_ar_bits_addr(bus_auto_out_11_ar_bits_addr),
    .auto_out_11_ar_bits_size(bus_auto_out_11_ar_bits_size),
    .auto_out_11_r_ready(bus_auto_out_11_r_ready),
    .auto_out_11_r_valid(bus_auto_out_11_r_valid),
    .auto_out_11_r_bits_id(bus_auto_out_11_r_bits_id),
    .auto_out_11_r_bits_data(bus_auto_out_11_r_bits_data),
    .auto_out_11_r_bits_resp(bus_auto_out_11_r_bits_resp),
    .auto_out_11_r_bits_last(bus_auto_out_11_r_bits_last),
    .auto_out_10_aw_ready(bus_auto_out_10_aw_ready),
    .auto_out_10_aw_valid(bus_auto_out_10_aw_valid),
    .auto_out_10_aw_bits_id(bus_auto_out_10_aw_bits_id),
    .auto_out_10_aw_bits_addr(bus_auto_out_10_aw_bits_addr),
    .auto_out_10_aw_bits_size(bus_auto_out_10_aw_bits_size),
    .auto_out_10_w_ready(bus_auto_out_10_w_ready),
    .auto_out_10_w_valid(bus_auto_out_10_w_valid),
    .auto_out_10_w_bits_data(bus_auto_out_10_w_bits_data),
    .auto_out_10_w_bits_strb(bus_auto_out_10_w_bits_strb),
    .auto_out_10_w_bits_last(bus_auto_out_10_w_bits_last),
    .auto_out_10_b_ready(bus_auto_out_10_b_ready),
    .auto_out_10_b_valid(bus_auto_out_10_b_valid),
    .auto_out_10_b_bits_id(bus_auto_out_10_b_bits_id),
    .auto_out_10_b_bits_resp(bus_auto_out_10_b_bits_resp),
    .auto_out_10_ar_ready(bus_auto_out_10_ar_ready),
    .auto_out_10_ar_valid(bus_auto_out_10_ar_valid),
    .auto_out_10_ar_bits_id(bus_auto_out_10_ar_bits_id),
    .auto_out_10_ar_bits_addr(bus_auto_out_10_ar_bits_addr),
    .auto_out_10_ar_bits_size(bus_auto_out_10_ar_bits_size),
    .auto_out_10_r_ready(bus_auto_out_10_r_ready),
    .auto_out_10_r_valid(bus_auto_out_10_r_valid),
    .auto_out_10_r_bits_id(bus_auto_out_10_r_bits_id),
    .auto_out_10_r_bits_data(bus_auto_out_10_r_bits_data),
    .auto_out_10_r_bits_resp(bus_auto_out_10_r_bits_resp),
    .auto_out_10_r_bits_last(bus_auto_out_10_r_bits_last),
    .auto_out_9_aw_ready(bus_auto_out_9_aw_ready),
    .auto_out_9_aw_valid(bus_auto_out_9_aw_valid),
    .auto_out_9_aw_bits_id(bus_auto_out_9_aw_bits_id),
    .auto_out_9_aw_bits_addr(bus_auto_out_9_aw_bits_addr),
    .auto_out_9_aw_bits_size(bus_auto_out_9_aw_bits_size),
    .auto_out_9_w_ready(bus_auto_out_9_w_ready),
    .auto_out_9_w_valid(bus_auto_out_9_w_valid),
    .auto_out_9_w_bits_data(bus_auto_out_9_w_bits_data),
    .auto_out_9_w_bits_strb(bus_auto_out_9_w_bits_strb),
    .auto_out_9_w_bits_last(bus_auto_out_9_w_bits_last),
    .auto_out_9_b_ready(bus_auto_out_9_b_ready),
    .auto_out_9_b_valid(bus_auto_out_9_b_valid),
    .auto_out_9_b_bits_id(bus_auto_out_9_b_bits_id),
    .auto_out_9_b_bits_resp(bus_auto_out_9_b_bits_resp),
    .auto_out_9_ar_ready(bus_auto_out_9_ar_ready),
    .auto_out_9_ar_valid(bus_auto_out_9_ar_valid),
    .auto_out_9_ar_bits_id(bus_auto_out_9_ar_bits_id),
    .auto_out_9_ar_bits_addr(bus_auto_out_9_ar_bits_addr),
    .auto_out_9_ar_bits_size(bus_auto_out_9_ar_bits_size),
    .auto_out_9_r_ready(bus_auto_out_9_r_ready),
    .auto_out_9_r_valid(bus_auto_out_9_r_valid),
    .auto_out_9_r_bits_id(bus_auto_out_9_r_bits_id),
    .auto_out_9_r_bits_data(bus_auto_out_9_r_bits_data),
    .auto_out_9_r_bits_resp(bus_auto_out_9_r_bits_resp),
    .auto_out_9_r_bits_last(bus_auto_out_9_r_bits_last),
    .auto_out_8_aw_ready(bus_auto_out_8_aw_ready),
    .auto_out_8_aw_valid(bus_auto_out_8_aw_valid),
    .auto_out_8_aw_bits_id(bus_auto_out_8_aw_bits_id),
    .auto_out_8_aw_bits_addr(bus_auto_out_8_aw_bits_addr),
    .auto_out_8_aw_bits_size(bus_auto_out_8_aw_bits_size),
    .auto_out_8_w_ready(bus_auto_out_8_w_ready),
    .auto_out_8_w_valid(bus_auto_out_8_w_valid),
    .auto_out_8_w_bits_data(bus_auto_out_8_w_bits_data),
    .auto_out_8_w_bits_strb(bus_auto_out_8_w_bits_strb),
    .auto_out_8_w_bits_last(bus_auto_out_8_w_bits_last),
    .auto_out_8_b_ready(bus_auto_out_8_b_ready),
    .auto_out_8_b_valid(bus_auto_out_8_b_valid),
    .auto_out_8_b_bits_id(bus_auto_out_8_b_bits_id),
    .auto_out_8_b_bits_resp(bus_auto_out_8_b_bits_resp),
    .auto_out_8_ar_ready(bus_auto_out_8_ar_ready),
    .auto_out_8_ar_valid(bus_auto_out_8_ar_valid),
    .auto_out_8_ar_bits_id(bus_auto_out_8_ar_bits_id),
    .auto_out_8_ar_bits_addr(bus_auto_out_8_ar_bits_addr),
    .auto_out_8_ar_bits_size(bus_auto_out_8_ar_bits_size),
    .auto_out_8_r_ready(bus_auto_out_8_r_ready),
    .auto_out_8_r_valid(bus_auto_out_8_r_valid),
    .auto_out_8_r_bits_id(bus_auto_out_8_r_bits_id),
    .auto_out_8_r_bits_data(bus_auto_out_8_r_bits_data),
    .auto_out_8_r_bits_resp(bus_auto_out_8_r_bits_resp),
    .auto_out_8_r_bits_last(bus_auto_out_8_r_bits_last),
    .auto_out_7_aw_ready(bus_auto_out_7_aw_ready),
    .auto_out_7_aw_valid(bus_auto_out_7_aw_valid),
    .auto_out_7_aw_bits_id(bus_auto_out_7_aw_bits_id),
    .auto_out_7_aw_bits_addr(bus_auto_out_7_aw_bits_addr),
    .auto_out_7_aw_bits_size(bus_auto_out_7_aw_bits_size),
    .auto_out_7_w_ready(bus_auto_out_7_w_ready),
    .auto_out_7_w_valid(bus_auto_out_7_w_valid),
    .auto_out_7_w_bits_data(bus_auto_out_7_w_bits_data),
    .auto_out_7_w_bits_strb(bus_auto_out_7_w_bits_strb),
    .auto_out_7_w_bits_last(bus_auto_out_7_w_bits_last),
    .auto_out_7_b_ready(bus_auto_out_7_b_ready),
    .auto_out_7_b_valid(bus_auto_out_7_b_valid),
    .auto_out_7_b_bits_id(bus_auto_out_7_b_bits_id),
    .auto_out_7_b_bits_resp(bus_auto_out_7_b_bits_resp),
    .auto_out_7_ar_ready(bus_auto_out_7_ar_ready),
    .auto_out_7_ar_valid(bus_auto_out_7_ar_valid),
    .auto_out_7_ar_bits_id(bus_auto_out_7_ar_bits_id),
    .auto_out_7_ar_bits_addr(bus_auto_out_7_ar_bits_addr),
    .auto_out_7_ar_bits_size(bus_auto_out_7_ar_bits_size),
    .auto_out_7_r_ready(bus_auto_out_7_r_ready),
    .auto_out_7_r_valid(bus_auto_out_7_r_valid),
    .auto_out_7_r_bits_id(bus_auto_out_7_r_bits_id),
    .auto_out_7_r_bits_data(bus_auto_out_7_r_bits_data),
    .auto_out_7_r_bits_resp(bus_auto_out_7_r_bits_resp),
    .auto_out_7_r_bits_last(bus_auto_out_7_r_bits_last),
    .auto_out_6_aw_ready(bus_auto_out_6_aw_ready),
    .auto_out_6_aw_valid(bus_auto_out_6_aw_valid),
    .auto_out_6_aw_bits_id(bus_auto_out_6_aw_bits_id),
    .auto_out_6_aw_bits_addr(bus_auto_out_6_aw_bits_addr),
    .auto_out_6_aw_bits_size(bus_auto_out_6_aw_bits_size),
    .auto_out_6_w_ready(bus_auto_out_6_w_ready),
    .auto_out_6_w_valid(bus_auto_out_6_w_valid),
    .auto_out_6_w_bits_data(bus_auto_out_6_w_bits_data),
    .auto_out_6_w_bits_strb(bus_auto_out_6_w_bits_strb),
    .auto_out_6_w_bits_last(bus_auto_out_6_w_bits_last),
    .auto_out_6_b_ready(bus_auto_out_6_b_ready),
    .auto_out_6_b_valid(bus_auto_out_6_b_valid),
    .auto_out_6_b_bits_id(bus_auto_out_6_b_bits_id),
    .auto_out_6_b_bits_resp(bus_auto_out_6_b_bits_resp),
    .auto_out_6_ar_ready(bus_auto_out_6_ar_ready),
    .auto_out_6_ar_valid(bus_auto_out_6_ar_valid),
    .auto_out_6_ar_bits_id(bus_auto_out_6_ar_bits_id),
    .auto_out_6_ar_bits_addr(bus_auto_out_6_ar_bits_addr),
    .auto_out_6_ar_bits_size(bus_auto_out_6_ar_bits_size),
    .auto_out_6_r_ready(bus_auto_out_6_r_ready),
    .auto_out_6_r_valid(bus_auto_out_6_r_valid),
    .auto_out_6_r_bits_id(bus_auto_out_6_r_bits_id),
    .auto_out_6_r_bits_data(bus_auto_out_6_r_bits_data),
    .auto_out_6_r_bits_resp(bus_auto_out_6_r_bits_resp),
    .auto_out_6_r_bits_last(bus_auto_out_6_r_bits_last),
    .auto_out_5_aw_ready(bus_auto_out_5_aw_ready),
    .auto_out_5_aw_valid(bus_auto_out_5_aw_valid),
    .auto_out_5_aw_bits_id(bus_auto_out_5_aw_bits_id),
    .auto_out_5_aw_bits_addr(bus_auto_out_5_aw_bits_addr),
    .auto_out_5_aw_bits_size(bus_auto_out_5_aw_bits_size),
    .auto_out_5_w_ready(bus_auto_out_5_w_ready),
    .auto_out_5_w_valid(bus_auto_out_5_w_valid),
    .auto_out_5_w_bits_data(bus_auto_out_5_w_bits_data),
    .auto_out_5_w_bits_strb(bus_auto_out_5_w_bits_strb),
    .auto_out_5_w_bits_last(bus_auto_out_5_w_bits_last),
    .auto_out_5_b_ready(bus_auto_out_5_b_ready),
    .auto_out_5_b_valid(bus_auto_out_5_b_valid),
    .auto_out_5_b_bits_id(bus_auto_out_5_b_bits_id),
    .auto_out_5_b_bits_resp(bus_auto_out_5_b_bits_resp),
    .auto_out_5_ar_ready(bus_auto_out_5_ar_ready),
    .auto_out_5_ar_valid(bus_auto_out_5_ar_valid),
    .auto_out_5_ar_bits_id(bus_auto_out_5_ar_bits_id),
    .auto_out_5_ar_bits_addr(bus_auto_out_5_ar_bits_addr),
    .auto_out_5_ar_bits_size(bus_auto_out_5_ar_bits_size),
    .auto_out_5_r_ready(bus_auto_out_5_r_ready),
    .auto_out_5_r_valid(bus_auto_out_5_r_valid),
    .auto_out_5_r_bits_id(bus_auto_out_5_r_bits_id),
    .auto_out_5_r_bits_data(bus_auto_out_5_r_bits_data),
    .auto_out_5_r_bits_resp(bus_auto_out_5_r_bits_resp),
    .auto_out_5_r_bits_last(bus_auto_out_5_r_bits_last),
    .auto_out_4_aw_ready(bus_auto_out_4_aw_ready),
    .auto_out_4_aw_valid(bus_auto_out_4_aw_valid),
    .auto_out_4_aw_bits_id(bus_auto_out_4_aw_bits_id),
    .auto_out_4_aw_bits_addr(bus_auto_out_4_aw_bits_addr),
    .auto_out_4_aw_bits_size(bus_auto_out_4_aw_bits_size),
    .auto_out_4_w_ready(bus_auto_out_4_w_ready),
    .auto_out_4_w_valid(bus_auto_out_4_w_valid),
    .auto_out_4_w_bits_data(bus_auto_out_4_w_bits_data),
    .auto_out_4_w_bits_strb(bus_auto_out_4_w_bits_strb),
    .auto_out_4_w_bits_last(bus_auto_out_4_w_bits_last),
    .auto_out_4_b_ready(bus_auto_out_4_b_ready),
    .auto_out_4_b_valid(bus_auto_out_4_b_valid),
    .auto_out_4_b_bits_id(bus_auto_out_4_b_bits_id),
    .auto_out_4_b_bits_resp(bus_auto_out_4_b_bits_resp),
    .auto_out_4_ar_ready(bus_auto_out_4_ar_ready),
    .auto_out_4_ar_valid(bus_auto_out_4_ar_valid),
    .auto_out_4_ar_bits_id(bus_auto_out_4_ar_bits_id),
    .auto_out_4_ar_bits_addr(bus_auto_out_4_ar_bits_addr),
    .auto_out_4_ar_bits_size(bus_auto_out_4_ar_bits_size),
    .auto_out_4_r_ready(bus_auto_out_4_r_ready),
    .auto_out_4_r_valid(bus_auto_out_4_r_valid),
    .auto_out_4_r_bits_id(bus_auto_out_4_r_bits_id),
    .auto_out_4_r_bits_data(bus_auto_out_4_r_bits_data),
    .auto_out_4_r_bits_resp(bus_auto_out_4_r_bits_resp),
    .auto_out_4_r_bits_last(bus_auto_out_4_r_bits_last),
    .auto_out_3_aw_ready(bus_auto_out_3_aw_ready),
    .auto_out_3_aw_valid(bus_auto_out_3_aw_valid),
    .auto_out_3_aw_bits_id(bus_auto_out_3_aw_bits_id),
    .auto_out_3_aw_bits_addr(bus_auto_out_3_aw_bits_addr),
    .auto_out_3_aw_bits_size(bus_auto_out_3_aw_bits_size),
    .auto_out_3_w_ready(bus_auto_out_3_w_ready),
    .auto_out_3_w_valid(bus_auto_out_3_w_valid),
    .auto_out_3_w_bits_data(bus_auto_out_3_w_bits_data),
    .auto_out_3_w_bits_strb(bus_auto_out_3_w_bits_strb),
    .auto_out_3_w_bits_last(bus_auto_out_3_w_bits_last),
    .auto_out_3_b_ready(bus_auto_out_3_b_ready),
    .auto_out_3_b_valid(bus_auto_out_3_b_valid),
    .auto_out_3_b_bits_id(bus_auto_out_3_b_bits_id),
    .auto_out_3_b_bits_resp(bus_auto_out_3_b_bits_resp),
    .auto_out_3_ar_ready(bus_auto_out_3_ar_ready),
    .auto_out_3_ar_valid(bus_auto_out_3_ar_valid),
    .auto_out_3_ar_bits_id(bus_auto_out_3_ar_bits_id),
    .auto_out_3_ar_bits_addr(bus_auto_out_3_ar_bits_addr),
    .auto_out_3_ar_bits_size(bus_auto_out_3_ar_bits_size),
    .auto_out_3_r_ready(bus_auto_out_3_r_ready),
    .auto_out_3_r_valid(bus_auto_out_3_r_valid),
    .auto_out_3_r_bits_id(bus_auto_out_3_r_bits_id),
    .auto_out_3_r_bits_data(bus_auto_out_3_r_bits_data),
    .auto_out_3_r_bits_resp(bus_auto_out_3_r_bits_resp),
    .auto_out_3_r_bits_last(bus_auto_out_3_r_bits_last),
    .auto_out_2_aw_ready(bus_auto_out_2_aw_ready),
    .auto_out_2_aw_valid(bus_auto_out_2_aw_valid),
    .auto_out_2_aw_bits_id(bus_auto_out_2_aw_bits_id),
    .auto_out_2_aw_bits_addr(bus_auto_out_2_aw_bits_addr),
    .auto_out_2_aw_bits_size(bus_auto_out_2_aw_bits_size),
    .auto_out_2_w_ready(bus_auto_out_2_w_ready),
    .auto_out_2_w_valid(bus_auto_out_2_w_valid),
    .auto_out_2_w_bits_data(bus_auto_out_2_w_bits_data),
    .auto_out_2_w_bits_strb(bus_auto_out_2_w_bits_strb),
    .auto_out_2_w_bits_last(bus_auto_out_2_w_bits_last),
    .auto_out_2_b_ready(bus_auto_out_2_b_ready),
    .auto_out_2_b_valid(bus_auto_out_2_b_valid),
    .auto_out_2_b_bits_id(bus_auto_out_2_b_bits_id),
    .auto_out_2_b_bits_resp(bus_auto_out_2_b_bits_resp),
    .auto_out_2_ar_ready(bus_auto_out_2_ar_ready),
    .auto_out_2_ar_valid(bus_auto_out_2_ar_valid),
    .auto_out_2_ar_bits_id(bus_auto_out_2_ar_bits_id),
    .auto_out_2_ar_bits_addr(bus_auto_out_2_ar_bits_addr),
    .auto_out_2_ar_bits_size(bus_auto_out_2_ar_bits_size),
    .auto_out_2_r_ready(bus_auto_out_2_r_ready),
    .auto_out_2_r_valid(bus_auto_out_2_r_valid),
    .auto_out_2_r_bits_id(bus_auto_out_2_r_bits_id),
    .auto_out_2_r_bits_data(bus_auto_out_2_r_bits_data),
    .auto_out_2_r_bits_resp(bus_auto_out_2_r_bits_resp),
    .auto_out_2_r_bits_last(bus_auto_out_2_r_bits_last),
    .auto_out_1_aw_ready(bus_auto_out_1_aw_ready),
    .auto_out_1_aw_valid(bus_auto_out_1_aw_valid),
    .auto_out_1_aw_bits_id(bus_auto_out_1_aw_bits_id),
    .auto_out_1_aw_bits_addr(bus_auto_out_1_aw_bits_addr),
    .auto_out_1_aw_bits_size(bus_auto_out_1_aw_bits_size),
    .auto_out_1_w_ready(bus_auto_out_1_w_ready),
    .auto_out_1_w_valid(bus_auto_out_1_w_valid),
    .auto_out_1_w_bits_data(bus_auto_out_1_w_bits_data),
    .auto_out_1_w_bits_strb(bus_auto_out_1_w_bits_strb),
    .auto_out_1_w_bits_last(bus_auto_out_1_w_bits_last),
    .auto_out_1_b_ready(bus_auto_out_1_b_ready),
    .auto_out_1_b_valid(bus_auto_out_1_b_valid),
    .auto_out_1_b_bits_id(bus_auto_out_1_b_bits_id),
    .auto_out_1_b_bits_resp(bus_auto_out_1_b_bits_resp),
    .auto_out_1_ar_ready(bus_auto_out_1_ar_ready),
    .auto_out_1_ar_valid(bus_auto_out_1_ar_valid),
    .auto_out_1_ar_bits_id(bus_auto_out_1_ar_bits_id),
    .auto_out_1_ar_bits_addr(bus_auto_out_1_ar_bits_addr),
    .auto_out_1_ar_bits_size(bus_auto_out_1_ar_bits_size),
    .auto_out_1_r_ready(bus_auto_out_1_r_ready),
    .auto_out_1_r_valid(bus_auto_out_1_r_valid),
    .auto_out_1_r_bits_id(bus_auto_out_1_r_bits_id),
    .auto_out_1_r_bits_data(bus_auto_out_1_r_bits_data),
    .auto_out_1_r_bits_resp(bus_auto_out_1_r_bits_resp),
    .auto_out_1_r_bits_last(bus_auto_out_1_r_bits_last),
    .auto_out_0_aw_ready(bus_auto_out_0_aw_ready),
    .auto_out_0_aw_valid(bus_auto_out_0_aw_valid),
    .auto_out_0_aw_bits_id(bus_auto_out_0_aw_bits_id),
    .auto_out_0_aw_bits_addr(bus_auto_out_0_aw_bits_addr),
    .auto_out_0_aw_bits_size(bus_auto_out_0_aw_bits_size),
    .auto_out_0_w_ready(bus_auto_out_0_w_ready),
    .auto_out_0_w_valid(bus_auto_out_0_w_valid),
    .auto_out_0_w_bits_data(bus_auto_out_0_w_bits_data),
    .auto_out_0_w_bits_strb(bus_auto_out_0_w_bits_strb),
    .auto_out_0_w_bits_last(bus_auto_out_0_w_bits_last),
    .auto_out_0_b_ready(bus_auto_out_0_b_ready),
    .auto_out_0_b_valid(bus_auto_out_0_b_valid),
    .auto_out_0_b_bits_id(bus_auto_out_0_b_bits_id),
    .auto_out_0_b_bits_resp(bus_auto_out_0_b_bits_resp),
    .auto_out_0_ar_ready(bus_auto_out_0_ar_ready),
    .auto_out_0_ar_valid(bus_auto_out_0_ar_valid),
    .auto_out_0_ar_bits_id(bus_auto_out_0_ar_bits_id),
    .auto_out_0_ar_bits_addr(bus_auto_out_0_ar_bits_addr),
    .auto_out_0_ar_bits_size(bus_auto_out_0_ar_bits_size),
    .auto_out_0_r_ready(bus_auto_out_0_r_ready),
    .auto_out_0_r_valid(bus_auto_out_0_r_valid),
    .auto_out_0_r_bits_id(bus_auto_out_0_r_bits_id),
    .auto_out_0_r_bits_data(bus_auto_out_0_r_bits_data),
    .auto_out_0_r_bits_resp(bus_auto_out_0_r_bits_resp),
    .auto_out_0_r_bits_last(bus_auto_out_0_r_bits_last)
  );
  AXI4Buffer axi4buf ( // @[Buffer.scala 58:29]
    .clock(axi4buf_clock),
    .reset(axi4buf_reset),
    .auto_in_aw_ready(axi4buf_auto_in_aw_ready),
    .auto_in_aw_valid(axi4buf_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4buf_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4buf_auto_in_aw_bits_addr),
    .auto_in_aw_bits_size(axi4buf_auto_in_aw_bits_size),
    .auto_in_w_ready(axi4buf_auto_in_w_ready),
    .auto_in_w_valid(axi4buf_auto_in_w_valid),
    .auto_in_w_bits_data(axi4buf_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi4buf_auto_in_w_bits_strb),
    .auto_in_w_bits_last(axi4buf_auto_in_w_bits_last),
    .auto_in_b_ready(axi4buf_auto_in_b_ready),
    .auto_in_b_valid(axi4buf_auto_in_b_valid),
    .auto_in_b_bits_id(axi4buf_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi4buf_auto_in_b_bits_resp),
    .auto_in_ar_ready(axi4buf_auto_in_ar_ready),
    .auto_in_ar_valid(axi4buf_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4buf_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4buf_auto_in_ar_bits_addr),
    .auto_in_ar_bits_size(axi4buf_auto_in_ar_bits_size),
    .auto_in_r_ready(axi4buf_auto_in_r_ready),
    .auto_in_r_valid(axi4buf_auto_in_r_valid),
    .auto_in_r_bits_id(axi4buf_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4buf_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4buf_auto_in_r_bits_resp),
    .auto_in_r_bits_last(axi4buf_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4buf_auto_out_aw_ready),
    .auto_out_aw_valid(axi4buf_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4buf_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4buf_auto_out_aw_bits_addr),
    .auto_out_w_ready(axi4buf_auto_out_w_ready),
    .auto_out_w_valid(axi4buf_auto_out_w_valid),
    .auto_out_w_bits_data(axi4buf_auto_out_w_bits_data),
    .auto_out_w_bits_strb(axi4buf_auto_out_w_bits_strb),
    .auto_out_w_bits_last(axi4buf_auto_out_w_bits_last),
    .auto_out_b_ready(axi4buf_auto_out_b_ready),
    .auto_out_b_valid(axi4buf_auto_out_b_valid),
    .auto_out_b_bits_id(axi4buf_auto_out_b_bits_id),
    .auto_out_b_bits_resp(axi4buf_auto_out_b_bits_resp),
    .auto_out_ar_ready(axi4buf_auto_out_ar_ready),
    .auto_out_ar_valid(axi4buf_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4buf_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4buf_auto_out_ar_bits_addr),
    .auto_out_ar_bits_size(axi4buf_auto_out_ar_bits_size),
    .auto_out_r_ready(axi4buf_auto_out_r_ready),
    .auto_out_r_valid(axi4buf_auto_out_r_valid),
    .auto_out_r_bits_id(axi4buf_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4buf_auto_out_r_bits_data),
    .auto_out_r_bits_resp(axi4buf_auto_out_r_bits_resp),
    .auto_out_r_bits_last(axi4buf_auto_out_r_bits_last)
  );
  AXI4Buffer axi4buf_1 ( // @[Buffer.scala 58:29]
    .clock(axi4buf_1_clock),
    .reset(axi4buf_1_reset),
    .auto_in_aw_ready(axi4buf_1_auto_in_aw_ready),
    .auto_in_aw_valid(axi4buf_1_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4buf_1_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4buf_1_auto_in_aw_bits_addr),
    .auto_in_aw_bits_size(axi4buf_1_auto_in_aw_bits_size),
    .auto_in_w_ready(axi4buf_1_auto_in_w_ready),
    .auto_in_w_valid(axi4buf_1_auto_in_w_valid),
    .auto_in_w_bits_data(axi4buf_1_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi4buf_1_auto_in_w_bits_strb),
    .auto_in_w_bits_last(axi4buf_1_auto_in_w_bits_last),
    .auto_in_b_ready(axi4buf_1_auto_in_b_ready),
    .auto_in_b_valid(axi4buf_1_auto_in_b_valid),
    .auto_in_b_bits_id(axi4buf_1_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi4buf_1_auto_in_b_bits_resp),
    .auto_in_ar_ready(axi4buf_1_auto_in_ar_ready),
    .auto_in_ar_valid(axi4buf_1_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4buf_1_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4buf_1_auto_in_ar_bits_addr),
    .auto_in_ar_bits_size(axi4buf_1_auto_in_ar_bits_size),
    .auto_in_r_ready(axi4buf_1_auto_in_r_ready),
    .auto_in_r_valid(axi4buf_1_auto_in_r_valid),
    .auto_in_r_bits_id(axi4buf_1_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4buf_1_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4buf_1_auto_in_r_bits_resp),
    .auto_in_r_bits_last(axi4buf_1_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4buf_1_auto_out_aw_ready),
    .auto_out_aw_valid(axi4buf_1_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4buf_1_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4buf_1_auto_out_aw_bits_addr),
    .auto_out_w_ready(axi4buf_1_auto_out_w_ready),
    .auto_out_w_valid(axi4buf_1_auto_out_w_valid),
    .auto_out_w_bits_data(axi4buf_1_auto_out_w_bits_data),
    .auto_out_w_bits_strb(axi4buf_1_auto_out_w_bits_strb),
    .auto_out_w_bits_last(axi4buf_1_auto_out_w_bits_last),
    .auto_out_b_ready(axi4buf_1_auto_out_b_ready),
    .auto_out_b_valid(axi4buf_1_auto_out_b_valid),
    .auto_out_b_bits_id(axi4buf_1_auto_out_b_bits_id),
    .auto_out_b_bits_resp(axi4buf_1_auto_out_b_bits_resp),
    .auto_out_ar_ready(axi4buf_1_auto_out_ar_ready),
    .auto_out_ar_valid(axi4buf_1_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4buf_1_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4buf_1_auto_out_ar_bits_addr),
    .auto_out_ar_bits_size(axi4buf_1_auto_out_ar_bits_size),
    .auto_out_r_ready(axi4buf_1_auto_out_r_ready),
    .auto_out_r_valid(axi4buf_1_auto_out_r_valid),
    .auto_out_r_bits_id(axi4buf_1_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4buf_1_auto_out_r_bits_data),
    .auto_out_r_bits_resp(axi4buf_1_auto_out_r_bits_resp),
    .auto_out_r_bits_last(axi4buf_1_auto_out_r_bits_last)
  );
  AXI4Buffer axi4buf_2 ( // @[Buffer.scala 58:29]
    .clock(axi4buf_2_clock),
    .reset(axi4buf_2_reset),
    .auto_in_aw_ready(axi4buf_2_auto_in_aw_ready),
    .auto_in_aw_valid(axi4buf_2_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4buf_2_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4buf_2_auto_in_aw_bits_addr),
    .auto_in_aw_bits_size(axi4buf_2_auto_in_aw_bits_size),
    .auto_in_w_ready(axi4buf_2_auto_in_w_ready),
    .auto_in_w_valid(axi4buf_2_auto_in_w_valid),
    .auto_in_w_bits_data(axi4buf_2_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi4buf_2_auto_in_w_bits_strb),
    .auto_in_w_bits_last(axi4buf_2_auto_in_w_bits_last),
    .auto_in_b_ready(axi4buf_2_auto_in_b_ready),
    .auto_in_b_valid(axi4buf_2_auto_in_b_valid),
    .auto_in_b_bits_id(axi4buf_2_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi4buf_2_auto_in_b_bits_resp),
    .auto_in_ar_ready(axi4buf_2_auto_in_ar_ready),
    .auto_in_ar_valid(axi4buf_2_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4buf_2_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4buf_2_auto_in_ar_bits_addr),
    .auto_in_ar_bits_size(axi4buf_2_auto_in_ar_bits_size),
    .auto_in_r_ready(axi4buf_2_auto_in_r_ready),
    .auto_in_r_valid(axi4buf_2_auto_in_r_valid),
    .auto_in_r_bits_id(axi4buf_2_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4buf_2_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4buf_2_auto_in_r_bits_resp),
    .auto_in_r_bits_last(axi4buf_2_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4buf_2_auto_out_aw_ready),
    .auto_out_aw_valid(axi4buf_2_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4buf_2_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4buf_2_auto_out_aw_bits_addr),
    .auto_out_w_ready(axi4buf_2_auto_out_w_ready),
    .auto_out_w_valid(axi4buf_2_auto_out_w_valid),
    .auto_out_w_bits_data(axi4buf_2_auto_out_w_bits_data),
    .auto_out_w_bits_strb(axi4buf_2_auto_out_w_bits_strb),
    .auto_out_w_bits_last(axi4buf_2_auto_out_w_bits_last),
    .auto_out_b_ready(axi4buf_2_auto_out_b_ready),
    .auto_out_b_valid(axi4buf_2_auto_out_b_valid),
    .auto_out_b_bits_id(axi4buf_2_auto_out_b_bits_id),
    .auto_out_b_bits_resp(axi4buf_2_auto_out_b_bits_resp),
    .auto_out_ar_ready(axi4buf_2_auto_out_ar_ready),
    .auto_out_ar_valid(axi4buf_2_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4buf_2_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4buf_2_auto_out_ar_bits_addr),
    .auto_out_ar_bits_size(axi4buf_2_auto_out_ar_bits_size),
    .auto_out_r_ready(axi4buf_2_auto_out_r_ready),
    .auto_out_r_valid(axi4buf_2_auto_out_r_valid),
    .auto_out_r_bits_id(axi4buf_2_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4buf_2_auto_out_r_bits_data),
    .auto_out_r_bits_resp(axi4buf_2_auto_out_r_bits_resp),
    .auto_out_r_bits_last(axi4buf_2_auto_out_r_bits_last)
  );
  AXI4Buffer axi4buf_3 ( // @[Buffer.scala 58:29]
    .clock(axi4buf_3_clock),
    .reset(axi4buf_3_reset),
    .auto_in_aw_ready(axi4buf_3_auto_in_aw_ready),
    .auto_in_aw_valid(axi4buf_3_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4buf_3_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4buf_3_auto_in_aw_bits_addr),
    .auto_in_aw_bits_size(axi4buf_3_auto_in_aw_bits_size),
    .auto_in_w_ready(axi4buf_3_auto_in_w_ready),
    .auto_in_w_valid(axi4buf_3_auto_in_w_valid),
    .auto_in_w_bits_data(axi4buf_3_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi4buf_3_auto_in_w_bits_strb),
    .auto_in_w_bits_last(axi4buf_3_auto_in_w_bits_last),
    .auto_in_b_ready(axi4buf_3_auto_in_b_ready),
    .auto_in_b_valid(axi4buf_3_auto_in_b_valid),
    .auto_in_b_bits_id(axi4buf_3_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi4buf_3_auto_in_b_bits_resp),
    .auto_in_ar_ready(axi4buf_3_auto_in_ar_ready),
    .auto_in_ar_valid(axi4buf_3_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4buf_3_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4buf_3_auto_in_ar_bits_addr),
    .auto_in_ar_bits_size(axi4buf_3_auto_in_ar_bits_size),
    .auto_in_r_ready(axi4buf_3_auto_in_r_ready),
    .auto_in_r_valid(axi4buf_3_auto_in_r_valid),
    .auto_in_r_bits_id(axi4buf_3_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4buf_3_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4buf_3_auto_in_r_bits_resp),
    .auto_in_r_bits_last(axi4buf_3_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4buf_3_auto_out_aw_ready),
    .auto_out_aw_valid(axi4buf_3_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4buf_3_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4buf_3_auto_out_aw_bits_addr),
    .auto_out_w_ready(axi4buf_3_auto_out_w_ready),
    .auto_out_w_valid(axi4buf_3_auto_out_w_valid),
    .auto_out_w_bits_data(axi4buf_3_auto_out_w_bits_data),
    .auto_out_w_bits_strb(axi4buf_3_auto_out_w_bits_strb),
    .auto_out_w_bits_last(axi4buf_3_auto_out_w_bits_last),
    .auto_out_b_ready(axi4buf_3_auto_out_b_ready),
    .auto_out_b_valid(axi4buf_3_auto_out_b_valid),
    .auto_out_b_bits_id(axi4buf_3_auto_out_b_bits_id),
    .auto_out_b_bits_resp(axi4buf_3_auto_out_b_bits_resp),
    .auto_out_ar_ready(axi4buf_3_auto_out_ar_ready),
    .auto_out_ar_valid(axi4buf_3_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4buf_3_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4buf_3_auto_out_ar_bits_addr),
    .auto_out_ar_bits_size(axi4buf_3_auto_out_ar_bits_size),
    .auto_out_r_ready(axi4buf_3_auto_out_r_ready),
    .auto_out_r_valid(axi4buf_3_auto_out_r_valid),
    .auto_out_r_bits_id(axi4buf_3_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4buf_3_auto_out_r_bits_data),
    .auto_out_r_bits_resp(axi4buf_3_auto_out_r_bits_resp),
    .auto_out_r_bits_last(axi4buf_3_auto_out_r_bits_last)
  );
  AXI4Buffer axi4buf_4 ( // @[Buffer.scala 58:29]
    .clock(axi4buf_4_clock),
    .reset(axi4buf_4_reset),
    .auto_in_aw_ready(axi4buf_4_auto_in_aw_ready),
    .auto_in_aw_valid(axi4buf_4_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4buf_4_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4buf_4_auto_in_aw_bits_addr),
    .auto_in_aw_bits_size(axi4buf_4_auto_in_aw_bits_size),
    .auto_in_w_ready(axi4buf_4_auto_in_w_ready),
    .auto_in_w_valid(axi4buf_4_auto_in_w_valid),
    .auto_in_w_bits_data(axi4buf_4_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi4buf_4_auto_in_w_bits_strb),
    .auto_in_w_bits_last(axi4buf_4_auto_in_w_bits_last),
    .auto_in_b_ready(axi4buf_4_auto_in_b_ready),
    .auto_in_b_valid(axi4buf_4_auto_in_b_valid),
    .auto_in_b_bits_id(axi4buf_4_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi4buf_4_auto_in_b_bits_resp),
    .auto_in_ar_ready(axi4buf_4_auto_in_ar_ready),
    .auto_in_ar_valid(axi4buf_4_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4buf_4_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4buf_4_auto_in_ar_bits_addr),
    .auto_in_ar_bits_size(axi4buf_4_auto_in_ar_bits_size),
    .auto_in_r_ready(axi4buf_4_auto_in_r_ready),
    .auto_in_r_valid(axi4buf_4_auto_in_r_valid),
    .auto_in_r_bits_id(axi4buf_4_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4buf_4_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4buf_4_auto_in_r_bits_resp),
    .auto_in_r_bits_last(axi4buf_4_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4buf_4_auto_out_aw_ready),
    .auto_out_aw_valid(axi4buf_4_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4buf_4_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4buf_4_auto_out_aw_bits_addr),
    .auto_out_w_ready(axi4buf_4_auto_out_w_ready),
    .auto_out_w_valid(axi4buf_4_auto_out_w_valid),
    .auto_out_w_bits_data(axi4buf_4_auto_out_w_bits_data),
    .auto_out_w_bits_strb(axi4buf_4_auto_out_w_bits_strb),
    .auto_out_w_bits_last(axi4buf_4_auto_out_w_bits_last),
    .auto_out_b_ready(axi4buf_4_auto_out_b_ready),
    .auto_out_b_valid(axi4buf_4_auto_out_b_valid),
    .auto_out_b_bits_id(axi4buf_4_auto_out_b_bits_id),
    .auto_out_b_bits_resp(axi4buf_4_auto_out_b_bits_resp),
    .auto_out_ar_ready(axi4buf_4_auto_out_ar_ready),
    .auto_out_ar_valid(axi4buf_4_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4buf_4_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4buf_4_auto_out_ar_bits_addr),
    .auto_out_ar_bits_size(axi4buf_4_auto_out_ar_bits_size),
    .auto_out_r_ready(axi4buf_4_auto_out_r_ready),
    .auto_out_r_valid(axi4buf_4_auto_out_r_valid),
    .auto_out_r_bits_id(axi4buf_4_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4buf_4_auto_out_r_bits_data),
    .auto_out_r_bits_resp(axi4buf_4_auto_out_r_bits_resp),
    .auto_out_r_bits_last(axi4buf_4_auto_out_r_bits_last)
  );
  AXI4Buffer axi4buf_5 ( // @[Buffer.scala 58:29]
    .clock(axi4buf_5_clock),
    .reset(axi4buf_5_reset),
    .auto_in_aw_ready(axi4buf_5_auto_in_aw_ready),
    .auto_in_aw_valid(axi4buf_5_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4buf_5_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4buf_5_auto_in_aw_bits_addr),
    .auto_in_aw_bits_size(axi4buf_5_auto_in_aw_bits_size),
    .auto_in_w_ready(axi4buf_5_auto_in_w_ready),
    .auto_in_w_valid(axi4buf_5_auto_in_w_valid),
    .auto_in_w_bits_data(axi4buf_5_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi4buf_5_auto_in_w_bits_strb),
    .auto_in_w_bits_last(axi4buf_5_auto_in_w_bits_last),
    .auto_in_b_ready(axi4buf_5_auto_in_b_ready),
    .auto_in_b_valid(axi4buf_5_auto_in_b_valid),
    .auto_in_b_bits_id(axi4buf_5_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi4buf_5_auto_in_b_bits_resp),
    .auto_in_ar_ready(axi4buf_5_auto_in_ar_ready),
    .auto_in_ar_valid(axi4buf_5_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4buf_5_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4buf_5_auto_in_ar_bits_addr),
    .auto_in_ar_bits_size(axi4buf_5_auto_in_ar_bits_size),
    .auto_in_r_ready(axi4buf_5_auto_in_r_ready),
    .auto_in_r_valid(axi4buf_5_auto_in_r_valid),
    .auto_in_r_bits_id(axi4buf_5_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4buf_5_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4buf_5_auto_in_r_bits_resp),
    .auto_in_r_bits_last(axi4buf_5_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4buf_5_auto_out_aw_ready),
    .auto_out_aw_valid(axi4buf_5_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4buf_5_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4buf_5_auto_out_aw_bits_addr),
    .auto_out_w_ready(axi4buf_5_auto_out_w_ready),
    .auto_out_w_valid(axi4buf_5_auto_out_w_valid),
    .auto_out_w_bits_data(axi4buf_5_auto_out_w_bits_data),
    .auto_out_w_bits_strb(axi4buf_5_auto_out_w_bits_strb),
    .auto_out_w_bits_last(axi4buf_5_auto_out_w_bits_last),
    .auto_out_b_ready(axi4buf_5_auto_out_b_ready),
    .auto_out_b_valid(axi4buf_5_auto_out_b_valid),
    .auto_out_b_bits_id(axi4buf_5_auto_out_b_bits_id),
    .auto_out_b_bits_resp(axi4buf_5_auto_out_b_bits_resp),
    .auto_out_ar_ready(axi4buf_5_auto_out_ar_ready),
    .auto_out_ar_valid(axi4buf_5_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4buf_5_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4buf_5_auto_out_ar_bits_addr),
    .auto_out_ar_bits_size(axi4buf_5_auto_out_ar_bits_size),
    .auto_out_r_ready(axi4buf_5_auto_out_r_ready),
    .auto_out_r_valid(axi4buf_5_auto_out_r_valid),
    .auto_out_r_bits_id(axi4buf_5_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4buf_5_auto_out_r_bits_data),
    .auto_out_r_bits_resp(axi4buf_5_auto_out_r_bits_resp),
    .auto_out_r_bits_last(axi4buf_5_auto_out_r_bits_last)
  );
  AXI4Buffer axi4buf_6 ( // @[Buffer.scala 58:29]
    .clock(axi4buf_6_clock),
    .reset(axi4buf_6_reset),
    .auto_in_aw_ready(axi4buf_6_auto_in_aw_ready),
    .auto_in_aw_valid(axi4buf_6_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4buf_6_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4buf_6_auto_in_aw_bits_addr),
    .auto_in_aw_bits_size(axi4buf_6_auto_in_aw_bits_size),
    .auto_in_w_ready(axi4buf_6_auto_in_w_ready),
    .auto_in_w_valid(axi4buf_6_auto_in_w_valid),
    .auto_in_w_bits_data(axi4buf_6_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi4buf_6_auto_in_w_bits_strb),
    .auto_in_w_bits_last(axi4buf_6_auto_in_w_bits_last),
    .auto_in_b_ready(axi4buf_6_auto_in_b_ready),
    .auto_in_b_valid(axi4buf_6_auto_in_b_valid),
    .auto_in_b_bits_id(axi4buf_6_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi4buf_6_auto_in_b_bits_resp),
    .auto_in_ar_ready(axi4buf_6_auto_in_ar_ready),
    .auto_in_ar_valid(axi4buf_6_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4buf_6_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4buf_6_auto_in_ar_bits_addr),
    .auto_in_ar_bits_size(axi4buf_6_auto_in_ar_bits_size),
    .auto_in_r_ready(axi4buf_6_auto_in_r_ready),
    .auto_in_r_valid(axi4buf_6_auto_in_r_valid),
    .auto_in_r_bits_id(axi4buf_6_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4buf_6_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4buf_6_auto_in_r_bits_resp),
    .auto_in_r_bits_last(axi4buf_6_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4buf_6_auto_out_aw_ready),
    .auto_out_aw_valid(axi4buf_6_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4buf_6_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4buf_6_auto_out_aw_bits_addr),
    .auto_out_w_ready(axi4buf_6_auto_out_w_ready),
    .auto_out_w_valid(axi4buf_6_auto_out_w_valid),
    .auto_out_w_bits_data(axi4buf_6_auto_out_w_bits_data),
    .auto_out_w_bits_strb(axi4buf_6_auto_out_w_bits_strb),
    .auto_out_w_bits_last(axi4buf_6_auto_out_w_bits_last),
    .auto_out_b_ready(axi4buf_6_auto_out_b_ready),
    .auto_out_b_valid(axi4buf_6_auto_out_b_valid),
    .auto_out_b_bits_id(axi4buf_6_auto_out_b_bits_id),
    .auto_out_b_bits_resp(axi4buf_6_auto_out_b_bits_resp),
    .auto_out_ar_ready(axi4buf_6_auto_out_ar_ready),
    .auto_out_ar_valid(axi4buf_6_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4buf_6_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4buf_6_auto_out_ar_bits_addr),
    .auto_out_ar_bits_size(axi4buf_6_auto_out_ar_bits_size),
    .auto_out_r_ready(axi4buf_6_auto_out_r_ready),
    .auto_out_r_valid(axi4buf_6_auto_out_r_valid),
    .auto_out_r_bits_id(axi4buf_6_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4buf_6_auto_out_r_bits_data),
    .auto_out_r_bits_resp(axi4buf_6_auto_out_r_bits_resp),
    .auto_out_r_bits_last(axi4buf_6_auto_out_r_bits_last)
  );
  AXI4Buffer axi4buf_7 ( // @[Buffer.scala 58:29]
    .clock(axi4buf_7_clock),
    .reset(axi4buf_7_reset),
    .auto_in_aw_ready(axi4buf_7_auto_in_aw_ready),
    .auto_in_aw_valid(axi4buf_7_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4buf_7_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4buf_7_auto_in_aw_bits_addr),
    .auto_in_aw_bits_size(axi4buf_7_auto_in_aw_bits_size),
    .auto_in_w_ready(axi4buf_7_auto_in_w_ready),
    .auto_in_w_valid(axi4buf_7_auto_in_w_valid),
    .auto_in_w_bits_data(axi4buf_7_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi4buf_7_auto_in_w_bits_strb),
    .auto_in_w_bits_last(axi4buf_7_auto_in_w_bits_last),
    .auto_in_b_ready(axi4buf_7_auto_in_b_ready),
    .auto_in_b_valid(axi4buf_7_auto_in_b_valid),
    .auto_in_b_bits_id(axi4buf_7_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi4buf_7_auto_in_b_bits_resp),
    .auto_in_ar_ready(axi4buf_7_auto_in_ar_ready),
    .auto_in_ar_valid(axi4buf_7_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4buf_7_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4buf_7_auto_in_ar_bits_addr),
    .auto_in_ar_bits_size(axi4buf_7_auto_in_ar_bits_size),
    .auto_in_r_ready(axi4buf_7_auto_in_r_ready),
    .auto_in_r_valid(axi4buf_7_auto_in_r_valid),
    .auto_in_r_bits_id(axi4buf_7_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4buf_7_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4buf_7_auto_in_r_bits_resp),
    .auto_in_r_bits_last(axi4buf_7_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4buf_7_auto_out_aw_ready),
    .auto_out_aw_valid(axi4buf_7_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4buf_7_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4buf_7_auto_out_aw_bits_addr),
    .auto_out_w_ready(axi4buf_7_auto_out_w_ready),
    .auto_out_w_valid(axi4buf_7_auto_out_w_valid),
    .auto_out_w_bits_data(axi4buf_7_auto_out_w_bits_data),
    .auto_out_w_bits_strb(axi4buf_7_auto_out_w_bits_strb),
    .auto_out_w_bits_last(axi4buf_7_auto_out_w_bits_last),
    .auto_out_b_ready(axi4buf_7_auto_out_b_ready),
    .auto_out_b_valid(axi4buf_7_auto_out_b_valid),
    .auto_out_b_bits_id(axi4buf_7_auto_out_b_bits_id),
    .auto_out_b_bits_resp(axi4buf_7_auto_out_b_bits_resp),
    .auto_out_ar_ready(axi4buf_7_auto_out_ar_ready),
    .auto_out_ar_valid(axi4buf_7_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4buf_7_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4buf_7_auto_out_ar_bits_addr),
    .auto_out_ar_bits_size(axi4buf_7_auto_out_ar_bits_size),
    .auto_out_r_ready(axi4buf_7_auto_out_r_ready),
    .auto_out_r_valid(axi4buf_7_auto_out_r_valid),
    .auto_out_r_bits_id(axi4buf_7_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4buf_7_auto_out_r_bits_data),
    .auto_out_r_bits_resp(axi4buf_7_auto_out_r_bits_resp),
    .auto_out_r_bits_last(axi4buf_7_auto_out_r_bits_last)
  );
  AXI4Buffer axi4buf_8 ( // @[Buffer.scala 58:29]
    .clock(axi4buf_8_clock),
    .reset(axi4buf_8_reset),
    .auto_in_aw_ready(axi4buf_8_auto_in_aw_ready),
    .auto_in_aw_valid(axi4buf_8_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4buf_8_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4buf_8_auto_in_aw_bits_addr),
    .auto_in_aw_bits_size(axi4buf_8_auto_in_aw_bits_size),
    .auto_in_w_ready(axi4buf_8_auto_in_w_ready),
    .auto_in_w_valid(axi4buf_8_auto_in_w_valid),
    .auto_in_w_bits_data(axi4buf_8_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi4buf_8_auto_in_w_bits_strb),
    .auto_in_w_bits_last(axi4buf_8_auto_in_w_bits_last),
    .auto_in_b_ready(axi4buf_8_auto_in_b_ready),
    .auto_in_b_valid(axi4buf_8_auto_in_b_valid),
    .auto_in_b_bits_id(axi4buf_8_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi4buf_8_auto_in_b_bits_resp),
    .auto_in_ar_ready(axi4buf_8_auto_in_ar_ready),
    .auto_in_ar_valid(axi4buf_8_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4buf_8_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4buf_8_auto_in_ar_bits_addr),
    .auto_in_ar_bits_size(axi4buf_8_auto_in_ar_bits_size),
    .auto_in_r_ready(axi4buf_8_auto_in_r_ready),
    .auto_in_r_valid(axi4buf_8_auto_in_r_valid),
    .auto_in_r_bits_id(axi4buf_8_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4buf_8_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4buf_8_auto_in_r_bits_resp),
    .auto_in_r_bits_last(axi4buf_8_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4buf_8_auto_out_aw_ready),
    .auto_out_aw_valid(axi4buf_8_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4buf_8_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4buf_8_auto_out_aw_bits_addr),
    .auto_out_w_ready(axi4buf_8_auto_out_w_ready),
    .auto_out_w_valid(axi4buf_8_auto_out_w_valid),
    .auto_out_w_bits_data(axi4buf_8_auto_out_w_bits_data),
    .auto_out_w_bits_strb(axi4buf_8_auto_out_w_bits_strb),
    .auto_out_w_bits_last(axi4buf_8_auto_out_w_bits_last),
    .auto_out_b_ready(axi4buf_8_auto_out_b_ready),
    .auto_out_b_valid(axi4buf_8_auto_out_b_valid),
    .auto_out_b_bits_id(axi4buf_8_auto_out_b_bits_id),
    .auto_out_b_bits_resp(axi4buf_8_auto_out_b_bits_resp),
    .auto_out_ar_ready(axi4buf_8_auto_out_ar_ready),
    .auto_out_ar_valid(axi4buf_8_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4buf_8_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4buf_8_auto_out_ar_bits_addr),
    .auto_out_ar_bits_size(axi4buf_8_auto_out_ar_bits_size),
    .auto_out_r_ready(axi4buf_8_auto_out_r_ready),
    .auto_out_r_valid(axi4buf_8_auto_out_r_valid),
    .auto_out_r_bits_id(axi4buf_8_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4buf_8_auto_out_r_bits_data),
    .auto_out_r_bits_resp(axi4buf_8_auto_out_r_bits_resp),
    .auto_out_r_bits_last(axi4buf_8_auto_out_r_bits_last)
  );
  AXI4Buffer axi4buf_9 ( // @[Buffer.scala 58:29]
    .clock(axi4buf_9_clock),
    .reset(axi4buf_9_reset),
    .auto_in_aw_ready(axi4buf_9_auto_in_aw_ready),
    .auto_in_aw_valid(axi4buf_9_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4buf_9_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4buf_9_auto_in_aw_bits_addr),
    .auto_in_aw_bits_size(axi4buf_9_auto_in_aw_bits_size),
    .auto_in_w_ready(axi4buf_9_auto_in_w_ready),
    .auto_in_w_valid(axi4buf_9_auto_in_w_valid),
    .auto_in_w_bits_data(axi4buf_9_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi4buf_9_auto_in_w_bits_strb),
    .auto_in_w_bits_last(axi4buf_9_auto_in_w_bits_last),
    .auto_in_b_ready(axi4buf_9_auto_in_b_ready),
    .auto_in_b_valid(axi4buf_9_auto_in_b_valid),
    .auto_in_b_bits_id(axi4buf_9_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi4buf_9_auto_in_b_bits_resp),
    .auto_in_ar_ready(axi4buf_9_auto_in_ar_ready),
    .auto_in_ar_valid(axi4buf_9_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4buf_9_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4buf_9_auto_in_ar_bits_addr),
    .auto_in_ar_bits_size(axi4buf_9_auto_in_ar_bits_size),
    .auto_in_r_ready(axi4buf_9_auto_in_r_ready),
    .auto_in_r_valid(axi4buf_9_auto_in_r_valid),
    .auto_in_r_bits_id(axi4buf_9_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4buf_9_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4buf_9_auto_in_r_bits_resp),
    .auto_in_r_bits_last(axi4buf_9_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4buf_9_auto_out_aw_ready),
    .auto_out_aw_valid(axi4buf_9_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4buf_9_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4buf_9_auto_out_aw_bits_addr),
    .auto_out_w_ready(axi4buf_9_auto_out_w_ready),
    .auto_out_w_valid(axi4buf_9_auto_out_w_valid),
    .auto_out_w_bits_data(axi4buf_9_auto_out_w_bits_data),
    .auto_out_w_bits_strb(axi4buf_9_auto_out_w_bits_strb),
    .auto_out_w_bits_last(axi4buf_9_auto_out_w_bits_last),
    .auto_out_b_ready(axi4buf_9_auto_out_b_ready),
    .auto_out_b_valid(axi4buf_9_auto_out_b_valid),
    .auto_out_b_bits_id(axi4buf_9_auto_out_b_bits_id),
    .auto_out_b_bits_resp(axi4buf_9_auto_out_b_bits_resp),
    .auto_out_ar_ready(axi4buf_9_auto_out_ar_ready),
    .auto_out_ar_valid(axi4buf_9_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4buf_9_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4buf_9_auto_out_ar_bits_addr),
    .auto_out_ar_bits_size(axi4buf_9_auto_out_ar_bits_size),
    .auto_out_r_ready(axi4buf_9_auto_out_r_ready),
    .auto_out_r_valid(axi4buf_9_auto_out_r_valid),
    .auto_out_r_bits_id(axi4buf_9_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4buf_9_auto_out_r_bits_data),
    .auto_out_r_bits_resp(axi4buf_9_auto_out_r_bits_resp),
    .auto_out_r_bits_last(axi4buf_9_auto_out_r_bits_last)
  );
  AXI4Buffer axi4buf_10 ( // @[Buffer.scala 58:29]
    .clock(axi4buf_10_clock),
    .reset(axi4buf_10_reset),
    .auto_in_aw_ready(axi4buf_10_auto_in_aw_ready),
    .auto_in_aw_valid(axi4buf_10_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4buf_10_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4buf_10_auto_in_aw_bits_addr),
    .auto_in_aw_bits_size(axi4buf_10_auto_in_aw_bits_size),
    .auto_in_w_ready(axi4buf_10_auto_in_w_ready),
    .auto_in_w_valid(axi4buf_10_auto_in_w_valid),
    .auto_in_w_bits_data(axi4buf_10_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi4buf_10_auto_in_w_bits_strb),
    .auto_in_w_bits_last(axi4buf_10_auto_in_w_bits_last),
    .auto_in_b_ready(axi4buf_10_auto_in_b_ready),
    .auto_in_b_valid(axi4buf_10_auto_in_b_valid),
    .auto_in_b_bits_id(axi4buf_10_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi4buf_10_auto_in_b_bits_resp),
    .auto_in_ar_ready(axi4buf_10_auto_in_ar_ready),
    .auto_in_ar_valid(axi4buf_10_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4buf_10_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4buf_10_auto_in_ar_bits_addr),
    .auto_in_ar_bits_size(axi4buf_10_auto_in_ar_bits_size),
    .auto_in_r_ready(axi4buf_10_auto_in_r_ready),
    .auto_in_r_valid(axi4buf_10_auto_in_r_valid),
    .auto_in_r_bits_id(axi4buf_10_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4buf_10_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4buf_10_auto_in_r_bits_resp),
    .auto_in_r_bits_last(axi4buf_10_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4buf_10_auto_out_aw_ready),
    .auto_out_aw_valid(axi4buf_10_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4buf_10_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4buf_10_auto_out_aw_bits_addr),
    .auto_out_w_ready(axi4buf_10_auto_out_w_ready),
    .auto_out_w_valid(axi4buf_10_auto_out_w_valid),
    .auto_out_w_bits_data(axi4buf_10_auto_out_w_bits_data),
    .auto_out_w_bits_strb(axi4buf_10_auto_out_w_bits_strb),
    .auto_out_w_bits_last(axi4buf_10_auto_out_w_bits_last),
    .auto_out_b_ready(axi4buf_10_auto_out_b_ready),
    .auto_out_b_valid(axi4buf_10_auto_out_b_valid),
    .auto_out_b_bits_id(axi4buf_10_auto_out_b_bits_id),
    .auto_out_b_bits_resp(axi4buf_10_auto_out_b_bits_resp),
    .auto_out_ar_ready(axi4buf_10_auto_out_ar_ready),
    .auto_out_ar_valid(axi4buf_10_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4buf_10_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4buf_10_auto_out_ar_bits_addr),
    .auto_out_ar_bits_size(axi4buf_10_auto_out_ar_bits_size),
    .auto_out_r_ready(axi4buf_10_auto_out_r_ready),
    .auto_out_r_valid(axi4buf_10_auto_out_r_valid),
    .auto_out_r_bits_id(axi4buf_10_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4buf_10_auto_out_r_bits_data),
    .auto_out_r_bits_resp(axi4buf_10_auto_out_r_bits_resp),
    .auto_out_r_bits_last(axi4buf_10_auto_out_r_bits_last)
  );
  AXI4Buffer axi4buf_11 ( // @[Buffer.scala 58:29]
    .clock(axi4buf_11_clock),
    .reset(axi4buf_11_reset),
    .auto_in_aw_ready(axi4buf_11_auto_in_aw_ready),
    .auto_in_aw_valid(axi4buf_11_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4buf_11_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4buf_11_auto_in_aw_bits_addr),
    .auto_in_aw_bits_size(axi4buf_11_auto_in_aw_bits_size),
    .auto_in_w_ready(axi4buf_11_auto_in_w_ready),
    .auto_in_w_valid(axi4buf_11_auto_in_w_valid),
    .auto_in_w_bits_data(axi4buf_11_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi4buf_11_auto_in_w_bits_strb),
    .auto_in_w_bits_last(axi4buf_11_auto_in_w_bits_last),
    .auto_in_b_ready(axi4buf_11_auto_in_b_ready),
    .auto_in_b_valid(axi4buf_11_auto_in_b_valid),
    .auto_in_b_bits_id(axi4buf_11_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi4buf_11_auto_in_b_bits_resp),
    .auto_in_ar_ready(axi4buf_11_auto_in_ar_ready),
    .auto_in_ar_valid(axi4buf_11_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4buf_11_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4buf_11_auto_in_ar_bits_addr),
    .auto_in_ar_bits_size(axi4buf_11_auto_in_ar_bits_size),
    .auto_in_r_ready(axi4buf_11_auto_in_r_ready),
    .auto_in_r_valid(axi4buf_11_auto_in_r_valid),
    .auto_in_r_bits_id(axi4buf_11_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4buf_11_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4buf_11_auto_in_r_bits_resp),
    .auto_in_r_bits_last(axi4buf_11_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4buf_11_auto_out_aw_ready),
    .auto_out_aw_valid(axi4buf_11_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4buf_11_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4buf_11_auto_out_aw_bits_addr),
    .auto_out_w_ready(axi4buf_11_auto_out_w_ready),
    .auto_out_w_valid(axi4buf_11_auto_out_w_valid),
    .auto_out_w_bits_data(axi4buf_11_auto_out_w_bits_data),
    .auto_out_w_bits_strb(axi4buf_11_auto_out_w_bits_strb),
    .auto_out_w_bits_last(axi4buf_11_auto_out_w_bits_last),
    .auto_out_b_ready(axi4buf_11_auto_out_b_ready),
    .auto_out_b_valid(axi4buf_11_auto_out_b_valid),
    .auto_out_b_bits_id(axi4buf_11_auto_out_b_bits_id),
    .auto_out_b_bits_resp(axi4buf_11_auto_out_b_bits_resp),
    .auto_out_ar_ready(axi4buf_11_auto_out_ar_ready),
    .auto_out_ar_valid(axi4buf_11_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4buf_11_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4buf_11_auto_out_ar_bits_addr),
    .auto_out_ar_bits_size(axi4buf_11_auto_out_ar_bits_size),
    .auto_out_r_ready(axi4buf_11_auto_out_r_ready),
    .auto_out_r_valid(axi4buf_11_auto_out_r_valid),
    .auto_out_r_bits_id(axi4buf_11_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4buf_11_auto_out_r_bits_data),
    .auto_out_r_bits_resp(axi4buf_11_auto_out_r_bits_resp),
    .auto_out_r_bits_last(axi4buf_11_auto_out_r_bits_last)
  );
  AXI4Buffer axi4buf_12 ( // @[Buffer.scala 58:29]
    .clock(axi4buf_12_clock),
    .reset(axi4buf_12_reset),
    .auto_in_aw_ready(axi4buf_12_auto_in_aw_ready),
    .auto_in_aw_valid(axi4buf_12_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4buf_12_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4buf_12_auto_in_aw_bits_addr),
    .auto_in_aw_bits_size(axi4buf_12_auto_in_aw_bits_size),
    .auto_in_w_ready(axi4buf_12_auto_in_w_ready),
    .auto_in_w_valid(axi4buf_12_auto_in_w_valid),
    .auto_in_w_bits_data(axi4buf_12_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi4buf_12_auto_in_w_bits_strb),
    .auto_in_w_bits_last(axi4buf_12_auto_in_w_bits_last),
    .auto_in_b_ready(axi4buf_12_auto_in_b_ready),
    .auto_in_b_valid(axi4buf_12_auto_in_b_valid),
    .auto_in_b_bits_id(axi4buf_12_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi4buf_12_auto_in_b_bits_resp),
    .auto_in_ar_ready(axi4buf_12_auto_in_ar_ready),
    .auto_in_ar_valid(axi4buf_12_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4buf_12_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4buf_12_auto_in_ar_bits_addr),
    .auto_in_ar_bits_size(axi4buf_12_auto_in_ar_bits_size),
    .auto_in_r_ready(axi4buf_12_auto_in_r_ready),
    .auto_in_r_valid(axi4buf_12_auto_in_r_valid),
    .auto_in_r_bits_id(axi4buf_12_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4buf_12_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4buf_12_auto_in_r_bits_resp),
    .auto_in_r_bits_last(axi4buf_12_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4buf_12_auto_out_aw_ready),
    .auto_out_aw_valid(axi4buf_12_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4buf_12_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4buf_12_auto_out_aw_bits_addr),
    .auto_out_w_ready(axi4buf_12_auto_out_w_ready),
    .auto_out_w_valid(axi4buf_12_auto_out_w_valid),
    .auto_out_w_bits_data(axi4buf_12_auto_out_w_bits_data),
    .auto_out_w_bits_strb(axi4buf_12_auto_out_w_bits_strb),
    .auto_out_w_bits_last(axi4buf_12_auto_out_w_bits_last),
    .auto_out_b_ready(axi4buf_12_auto_out_b_ready),
    .auto_out_b_valid(axi4buf_12_auto_out_b_valid),
    .auto_out_b_bits_id(axi4buf_12_auto_out_b_bits_id),
    .auto_out_b_bits_resp(axi4buf_12_auto_out_b_bits_resp),
    .auto_out_ar_ready(axi4buf_12_auto_out_ar_ready),
    .auto_out_ar_valid(axi4buf_12_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4buf_12_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4buf_12_auto_out_ar_bits_addr),
    .auto_out_ar_bits_size(axi4buf_12_auto_out_ar_bits_size),
    .auto_out_r_ready(axi4buf_12_auto_out_r_ready),
    .auto_out_r_valid(axi4buf_12_auto_out_r_valid),
    .auto_out_r_bits_id(axi4buf_12_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4buf_12_auto_out_r_bits_data),
    .auto_out_r_bits_resp(axi4buf_12_auto_out_r_bits_resp),
    .auto_out_r_bits_last(axi4buf_12_auto_out_r_bits_last)
  );
  AXI4Buffer axi4buf_13 ( // @[Buffer.scala 58:29]
    .clock(axi4buf_13_clock),
    .reset(axi4buf_13_reset),
    .auto_in_aw_ready(axi4buf_13_auto_in_aw_ready),
    .auto_in_aw_valid(axi4buf_13_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4buf_13_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4buf_13_auto_in_aw_bits_addr),
    .auto_in_aw_bits_size(axi4buf_13_auto_in_aw_bits_size),
    .auto_in_w_ready(axi4buf_13_auto_in_w_ready),
    .auto_in_w_valid(axi4buf_13_auto_in_w_valid),
    .auto_in_w_bits_data(axi4buf_13_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi4buf_13_auto_in_w_bits_strb),
    .auto_in_w_bits_last(axi4buf_13_auto_in_w_bits_last),
    .auto_in_b_ready(axi4buf_13_auto_in_b_ready),
    .auto_in_b_valid(axi4buf_13_auto_in_b_valid),
    .auto_in_b_bits_id(axi4buf_13_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi4buf_13_auto_in_b_bits_resp),
    .auto_in_ar_ready(axi4buf_13_auto_in_ar_ready),
    .auto_in_ar_valid(axi4buf_13_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4buf_13_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4buf_13_auto_in_ar_bits_addr),
    .auto_in_ar_bits_size(axi4buf_13_auto_in_ar_bits_size),
    .auto_in_r_ready(axi4buf_13_auto_in_r_ready),
    .auto_in_r_valid(axi4buf_13_auto_in_r_valid),
    .auto_in_r_bits_id(axi4buf_13_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4buf_13_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4buf_13_auto_in_r_bits_resp),
    .auto_in_r_bits_last(axi4buf_13_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4buf_13_auto_out_aw_ready),
    .auto_out_aw_valid(axi4buf_13_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4buf_13_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4buf_13_auto_out_aw_bits_addr),
    .auto_out_w_ready(axi4buf_13_auto_out_w_ready),
    .auto_out_w_valid(axi4buf_13_auto_out_w_valid),
    .auto_out_w_bits_data(axi4buf_13_auto_out_w_bits_data),
    .auto_out_w_bits_strb(axi4buf_13_auto_out_w_bits_strb),
    .auto_out_w_bits_last(axi4buf_13_auto_out_w_bits_last),
    .auto_out_b_ready(axi4buf_13_auto_out_b_ready),
    .auto_out_b_valid(axi4buf_13_auto_out_b_valid),
    .auto_out_b_bits_id(axi4buf_13_auto_out_b_bits_id),
    .auto_out_b_bits_resp(axi4buf_13_auto_out_b_bits_resp),
    .auto_out_ar_ready(axi4buf_13_auto_out_ar_ready),
    .auto_out_ar_valid(axi4buf_13_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4buf_13_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4buf_13_auto_out_ar_bits_addr),
    .auto_out_ar_bits_size(axi4buf_13_auto_out_ar_bits_size),
    .auto_out_r_ready(axi4buf_13_auto_out_r_ready),
    .auto_out_r_valid(axi4buf_13_auto_out_r_valid),
    .auto_out_r_bits_id(axi4buf_13_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4buf_13_auto_out_r_bits_data),
    .auto_out_r_bits_resp(axi4buf_13_auto_out_r_bits_resp),
    .auto_out_r_bits_last(axi4buf_13_auto_out_r_bits_last)
  );
  AXI4Buffer axi4buf_14 ( // @[Buffer.scala 58:29]
    .clock(axi4buf_14_clock),
    .reset(axi4buf_14_reset),
    .auto_in_aw_ready(axi4buf_14_auto_in_aw_ready),
    .auto_in_aw_valid(axi4buf_14_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4buf_14_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4buf_14_auto_in_aw_bits_addr),
    .auto_in_aw_bits_size(axi4buf_14_auto_in_aw_bits_size),
    .auto_in_w_ready(axi4buf_14_auto_in_w_ready),
    .auto_in_w_valid(axi4buf_14_auto_in_w_valid),
    .auto_in_w_bits_data(axi4buf_14_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi4buf_14_auto_in_w_bits_strb),
    .auto_in_w_bits_last(axi4buf_14_auto_in_w_bits_last),
    .auto_in_b_ready(axi4buf_14_auto_in_b_ready),
    .auto_in_b_valid(axi4buf_14_auto_in_b_valid),
    .auto_in_b_bits_id(axi4buf_14_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi4buf_14_auto_in_b_bits_resp),
    .auto_in_ar_ready(axi4buf_14_auto_in_ar_ready),
    .auto_in_ar_valid(axi4buf_14_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4buf_14_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4buf_14_auto_in_ar_bits_addr),
    .auto_in_ar_bits_size(axi4buf_14_auto_in_ar_bits_size),
    .auto_in_r_ready(axi4buf_14_auto_in_r_ready),
    .auto_in_r_valid(axi4buf_14_auto_in_r_valid),
    .auto_in_r_bits_id(axi4buf_14_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4buf_14_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4buf_14_auto_in_r_bits_resp),
    .auto_in_r_bits_last(axi4buf_14_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4buf_14_auto_out_aw_ready),
    .auto_out_aw_valid(axi4buf_14_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4buf_14_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4buf_14_auto_out_aw_bits_addr),
    .auto_out_w_ready(axi4buf_14_auto_out_w_ready),
    .auto_out_w_valid(axi4buf_14_auto_out_w_valid),
    .auto_out_w_bits_data(axi4buf_14_auto_out_w_bits_data),
    .auto_out_w_bits_strb(axi4buf_14_auto_out_w_bits_strb),
    .auto_out_w_bits_last(axi4buf_14_auto_out_w_bits_last),
    .auto_out_b_ready(axi4buf_14_auto_out_b_ready),
    .auto_out_b_valid(axi4buf_14_auto_out_b_valid),
    .auto_out_b_bits_id(axi4buf_14_auto_out_b_bits_id),
    .auto_out_b_bits_resp(axi4buf_14_auto_out_b_bits_resp),
    .auto_out_ar_ready(axi4buf_14_auto_out_ar_ready),
    .auto_out_ar_valid(axi4buf_14_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4buf_14_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4buf_14_auto_out_ar_bits_addr),
    .auto_out_ar_bits_size(axi4buf_14_auto_out_ar_bits_size),
    .auto_out_r_ready(axi4buf_14_auto_out_r_ready),
    .auto_out_r_valid(axi4buf_14_auto_out_r_valid),
    .auto_out_r_bits_id(axi4buf_14_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4buf_14_auto_out_r_bits_data),
    .auto_out_r_bits_resp(axi4buf_14_auto_out_r_bits_resp),
    .auto_out_r_bits_last(axi4buf_14_auto_out_r_bits_last)
  );
  AXI4Buffer axi4buf_15 ( // @[Buffer.scala 58:29]
    .clock(axi4buf_15_clock),
    .reset(axi4buf_15_reset),
    .auto_in_aw_ready(axi4buf_15_auto_in_aw_ready),
    .auto_in_aw_valid(axi4buf_15_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4buf_15_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4buf_15_auto_in_aw_bits_addr),
    .auto_in_aw_bits_size(axi4buf_15_auto_in_aw_bits_size),
    .auto_in_w_ready(axi4buf_15_auto_in_w_ready),
    .auto_in_w_valid(axi4buf_15_auto_in_w_valid),
    .auto_in_w_bits_data(axi4buf_15_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi4buf_15_auto_in_w_bits_strb),
    .auto_in_w_bits_last(axi4buf_15_auto_in_w_bits_last),
    .auto_in_b_ready(axi4buf_15_auto_in_b_ready),
    .auto_in_b_valid(axi4buf_15_auto_in_b_valid),
    .auto_in_b_bits_id(axi4buf_15_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi4buf_15_auto_in_b_bits_resp),
    .auto_in_ar_ready(axi4buf_15_auto_in_ar_ready),
    .auto_in_ar_valid(axi4buf_15_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4buf_15_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4buf_15_auto_in_ar_bits_addr),
    .auto_in_ar_bits_size(axi4buf_15_auto_in_ar_bits_size),
    .auto_in_r_ready(axi4buf_15_auto_in_r_ready),
    .auto_in_r_valid(axi4buf_15_auto_in_r_valid),
    .auto_in_r_bits_id(axi4buf_15_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4buf_15_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4buf_15_auto_in_r_bits_resp),
    .auto_in_r_bits_last(axi4buf_15_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4buf_15_auto_out_aw_ready),
    .auto_out_aw_valid(axi4buf_15_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4buf_15_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4buf_15_auto_out_aw_bits_addr),
    .auto_out_w_ready(axi4buf_15_auto_out_w_ready),
    .auto_out_w_valid(axi4buf_15_auto_out_w_valid),
    .auto_out_w_bits_data(axi4buf_15_auto_out_w_bits_data),
    .auto_out_w_bits_strb(axi4buf_15_auto_out_w_bits_strb),
    .auto_out_w_bits_last(axi4buf_15_auto_out_w_bits_last),
    .auto_out_b_ready(axi4buf_15_auto_out_b_ready),
    .auto_out_b_valid(axi4buf_15_auto_out_b_valid),
    .auto_out_b_bits_id(axi4buf_15_auto_out_b_bits_id),
    .auto_out_b_bits_resp(axi4buf_15_auto_out_b_bits_resp),
    .auto_out_ar_ready(axi4buf_15_auto_out_ar_ready),
    .auto_out_ar_valid(axi4buf_15_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4buf_15_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4buf_15_auto_out_ar_bits_addr),
    .auto_out_ar_bits_size(axi4buf_15_auto_out_ar_bits_size),
    .auto_out_r_ready(axi4buf_15_auto_out_r_ready),
    .auto_out_r_valid(axi4buf_15_auto_out_r_valid),
    .auto_out_r_bits_id(axi4buf_15_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4buf_15_auto_out_r_bits_data),
    .auto_out_r_bits_resp(axi4buf_15_auto_out_r_bits_resp),
    .auto_out_r_bits_last(axi4buf_15_auto_out_r_bits_last)
  );
  AXI4Buffer axi4buf_16 ( // @[Buffer.scala 58:29]
    .clock(axi4buf_16_clock),
    .reset(axi4buf_16_reset),
    .auto_in_aw_ready(axi4buf_16_auto_in_aw_ready),
    .auto_in_aw_valid(axi4buf_16_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4buf_16_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4buf_16_auto_in_aw_bits_addr),
    .auto_in_aw_bits_size(axi4buf_16_auto_in_aw_bits_size),
    .auto_in_w_ready(axi4buf_16_auto_in_w_ready),
    .auto_in_w_valid(axi4buf_16_auto_in_w_valid),
    .auto_in_w_bits_data(axi4buf_16_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi4buf_16_auto_in_w_bits_strb),
    .auto_in_w_bits_last(axi4buf_16_auto_in_w_bits_last),
    .auto_in_b_ready(axi4buf_16_auto_in_b_ready),
    .auto_in_b_valid(axi4buf_16_auto_in_b_valid),
    .auto_in_b_bits_id(axi4buf_16_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi4buf_16_auto_in_b_bits_resp),
    .auto_in_ar_ready(axi4buf_16_auto_in_ar_ready),
    .auto_in_ar_valid(axi4buf_16_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4buf_16_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4buf_16_auto_in_ar_bits_addr),
    .auto_in_ar_bits_size(axi4buf_16_auto_in_ar_bits_size),
    .auto_in_r_ready(axi4buf_16_auto_in_r_ready),
    .auto_in_r_valid(axi4buf_16_auto_in_r_valid),
    .auto_in_r_bits_id(axi4buf_16_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4buf_16_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4buf_16_auto_in_r_bits_resp),
    .auto_in_r_bits_last(axi4buf_16_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4buf_16_auto_out_aw_ready),
    .auto_out_aw_valid(axi4buf_16_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4buf_16_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4buf_16_auto_out_aw_bits_addr),
    .auto_out_w_ready(axi4buf_16_auto_out_w_ready),
    .auto_out_w_valid(axi4buf_16_auto_out_w_valid),
    .auto_out_w_bits_data(axi4buf_16_auto_out_w_bits_data),
    .auto_out_w_bits_strb(axi4buf_16_auto_out_w_bits_strb),
    .auto_out_w_bits_last(axi4buf_16_auto_out_w_bits_last),
    .auto_out_b_ready(axi4buf_16_auto_out_b_ready),
    .auto_out_b_valid(axi4buf_16_auto_out_b_valid),
    .auto_out_b_bits_id(axi4buf_16_auto_out_b_bits_id),
    .auto_out_b_bits_resp(axi4buf_16_auto_out_b_bits_resp),
    .auto_out_ar_ready(axi4buf_16_auto_out_ar_ready),
    .auto_out_ar_valid(axi4buf_16_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4buf_16_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4buf_16_auto_out_ar_bits_addr),
    .auto_out_ar_bits_size(axi4buf_16_auto_out_ar_bits_size),
    .auto_out_r_ready(axi4buf_16_auto_out_r_ready),
    .auto_out_r_valid(axi4buf_16_auto_out_r_valid),
    .auto_out_r_bits_id(axi4buf_16_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4buf_16_auto_out_r_bits_data),
    .auto_out_r_bits_resp(axi4buf_16_auto_out_r_bits_resp),
    .auto_out_r_bits_last(axi4buf_16_auto_out_r_bits_last)
  );
  AXI4Buffer axi4buf_17 ( // @[Buffer.scala 58:29]
    .clock(axi4buf_17_clock),
    .reset(axi4buf_17_reset),
    .auto_in_aw_ready(axi4buf_17_auto_in_aw_ready),
    .auto_in_aw_valid(axi4buf_17_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4buf_17_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4buf_17_auto_in_aw_bits_addr),
    .auto_in_aw_bits_size(axi4buf_17_auto_in_aw_bits_size),
    .auto_in_w_ready(axi4buf_17_auto_in_w_ready),
    .auto_in_w_valid(axi4buf_17_auto_in_w_valid),
    .auto_in_w_bits_data(axi4buf_17_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi4buf_17_auto_in_w_bits_strb),
    .auto_in_w_bits_last(axi4buf_17_auto_in_w_bits_last),
    .auto_in_b_ready(axi4buf_17_auto_in_b_ready),
    .auto_in_b_valid(axi4buf_17_auto_in_b_valid),
    .auto_in_b_bits_id(axi4buf_17_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi4buf_17_auto_in_b_bits_resp),
    .auto_in_ar_ready(axi4buf_17_auto_in_ar_ready),
    .auto_in_ar_valid(axi4buf_17_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4buf_17_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4buf_17_auto_in_ar_bits_addr),
    .auto_in_ar_bits_size(axi4buf_17_auto_in_ar_bits_size),
    .auto_in_r_ready(axi4buf_17_auto_in_r_ready),
    .auto_in_r_valid(axi4buf_17_auto_in_r_valid),
    .auto_in_r_bits_id(axi4buf_17_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4buf_17_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4buf_17_auto_in_r_bits_resp),
    .auto_in_r_bits_last(axi4buf_17_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4buf_17_auto_out_aw_ready),
    .auto_out_aw_valid(axi4buf_17_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4buf_17_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4buf_17_auto_out_aw_bits_addr),
    .auto_out_w_ready(axi4buf_17_auto_out_w_ready),
    .auto_out_w_valid(axi4buf_17_auto_out_w_valid),
    .auto_out_w_bits_data(axi4buf_17_auto_out_w_bits_data),
    .auto_out_w_bits_strb(axi4buf_17_auto_out_w_bits_strb),
    .auto_out_w_bits_last(axi4buf_17_auto_out_w_bits_last),
    .auto_out_b_ready(axi4buf_17_auto_out_b_ready),
    .auto_out_b_valid(axi4buf_17_auto_out_b_valid),
    .auto_out_b_bits_id(axi4buf_17_auto_out_b_bits_id),
    .auto_out_b_bits_resp(axi4buf_17_auto_out_b_bits_resp),
    .auto_out_ar_ready(axi4buf_17_auto_out_ar_ready),
    .auto_out_ar_valid(axi4buf_17_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4buf_17_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4buf_17_auto_out_ar_bits_addr),
    .auto_out_ar_bits_size(axi4buf_17_auto_out_ar_bits_size),
    .auto_out_r_ready(axi4buf_17_auto_out_r_ready),
    .auto_out_r_valid(axi4buf_17_auto_out_r_valid),
    .auto_out_r_bits_id(axi4buf_17_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4buf_17_auto_out_r_bits_data),
    .auto_out_r_bits_resp(axi4buf_17_auto_out_r_bits_resp),
    .auto_out_r_bits_last(axi4buf_17_auto_out_r_bits_last)
  );
  AXI4Buffer axi4buf_18 ( // @[Buffer.scala 58:29]
    .clock(axi4buf_18_clock),
    .reset(axi4buf_18_reset),
    .auto_in_aw_ready(axi4buf_18_auto_in_aw_ready),
    .auto_in_aw_valid(axi4buf_18_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4buf_18_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4buf_18_auto_in_aw_bits_addr),
    .auto_in_aw_bits_size(axi4buf_18_auto_in_aw_bits_size),
    .auto_in_w_ready(axi4buf_18_auto_in_w_ready),
    .auto_in_w_valid(axi4buf_18_auto_in_w_valid),
    .auto_in_w_bits_data(axi4buf_18_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi4buf_18_auto_in_w_bits_strb),
    .auto_in_w_bits_last(axi4buf_18_auto_in_w_bits_last),
    .auto_in_b_ready(axi4buf_18_auto_in_b_ready),
    .auto_in_b_valid(axi4buf_18_auto_in_b_valid),
    .auto_in_b_bits_id(axi4buf_18_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi4buf_18_auto_in_b_bits_resp),
    .auto_in_ar_ready(axi4buf_18_auto_in_ar_ready),
    .auto_in_ar_valid(axi4buf_18_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4buf_18_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4buf_18_auto_in_ar_bits_addr),
    .auto_in_ar_bits_size(axi4buf_18_auto_in_ar_bits_size),
    .auto_in_r_ready(axi4buf_18_auto_in_r_ready),
    .auto_in_r_valid(axi4buf_18_auto_in_r_valid),
    .auto_in_r_bits_id(axi4buf_18_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4buf_18_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4buf_18_auto_in_r_bits_resp),
    .auto_in_r_bits_last(axi4buf_18_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4buf_18_auto_out_aw_ready),
    .auto_out_aw_valid(axi4buf_18_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4buf_18_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4buf_18_auto_out_aw_bits_addr),
    .auto_out_w_ready(axi4buf_18_auto_out_w_ready),
    .auto_out_w_valid(axi4buf_18_auto_out_w_valid),
    .auto_out_w_bits_data(axi4buf_18_auto_out_w_bits_data),
    .auto_out_w_bits_strb(axi4buf_18_auto_out_w_bits_strb),
    .auto_out_w_bits_last(axi4buf_18_auto_out_w_bits_last),
    .auto_out_b_ready(axi4buf_18_auto_out_b_ready),
    .auto_out_b_valid(axi4buf_18_auto_out_b_valid),
    .auto_out_b_bits_id(axi4buf_18_auto_out_b_bits_id),
    .auto_out_b_bits_resp(axi4buf_18_auto_out_b_bits_resp),
    .auto_out_ar_ready(axi4buf_18_auto_out_ar_ready),
    .auto_out_ar_valid(axi4buf_18_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4buf_18_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4buf_18_auto_out_ar_bits_addr),
    .auto_out_ar_bits_size(axi4buf_18_auto_out_ar_bits_size),
    .auto_out_r_ready(axi4buf_18_auto_out_r_ready),
    .auto_out_r_valid(axi4buf_18_auto_out_r_valid),
    .auto_out_r_bits_id(axi4buf_18_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4buf_18_auto_out_r_bits_data),
    .auto_out_r_bits_resp(axi4buf_18_auto_out_r_bits_resp),
    .auto_out_r_bits_last(axi4buf_18_auto_out_r_bits_last)
  );
  AXI4Buffer axi4buf_19 ( // @[Buffer.scala 58:29]
    .clock(axi4buf_19_clock),
    .reset(axi4buf_19_reset),
    .auto_in_aw_ready(axi4buf_19_auto_in_aw_ready),
    .auto_in_aw_valid(axi4buf_19_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4buf_19_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4buf_19_auto_in_aw_bits_addr),
    .auto_in_aw_bits_size(axi4buf_19_auto_in_aw_bits_size),
    .auto_in_w_ready(axi4buf_19_auto_in_w_ready),
    .auto_in_w_valid(axi4buf_19_auto_in_w_valid),
    .auto_in_w_bits_data(axi4buf_19_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi4buf_19_auto_in_w_bits_strb),
    .auto_in_w_bits_last(axi4buf_19_auto_in_w_bits_last),
    .auto_in_b_ready(axi4buf_19_auto_in_b_ready),
    .auto_in_b_valid(axi4buf_19_auto_in_b_valid),
    .auto_in_b_bits_id(axi4buf_19_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi4buf_19_auto_in_b_bits_resp),
    .auto_in_ar_ready(axi4buf_19_auto_in_ar_ready),
    .auto_in_ar_valid(axi4buf_19_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4buf_19_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4buf_19_auto_in_ar_bits_addr),
    .auto_in_ar_bits_size(axi4buf_19_auto_in_ar_bits_size),
    .auto_in_r_ready(axi4buf_19_auto_in_r_ready),
    .auto_in_r_valid(axi4buf_19_auto_in_r_valid),
    .auto_in_r_bits_id(axi4buf_19_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4buf_19_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4buf_19_auto_in_r_bits_resp),
    .auto_in_r_bits_last(axi4buf_19_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4buf_19_auto_out_aw_ready),
    .auto_out_aw_valid(axi4buf_19_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4buf_19_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4buf_19_auto_out_aw_bits_addr),
    .auto_out_w_ready(axi4buf_19_auto_out_w_ready),
    .auto_out_w_valid(axi4buf_19_auto_out_w_valid),
    .auto_out_w_bits_data(axi4buf_19_auto_out_w_bits_data),
    .auto_out_w_bits_strb(axi4buf_19_auto_out_w_bits_strb),
    .auto_out_w_bits_last(axi4buf_19_auto_out_w_bits_last),
    .auto_out_b_ready(axi4buf_19_auto_out_b_ready),
    .auto_out_b_valid(axi4buf_19_auto_out_b_valid),
    .auto_out_b_bits_id(axi4buf_19_auto_out_b_bits_id),
    .auto_out_b_bits_resp(axi4buf_19_auto_out_b_bits_resp),
    .auto_out_ar_ready(axi4buf_19_auto_out_ar_ready),
    .auto_out_ar_valid(axi4buf_19_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4buf_19_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4buf_19_auto_out_ar_bits_addr),
    .auto_out_ar_bits_size(axi4buf_19_auto_out_ar_bits_size),
    .auto_out_r_ready(axi4buf_19_auto_out_r_ready),
    .auto_out_r_valid(axi4buf_19_auto_out_r_valid),
    .auto_out_r_bits_id(axi4buf_19_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4buf_19_auto_out_r_bits_data),
    .auto_out_r_bits_resp(axi4buf_19_auto_out_r_bits_resp),
    .auto_out_r_bits_last(axi4buf_19_auto_out_r_bits_last)
  );
  AXI4StreamBuffer buffer ( // @[Buffer.scala 29:28]
    .clock(buffer_clock),
    .reset(buffer_reset),
    .auto_in_ready(buffer_auto_in_ready),
    .auto_in_valid(buffer_auto_in_valid),
    .auto_in_bits_data(buffer_auto_in_bits_data),
    .auto_in_bits_last(buffer_auto_in_bits_last),
    .auto_out_ready(buffer_auto_out_ready),
    .auto_out_valid(buffer_auto_out_valid),
    .auto_out_bits_data(buffer_auto_out_bits_data),
    .auto_out_bits_last(buffer_auto_out_bits_last)
  );
  AXI4StreamBuffer_1 buffer_1 ( // @[Buffer.scala 29:28]
    .clock(buffer_1_clock),
    .reset(buffer_1_reset),
    .auto_in_ready(buffer_1_auto_in_ready),
    .auto_in_valid(buffer_1_auto_in_valid),
    .auto_in_bits_data(buffer_1_auto_in_bits_data),
    .auto_in_bits_last(buffer_1_auto_in_bits_last),
    .auto_out_ready(buffer_1_auto_out_ready),
    .auto_out_valid(buffer_1_auto_out_valid),
    .auto_out_bits_data(buffer_1_auto_out_bits_data),
    .auto_out_bits_last(buffer_1_auto_out_bits_last)
  );
  AXI4StreamBuffer_2 buffer_2 ( // @[Buffer.scala 29:28]
    .clock(buffer_2_clock),
    .reset(buffer_2_reset),
    .auto_in_ready(buffer_2_auto_in_ready),
    .auto_in_valid(buffer_2_auto_in_valid),
    .auto_in_bits_data(buffer_2_auto_in_bits_data),
    .auto_in_bits_last(buffer_2_auto_in_bits_last),
    .auto_out_ready(buffer_2_auto_out_ready),
    .auto_out_valid(buffer_2_auto_out_valid),
    .auto_out_bits_data(buffer_2_auto_out_bits_data),
    .auto_out_bits_last(buffer_2_auto_out_bits_last)
  );
  AXI4StreamBuffer_1 buffer_3 ( // @[Buffer.scala 29:28]
    .clock(buffer_3_clock),
    .reset(buffer_3_reset),
    .auto_in_ready(buffer_3_auto_in_ready),
    .auto_in_valid(buffer_3_auto_in_valid),
    .auto_in_bits_data(buffer_3_auto_in_bits_data),
    .auto_in_bits_last(buffer_3_auto_in_bits_last),
    .auto_out_ready(buffer_3_auto_out_ready),
    .auto_out_valid(buffer_3_auto_out_valid),
    .auto_out_bits_data(buffer_3_auto_out_bits_data),
    .auto_out_bits_last(buffer_3_auto_out_bits_last)
  );
  AXI4StreamBuffer_4 buffer_4 ( // @[Buffer.scala 29:28]
    .clock(buffer_4_clock),
    .reset(buffer_4_reset),
    .auto_in_ready(buffer_4_auto_in_ready),
    .auto_in_valid(buffer_4_auto_in_valid),
    .auto_in_bits_data(buffer_4_auto_in_bits_data),
    .auto_in_bits_last(buffer_4_auto_in_bits_last),
    .auto_out_ready(buffer_4_auto_out_ready),
    .auto_out_valid(buffer_4_auto_out_valid),
    .auto_out_bits_data(buffer_4_auto_out_bits_data),
    .auto_out_bits_last(buffer_4_auto_out_bits_last)
  );
  AXI4StreamBuffer_5 buffer_5 ( // @[Buffer.scala 29:28]
    .clock(buffer_5_clock),
    .reset(buffer_5_reset),
    .auto_in_ready(buffer_5_auto_in_ready),
    .auto_in_valid(buffer_5_auto_in_valid),
    .auto_in_bits_data(buffer_5_auto_in_bits_data),
    .auto_in_bits_last(buffer_5_auto_in_bits_last),
    .auto_out_ready(buffer_5_auto_out_ready),
    .auto_out_valid(buffer_5_auto_out_valid),
    .auto_out_bits_data(buffer_5_auto_out_bits_data),
    .auto_out_bits_last(buffer_5_auto_out_bits_last)
  );
  AXI4StreamBuffer_5 buffer_6 ( // @[Buffer.scala 29:28]
    .clock(buffer_6_clock),
    .reset(buffer_6_reset),
    .auto_in_ready(buffer_6_auto_in_ready),
    .auto_in_valid(buffer_6_auto_in_valid),
    .auto_in_bits_data(buffer_6_auto_in_bits_data),
    .auto_in_bits_last(buffer_6_auto_in_bits_last),
    .auto_out_ready(buffer_6_auto_out_ready),
    .auto_out_valid(buffer_6_auto_out_valid),
    .auto_out_bits_data(buffer_6_auto_out_bits_data),
    .auto_out_bits_last(buffer_6_auto_out_bits_last)
  );
  AXI4StreamBuffer_5 buffer_7 ( // @[Buffer.scala 29:28]
    .clock(buffer_7_clock),
    .reset(buffer_7_reset),
    .auto_in_ready(buffer_7_auto_in_ready),
    .auto_in_valid(buffer_7_auto_in_valid),
    .auto_in_bits_data(buffer_7_auto_in_bits_data),
    .auto_in_bits_last(buffer_7_auto_in_bits_last),
    .auto_out_ready(buffer_7_auto_out_ready),
    .auto_out_valid(buffer_7_auto_out_valid),
    .auto_out_bits_data(buffer_7_auto_out_bits_data),
    .auto_out_bits_last(buffer_7_auto_out_bits_last)
  );
  AXI4StreamBuffer_5 buffer_8 ( // @[Buffer.scala 29:28]
    .clock(buffer_8_clock),
    .reset(buffer_8_reset),
    .auto_in_ready(buffer_8_auto_in_ready),
    .auto_in_valid(buffer_8_auto_in_valid),
    .auto_in_bits_data(buffer_8_auto_in_bits_data),
    .auto_in_bits_last(buffer_8_auto_in_bits_last),
    .auto_out_ready(buffer_8_auto_out_ready),
    .auto_out_valid(buffer_8_auto_out_valid),
    .auto_out_bits_data(buffer_8_auto_out_bits_data),
    .auto_out_bits_last(buffer_8_auto_out_bits_last)
  );
  AXI4StreamBuffer_9 buffer_9 ( // @[Buffer.scala 29:28]
    .clock(buffer_9_clock),
    .reset(buffer_9_reset),
    .auto_in_ready(buffer_9_auto_in_ready),
    .auto_in_valid(buffer_9_auto_in_valid),
    .auto_in_bits_data(buffer_9_auto_in_bits_data),
    .auto_in_bits_last(buffer_9_auto_in_bits_last),
    .auto_out_ready(buffer_9_auto_out_ready),
    .auto_out_valid(buffer_9_auto_out_valid),
    .auto_out_bits_data(buffer_9_auto_out_bits_data),
    .auto_out_bits_last(buffer_9_auto_out_bits_last)
  );
  BundleBridgeToAXI4 converter ( // @[Node.scala 65:31]
    .auto_in_aw_ready(converter_auto_in_aw_ready),
    .auto_in_aw_valid(converter_auto_in_aw_valid),
    .auto_in_aw_bits_id(converter_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(converter_auto_in_aw_bits_addr),
    .auto_in_aw_bits_size(converter_auto_in_aw_bits_size),
    .auto_in_w_ready(converter_auto_in_w_ready),
    .auto_in_w_valid(converter_auto_in_w_valid),
    .auto_in_w_bits_data(converter_auto_in_w_bits_data),
    .auto_in_w_bits_strb(converter_auto_in_w_bits_strb),
    .auto_in_w_bits_last(converter_auto_in_w_bits_last),
    .auto_in_b_ready(converter_auto_in_b_ready),
    .auto_in_b_valid(converter_auto_in_b_valid),
    .auto_in_b_bits_resp(converter_auto_in_b_bits_resp),
    .auto_in_ar_ready(converter_auto_in_ar_ready),
    .auto_in_ar_valid(converter_auto_in_ar_valid),
    .auto_in_ar_bits_id(converter_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(converter_auto_in_ar_bits_addr),
    .auto_in_ar_bits_size(converter_auto_in_ar_bits_size),
    .auto_in_r_ready(converter_auto_in_r_ready),
    .auto_in_r_valid(converter_auto_in_r_valid),
    .auto_in_r_bits_data(converter_auto_in_r_bits_data),
    .auto_in_r_bits_resp(converter_auto_in_r_bits_resp),
    .auto_in_r_bits_last(converter_auto_in_r_bits_last),
    .auto_out_aw_ready(converter_auto_out_aw_ready),
    .auto_out_aw_valid(converter_auto_out_aw_valid),
    .auto_out_aw_bits_id(converter_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(converter_auto_out_aw_bits_addr),
    .auto_out_aw_bits_size(converter_auto_out_aw_bits_size),
    .auto_out_w_ready(converter_auto_out_w_ready),
    .auto_out_w_valid(converter_auto_out_w_valid),
    .auto_out_w_bits_data(converter_auto_out_w_bits_data),
    .auto_out_w_bits_strb(converter_auto_out_w_bits_strb),
    .auto_out_w_bits_last(converter_auto_out_w_bits_last),
    .auto_out_b_ready(converter_auto_out_b_ready),
    .auto_out_b_valid(converter_auto_out_b_valid),
    .auto_out_b_bits_resp(converter_auto_out_b_bits_resp),
    .auto_out_ar_ready(converter_auto_out_ar_ready),
    .auto_out_ar_valid(converter_auto_out_ar_valid),
    .auto_out_ar_bits_id(converter_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(converter_auto_out_ar_bits_addr),
    .auto_out_ar_bits_size(converter_auto_out_ar_bits_size),
    .auto_out_r_ready(converter_auto_out_r_ready),
    .auto_out_r_valid(converter_auto_out_r_valid),
    .auto_out_r_bits_data(converter_auto_out_r_bits_data),
    .auto_out_r_bits_resp(converter_auto_out_r_bits_resp),
    .auto_out_r_bits_last(converter_auto_out_r_bits_last)
  );
  AXI4StreamToBundleBridge converter_1 ( // @[Nodes.scala 165:31]
    .auto_in_ready(converter_1_auto_in_ready),
    .auto_in_valid(converter_1_auto_in_valid),
    .auto_in_bits_data(converter_1_auto_in_bits_data),
    .auto_in_bits_last(converter_1_auto_in_bits_last),
    .auto_out_ready(converter_1_auto_out_ready),
    .auto_out_valid(converter_1_auto_out_valid),
    .auto_out_bits_data(converter_1_auto_out_bits_data),
    .auto_out_bits_last(converter_1_auto_out_bits_last)
  );
  AXI4StreamToBundleBridge converter_2 ( // @[Nodes.scala 201:31]
    .auto_in_ready(converter_2_auto_in_ready),
    .auto_in_valid(converter_2_auto_in_valid),
    .auto_in_bits_data(converter_2_auto_in_bits_data),
    .auto_in_bits_last(converter_2_auto_in_bits_last),
    .auto_out_ready(converter_2_auto_out_ready),
    .auto_out_valid(converter_2_auto_out_valid),
    .auto_out_bits_data(converter_2_auto_out_bits_data),
    .auto_out_bits_last(converter_2_auto_out_bits_last)
  );
  assign ioMem_0_aw_ready = converter_auto_in_aw_ready; // @[Nodes.scala 624:60]
  assign ioMem_0_w_ready = converter_auto_in_w_ready; // @[Nodes.scala 624:60]
  assign ioMem_0_b_valid = converter_auto_in_b_valid; // @[Nodes.scala 624:60]
  assign ioMem_0_b_bits_id = 1'h0; // @[Nodes.scala 624:60]
  assign ioMem_0_b_bits_resp = converter_auto_in_b_bits_resp; // @[Nodes.scala 624:60]
  assign ioMem_0_ar_ready = converter_auto_in_ar_ready; // @[Nodes.scala 624:60]
  assign ioMem_0_r_valid = converter_auto_in_r_valid; // @[Nodes.scala 624:60]
  assign ioMem_0_r_bits_id = 1'h0; // @[Nodes.scala 624:60]
  assign ioMem_0_r_bits_data = converter_auto_in_r_bits_data; // @[Nodes.scala 624:60]
  assign ioMem_0_r_bits_resp = converter_auto_in_r_bits_resp; // @[Nodes.scala 624:60]
  assign ioMem_0_r_bits_last = converter_auto_in_r_bits_last; // @[Nodes.scala 624:60]
  assign outStream_0_valid = converter_1_auto_out_valid; // @[Nodes.scala 649:56]
  assign outStream_0_bits_data = converter_1_auto_out_bits_data; // @[Nodes.scala 649:56]
  assign outStream_0_bits_last = converter_1_auto_out_bits_last; // @[Nodes.scala 649:56]
  assign inStream_0_ready = converter_2_auto_in_ready; // @[Nodes.scala 624:60]
  assign int_0 = uart_int_0; // @[SpectrometerTest.scala 259:9]
  assign uTx = uart_io_txd; // @[SpectrometerTest.scala 265:9]
  assign widthAdapter_clock = clock;
  assign widthAdapter_reset = reset;
  assign widthAdapter_auto_in_valid = in_queue_auto_out_out_valid; // @[LazyModule.scala 167:31]
  assign widthAdapter_auto_in_bits_data = in_queue_auto_out_out_bits_data; // @[LazyModule.scala 167:31]
  assign widthAdapter_auto_in_bits_last = in_queue_auto_out_out_bits_last; // @[LazyModule.scala 167:31]
  assign widthAdapter_auto_out_ready = in_split_auto_stream_in_ready; // @[LazyModule.scala 167:57]
  assign in_split_clock = clock;
  assign in_split_reset = reset;
  assign in_split_auto_mem_in_aw_valid = axi4buf_auto_out_aw_valid; // @[LazyModule.scala 167:31]
  assign in_split_auto_mem_in_aw_bits_id = axi4buf_auto_out_aw_bits_id; // @[LazyModule.scala 167:31]
  assign in_split_auto_mem_in_aw_bits_addr = axi4buf_auto_out_aw_bits_addr; // @[LazyModule.scala 167:31]
  assign in_split_auto_mem_in_w_valid = axi4buf_auto_out_w_valid; // @[LazyModule.scala 167:31]
  assign in_split_auto_mem_in_w_bits_data = axi4buf_auto_out_w_bits_data; // @[LazyModule.scala 167:31]
  assign in_split_auto_mem_in_w_bits_strb = axi4buf_auto_out_w_bits_strb; // @[LazyModule.scala 167:31]
  assign in_split_auto_mem_in_b_ready = axi4buf_auto_out_b_ready; // @[LazyModule.scala 167:31]
  assign in_split_auto_mem_in_ar_valid = axi4buf_auto_out_ar_valid; // @[LazyModule.scala 167:31]
  assign in_split_auto_mem_in_ar_bits_id = axi4buf_auto_out_ar_bits_id; // @[LazyModule.scala 167:31]
  assign in_split_auto_mem_in_ar_bits_addr = axi4buf_auto_out_ar_bits_addr; // @[LazyModule.scala 167:31]
  assign in_split_auto_mem_in_ar_bits_size = axi4buf_auto_out_ar_bits_size; // @[LazyModule.scala 167:31]
  assign in_split_auto_mem_in_r_ready = axi4buf_auto_out_r_ready; // @[LazyModule.scala 167:31]
  assign in_split_auto_stream_in_valid = widthAdapter_auto_out_valid; // @[LazyModule.scala 167:57]
  assign in_split_auto_stream_in_bits_data = widthAdapter_auto_out_bits_data; // @[LazyModule.scala 167:57]
  assign in_split_auto_stream_in_bits_last = widthAdapter_auto_out_bits_last; // @[LazyModule.scala 167:57]
  assign in_split_auto_stream_out_4_ready = buffer_7_auto_in_ready; // @[LazyModule.scala 167:57]
  assign in_split_auto_stream_out_3_ready = mag_mux_0_auto_stream_in_1_ready; // @[LazyModule.scala 167:57]
  assign in_split_auto_stream_out_2_ready = fft_mux_0_auto_stream_in_1_ready; // @[LazyModule.scala 167:57]
  assign in_split_auto_stream_out_1_ready = nco_mux_0_auto_stream_in_1_ready; // @[LazyModule.scala 167:57]
  assign in_split_auto_stream_out_0_ready = plfg_mux_0_auto_stream_in_1_ready; // @[LazyModule.scala 167:57]
  assign in_queue_clock = clock;
  assign in_queue_reset = reset;
  assign in_queue_auto_out_out_ready = widthAdapter_auto_in_ready; // @[LazyModule.scala 167:31]
  assign in_queue_auto_in_in_valid = converter_2_auto_out_valid; // @[LazyModule.scala 167:31]
  assign in_queue_auto_in_in_bits_data = converter_2_auto_out_bits_data; // @[LazyModule.scala 167:31]
  assign in_queue_auto_in_in_bits_last = converter_2_auto_out_bits_last; // @[LazyModule.scala 167:31]
  assign plfg_clock = clock;
  assign plfg_reset = reset;
  assign plfg_auto_mem_in_aw_valid = axi4buf_1_auto_out_aw_valid; // @[LazyModule.scala 167:31]
  assign plfg_auto_mem_in_aw_bits_id = axi4buf_1_auto_out_aw_bits_id; // @[LazyModule.scala 167:31]
  assign plfg_auto_mem_in_aw_bits_addr = axi4buf_1_auto_out_aw_bits_addr; // @[LazyModule.scala 167:31]
  assign plfg_auto_mem_in_w_valid = axi4buf_1_auto_out_w_valid; // @[LazyModule.scala 167:31]
  assign plfg_auto_mem_in_w_bits_data = axi4buf_1_auto_out_w_bits_data; // @[LazyModule.scala 167:31]
  assign plfg_auto_mem_in_w_bits_strb = axi4buf_1_auto_out_w_bits_strb; // @[LazyModule.scala 167:31]
  assign plfg_auto_mem_in_w_bits_last = axi4buf_1_auto_out_w_bits_last; // @[LazyModule.scala 167:31]
  assign plfg_auto_mem_in_b_ready = axi4buf_1_auto_out_b_ready; // @[LazyModule.scala 167:31]
  assign plfg_auto_mem_in_ar_valid = axi4buf_1_auto_out_ar_valid; // @[LazyModule.scala 167:31]
  assign plfg_auto_mem_in_ar_bits_id = axi4buf_1_auto_out_ar_bits_id; // @[LazyModule.scala 167:31]
  assign plfg_auto_mem_in_ar_bits_addr = axi4buf_1_auto_out_ar_bits_addr; // @[LazyModule.scala 167:31]
  assign plfg_auto_mem_in_ar_bits_size = axi4buf_1_auto_out_ar_bits_size; // @[LazyModule.scala 167:31]
  assign plfg_auto_mem_in_r_ready = axi4buf_1_auto_out_r_ready; // @[LazyModule.scala 167:31]
  assign plfg_auto_stream_out_ready = plfg_split_auto_stream_in_ready; // @[LazyModule.scala 167:57]
  assign plfg_split_clock = clock;
  assign plfg_split_reset = reset;
  assign plfg_split_auto_mem_in_aw_valid = axi4buf_2_auto_out_aw_valid; // @[LazyModule.scala 167:31]
  assign plfg_split_auto_mem_in_aw_bits_id = axi4buf_2_auto_out_aw_bits_id; // @[LazyModule.scala 167:31]
  assign plfg_split_auto_mem_in_aw_bits_addr = axi4buf_2_auto_out_aw_bits_addr; // @[LazyModule.scala 167:31]
  assign plfg_split_auto_mem_in_w_valid = axi4buf_2_auto_out_w_valid; // @[LazyModule.scala 167:31]
  assign plfg_split_auto_mem_in_w_bits_data = axi4buf_2_auto_out_w_bits_data; // @[LazyModule.scala 167:31]
  assign plfg_split_auto_mem_in_w_bits_strb = axi4buf_2_auto_out_w_bits_strb; // @[LazyModule.scala 167:31]
  assign plfg_split_auto_mem_in_b_ready = axi4buf_2_auto_out_b_ready; // @[LazyModule.scala 167:31]
  assign plfg_split_auto_mem_in_ar_valid = axi4buf_2_auto_out_ar_valid; // @[LazyModule.scala 167:31]
  assign plfg_split_auto_mem_in_ar_bits_id = axi4buf_2_auto_out_ar_bits_id; // @[LazyModule.scala 167:31]
  assign plfg_split_auto_mem_in_ar_bits_addr = axi4buf_2_auto_out_ar_bits_addr; // @[LazyModule.scala 167:31]
  assign plfg_split_auto_mem_in_ar_bits_size = axi4buf_2_auto_out_ar_bits_size; // @[LazyModule.scala 167:31]
  assign plfg_split_auto_mem_in_r_ready = axi4buf_2_auto_out_r_ready; // @[LazyModule.scala 167:31]
  assign plfg_split_auto_stream_in_valid = plfg_auto_stream_out_valid; // @[LazyModule.scala 167:57]
  assign plfg_split_auto_stream_in_bits_data = plfg_auto_stream_out_bits_data; // @[LazyModule.scala 167:57]
  assign plfg_split_auto_stream_in_bits_last = plfg_auto_stream_out_bits_last; // @[LazyModule.scala 167:57]
  assign plfg_split_auto_stream_out_1_ready = plfg_mux_0_auto_stream_in_0_ready; // @[LazyModule.scala 167:57]
  assign plfg_split_auto_stream_out_0_ready = plfg_mux_1_auto_stream_in_ready; // @[LazyModule.scala 167:57]
  assign plfg_mux_0_clock = clock;
  assign plfg_mux_0_reset = reset;
  assign plfg_mux_0_auto_register_in_aw_valid = axi4buf_3_auto_out_aw_valid; // @[LazyModule.scala 167:31]
  assign plfg_mux_0_auto_register_in_aw_bits_id = axi4buf_3_auto_out_aw_bits_id; // @[LazyModule.scala 167:31]
  assign plfg_mux_0_auto_register_in_aw_bits_addr = axi4buf_3_auto_out_aw_bits_addr; // @[LazyModule.scala 167:31]
  assign plfg_mux_0_auto_register_in_w_valid = axi4buf_3_auto_out_w_valid; // @[LazyModule.scala 167:31]
  assign plfg_mux_0_auto_register_in_w_bits_data = axi4buf_3_auto_out_w_bits_data; // @[LazyModule.scala 167:31]
  assign plfg_mux_0_auto_register_in_w_bits_strb = axi4buf_3_auto_out_w_bits_strb; // @[LazyModule.scala 167:31]
  assign plfg_mux_0_auto_register_in_b_ready = axi4buf_3_auto_out_b_ready; // @[LazyModule.scala 167:31]
  assign plfg_mux_0_auto_register_in_ar_valid = axi4buf_3_auto_out_ar_valid; // @[LazyModule.scala 167:31]
  assign plfg_mux_0_auto_register_in_ar_bits_id = axi4buf_3_auto_out_ar_bits_id; // @[LazyModule.scala 167:31]
  assign plfg_mux_0_auto_register_in_ar_bits_addr = axi4buf_3_auto_out_ar_bits_addr; // @[LazyModule.scala 167:31]
  assign plfg_mux_0_auto_register_in_ar_bits_size = axi4buf_3_auto_out_ar_bits_size; // @[LazyModule.scala 167:31]
  assign plfg_mux_0_auto_register_in_r_ready = axi4buf_3_auto_out_r_ready; // @[LazyModule.scala 167:31]
  assign plfg_mux_0_auto_stream_in_2_valid = uRx_split_auto_stream_out_0_valid; // @[LazyModule.scala 167:31]
  assign plfg_mux_0_auto_stream_in_2_bits_data = uRx_split_auto_stream_out_0_bits_data; // @[LazyModule.scala 167:31]
  assign plfg_mux_0_auto_stream_in_2_bits_last = uRx_split_auto_stream_out_0_bits_last; // @[LazyModule.scala 167:31]
  assign plfg_mux_0_auto_stream_in_1_valid = in_split_auto_stream_out_0_valid; // @[LazyModule.scala 167:57]
  assign plfg_mux_0_auto_stream_in_1_bits_data = in_split_auto_stream_out_0_bits_data; // @[LazyModule.scala 167:57]
  assign plfg_mux_0_auto_stream_in_1_bits_last = in_split_auto_stream_out_0_bits_last; // @[LazyModule.scala 167:57]
  assign plfg_mux_0_auto_stream_in_0_valid = plfg_split_auto_stream_out_1_valid; // @[LazyModule.scala 167:57]
  assign plfg_mux_0_auto_stream_in_0_bits_data = plfg_split_auto_stream_out_1_bits_data; // @[LazyModule.scala 167:57]
  assign plfg_mux_0_auto_stream_in_0_bits_last = plfg_split_auto_stream_out_1_bits_last; // @[LazyModule.scala 167:57]
  assign plfg_mux_0_auto_stream_out_0_ready = nco_auto_freq_in_ready; // @[LazyModule.scala 167:57]
  assign plfg_mux_1_clock = clock;
  assign plfg_mux_1_reset = reset;
  assign plfg_mux_1_auto_register_in_aw_valid = axi4buf_4_auto_out_aw_valid; // @[LazyModule.scala 167:31]
  assign plfg_mux_1_auto_register_in_aw_bits_id = axi4buf_4_auto_out_aw_bits_id; // @[LazyModule.scala 167:31]
  assign plfg_mux_1_auto_register_in_aw_bits_addr = axi4buf_4_auto_out_aw_bits_addr; // @[LazyModule.scala 167:31]
  assign plfg_mux_1_auto_register_in_w_valid = axi4buf_4_auto_out_w_valid; // @[LazyModule.scala 167:31]
  assign plfg_mux_1_auto_register_in_w_bits_data = axi4buf_4_auto_out_w_bits_data; // @[LazyModule.scala 167:31]
  assign plfg_mux_1_auto_register_in_w_bits_strb = axi4buf_4_auto_out_w_bits_strb; // @[LazyModule.scala 167:31]
  assign plfg_mux_1_auto_register_in_b_ready = axi4buf_4_auto_out_b_ready; // @[LazyModule.scala 167:31]
  assign plfg_mux_1_auto_register_in_ar_valid = axi4buf_4_auto_out_ar_valid; // @[LazyModule.scala 167:31]
  assign plfg_mux_1_auto_register_in_ar_bits_id = axi4buf_4_auto_out_ar_bits_id; // @[LazyModule.scala 167:31]
  assign plfg_mux_1_auto_register_in_ar_bits_addr = axi4buf_4_auto_out_ar_bits_addr; // @[LazyModule.scala 167:31]
  assign plfg_mux_1_auto_register_in_ar_bits_size = axi4buf_4_auto_out_ar_bits_size; // @[LazyModule.scala 167:31]
  assign plfg_mux_1_auto_register_in_r_ready = axi4buf_4_auto_out_r_ready; // @[LazyModule.scala 167:31]
  assign plfg_mux_1_auto_stream_in_valid = plfg_split_auto_stream_out_0_valid; // @[LazyModule.scala 167:57]
  assign plfg_mux_1_auto_stream_in_bits_data = plfg_split_auto_stream_out_0_bits_data; // @[LazyModule.scala 167:57]
  assign plfg_mux_1_auto_stream_in_bits_last = plfg_split_auto_stream_out_0_bits_last; // @[LazyModule.scala 167:57]
  assign plfg_mux_1_auto_stream_out_1_ready = buffer_6_auto_in_ready; // @[LazyModule.scala 167:57]
  assign nco_clock = clock;
  assign nco_reset = reset;
  assign nco_auto_stream_out_ready = nco_split_auto_stream_in_ready; // @[LazyModule.scala 167:57]
  assign nco_auto_freq_in_valid = plfg_mux_0_auto_stream_out_0_valid; // @[LazyModule.scala 167:57]
  assign nco_auto_freq_in_bits_data = plfg_mux_0_auto_stream_out_0_bits_data; // @[LazyModule.scala 167:57]
  assign nco_auto_freq_in_bits_last = plfg_mux_0_auto_stream_out_0_bits_last; // @[LazyModule.scala 167:57]
  assign nco_split_clock = clock;
  assign nco_split_reset = reset;
  assign nco_split_auto_mem_in_aw_valid = axi4buf_6_auto_out_aw_valid; // @[LazyModule.scala 167:31]
  assign nco_split_auto_mem_in_aw_bits_id = axi4buf_6_auto_out_aw_bits_id; // @[LazyModule.scala 167:31]
  assign nco_split_auto_mem_in_aw_bits_addr = axi4buf_6_auto_out_aw_bits_addr; // @[LazyModule.scala 167:31]
  assign nco_split_auto_mem_in_w_valid = axi4buf_6_auto_out_w_valid; // @[LazyModule.scala 167:31]
  assign nco_split_auto_mem_in_w_bits_data = axi4buf_6_auto_out_w_bits_data; // @[LazyModule.scala 167:31]
  assign nco_split_auto_mem_in_w_bits_strb = axi4buf_6_auto_out_w_bits_strb; // @[LazyModule.scala 167:31]
  assign nco_split_auto_mem_in_b_ready = axi4buf_6_auto_out_b_ready; // @[LazyModule.scala 167:31]
  assign nco_split_auto_mem_in_ar_valid = axi4buf_6_auto_out_ar_valid; // @[LazyModule.scala 167:31]
  assign nco_split_auto_mem_in_ar_bits_id = axi4buf_6_auto_out_ar_bits_id; // @[LazyModule.scala 167:31]
  assign nco_split_auto_mem_in_ar_bits_addr = axi4buf_6_auto_out_ar_bits_addr; // @[LazyModule.scala 167:31]
  assign nco_split_auto_mem_in_ar_bits_size = axi4buf_6_auto_out_ar_bits_size; // @[LazyModule.scala 167:31]
  assign nco_split_auto_mem_in_r_ready = axi4buf_6_auto_out_r_ready; // @[LazyModule.scala 167:31]
  assign nco_split_auto_stream_in_valid = nco_auto_stream_out_valid; // @[LazyModule.scala 167:57]
  assign nco_split_auto_stream_in_bits_data = nco_auto_stream_out_bits_data; // @[LazyModule.scala 167:57]
  assign nco_split_auto_stream_in_bits_last = nco_auto_stream_out_bits_last; // @[LazyModule.scala 167:57]
  assign nco_split_auto_stream_out_1_ready = nco_mux_0_auto_stream_in_0_ready; // @[LazyModule.scala 167:57]
  assign nco_split_auto_stream_out_0_ready = nco_mux_1_auto_stream_in_ready; // @[LazyModule.scala 167:57]
  assign nco_mux_0_clock = clock;
  assign nco_mux_0_reset = reset;
  assign nco_mux_0_auto_register_in_aw_valid = axi4buf_7_auto_out_aw_valid; // @[LazyModule.scala 167:31]
  assign nco_mux_0_auto_register_in_aw_bits_id = axi4buf_7_auto_out_aw_bits_id; // @[LazyModule.scala 167:31]
  assign nco_mux_0_auto_register_in_aw_bits_addr = axi4buf_7_auto_out_aw_bits_addr; // @[LazyModule.scala 167:31]
  assign nco_mux_0_auto_register_in_w_valid = axi4buf_7_auto_out_w_valid; // @[LazyModule.scala 167:31]
  assign nco_mux_0_auto_register_in_w_bits_data = axi4buf_7_auto_out_w_bits_data; // @[LazyModule.scala 167:31]
  assign nco_mux_0_auto_register_in_w_bits_strb = axi4buf_7_auto_out_w_bits_strb; // @[LazyModule.scala 167:31]
  assign nco_mux_0_auto_register_in_b_ready = axi4buf_7_auto_out_b_ready; // @[LazyModule.scala 167:31]
  assign nco_mux_0_auto_register_in_ar_valid = axi4buf_7_auto_out_ar_valid; // @[LazyModule.scala 167:31]
  assign nco_mux_0_auto_register_in_ar_bits_id = axi4buf_7_auto_out_ar_bits_id; // @[LazyModule.scala 167:31]
  assign nco_mux_0_auto_register_in_ar_bits_addr = axi4buf_7_auto_out_ar_bits_addr; // @[LazyModule.scala 167:31]
  assign nco_mux_0_auto_register_in_ar_bits_size = axi4buf_7_auto_out_ar_bits_size; // @[LazyModule.scala 167:31]
  assign nco_mux_0_auto_register_in_r_ready = axi4buf_7_auto_out_r_ready; // @[LazyModule.scala 167:31]
  assign nco_mux_0_auto_stream_in_2_valid = uRx_split_auto_stream_out_1_valid; // @[LazyModule.scala 167:31]
  assign nco_mux_0_auto_stream_in_2_bits_data = uRx_split_auto_stream_out_1_bits_data; // @[LazyModule.scala 167:31]
  assign nco_mux_0_auto_stream_in_2_bits_last = uRx_split_auto_stream_out_1_bits_last; // @[LazyModule.scala 167:31]
  assign nco_mux_0_auto_stream_in_1_valid = in_split_auto_stream_out_1_valid; // @[LazyModule.scala 167:57]
  assign nco_mux_0_auto_stream_in_1_bits_data = in_split_auto_stream_out_1_bits_data; // @[LazyModule.scala 167:57]
  assign nco_mux_0_auto_stream_in_1_bits_last = in_split_auto_stream_out_1_bits_last; // @[LazyModule.scala 167:57]
  assign nco_mux_0_auto_stream_in_0_valid = nco_split_auto_stream_out_1_valid; // @[LazyModule.scala 167:57]
  assign nco_mux_0_auto_stream_in_0_bits_data = nco_split_auto_stream_out_1_bits_data; // @[LazyModule.scala 167:57]
  assign nco_mux_0_auto_stream_in_0_bits_last = nco_split_auto_stream_out_1_bits_last; // @[LazyModule.scala 167:57]
  assign nco_mux_0_auto_stream_out_0_ready = buffer_auto_in_ready; // @[LazyModule.scala 167:57]
  assign nco_mux_1_clock = clock;
  assign nco_mux_1_reset = reset;
  assign nco_mux_1_auto_register_in_aw_valid = axi4buf_8_auto_out_aw_valid; // @[LazyModule.scala 167:31]
  assign nco_mux_1_auto_register_in_aw_bits_id = axi4buf_8_auto_out_aw_bits_id; // @[LazyModule.scala 167:31]
  assign nco_mux_1_auto_register_in_aw_bits_addr = axi4buf_8_auto_out_aw_bits_addr; // @[LazyModule.scala 167:31]
  assign nco_mux_1_auto_register_in_w_valid = axi4buf_8_auto_out_w_valid; // @[LazyModule.scala 167:31]
  assign nco_mux_1_auto_register_in_w_bits_data = axi4buf_8_auto_out_w_bits_data; // @[LazyModule.scala 167:31]
  assign nco_mux_1_auto_register_in_w_bits_strb = axi4buf_8_auto_out_w_bits_strb; // @[LazyModule.scala 167:31]
  assign nco_mux_1_auto_register_in_b_ready = axi4buf_8_auto_out_b_ready; // @[LazyModule.scala 167:31]
  assign nco_mux_1_auto_register_in_ar_valid = axi4buf_8_auto_out_ar_valid; // @[LazyModule.scala 167:31]
  assign nco_mux_1_auto_register_in_ar_bits_id = axi4buf_8_auto_out_ar_bits_id; // @[LazyModule.scala 167:31]
  assign nco_mux_1_auto_register_in_ar_bits_addr = axi4buf_8_auto_out_ar_bits_addr; // @[LazyModule.scala 167:31]
  assign nco_mux_1_auto_register_in_ar_bits_size = axi4buf_8_auto_out_ar_bits_size; // @[LazyModule.scala 167:31]
  assign nco_mux_1_auto_register_in_r_ready = axi4buf_8_auto_out_r_ready; // @[LazyModule.scala 167:31]
  assign nco_mux_1_auto_stream_in_valid = nco_split_auto_stream_out_0_valid; // @[LazyModule.scala 167:57]
  assign nco_mux_1_auto_stream_in_bits_data = nco_split_auto_stream_out_0_bits_data; // @[LazyModule.scala 167:57]
  assign nco_mux_1_auto_stream_in_bits_last = nco_split_auto_stream_out_0_bits_last; // @[LazyModule.scala 167:57]
  assign nco_mux_1_auto_stream_out_1_ready = buffer_5_auto_in_ready; // @[LazyModule.scala 167:57]
  assign fft_clock = clock;
  assign fft_reset = reset;
  assign fft_auto_mem_in_aw_valid = axi4buf_9_auto_out_aw_valid; // @[LazyModule.scala 167:31]
  assign fft_auto_mem_in_aw_bits_id = axi4buf_9_auto_out_aw_bits_id; // @[LazyModule.scala 167:31]
  assign fft_auto_mem_in_aw_bits_addr = axi4buf_9_auto_out_aw_bits_addr; // @[LazyModule.scala 167:31]
  assign fft_auto_mem_in_w_valid = axi4buf_9_auto_out_w_valid; // @[LazyModule.scala 167:31]
  assign fft_auto_mem_in_w_bits_data = axi4buf_9_auto_out_w_bits_data; // @[LazyModule.scala 167:31]
  assign fft_auto_mem_in_w_bits_strb = axi4buf_9_auto_out_w_bits_strb; // @[LazyModule.scala 167:31]
  assign fft_auto_mem_in_b_ready = axi4buf_9_auto_out_b_ready; // @[LazyModule.scala 167:31]
  assign fft_auto_mem_in_ar_valid = axi4buf_9_auto_out_ar_valid; // @[LazyModule.scala 167:31]
  assign fft_auto_mem_in_ar_bits_id = axi4buf_9_auto_out_ar_bits_id; // @[LazyModule.scala 167:31]
  assign fft_auto_mem_in_ar_bits_addr = axi4buf_9_auto_out_ar_bits_addr; // @[LazyModule.scala 167:31]
  assign fft_auto_mem_in_ar_bits_size = axi4buf_9_auto_out_ar_bits_size; // @[LazyModule.scala 167:31]
  assign fft_auto_mem_in_r_ready = axi4buf_9_auto_out_r_ready; // @[LazyModule.scala 167:31]
  assign fft_auto_stream_in_valid = buffer_auto_out_valid; // @[LazyModule.scala 167:31]
  assign fft_auto_stream_in_bits_data = buffer_auto_out_bits_data; // @[LazyModule.scala 167:31]
  assign fft_auto_stream_in_bits_last = buffer_auto_out_bits_last; // @[LazyModule.scala 167:31]
  assign fft_auto_stream_out_ready = fft_split_auto_stream_in_ready; // @[LazyModule.scala 167:57]
  assign fft_split_clock = clock;
  assign fft_split_reset = reset;
  assign fft_split_auto_mem_in_aw_valid = axi4buf_10_auto_out_aw_valid; // @[LazyModule.scala 167:31]
  assign fft_split_auto_mem_in_aw_bits_id = axi4buf_10_auto_out_aw_bits_id; // @[LazyModule.scala 167:31]
  assign fft_split_auto_mem_in_aw_bits_addr = axi4buf_10_auto_out_aw_bits_addr; // @[LazyModule.scala 167:31]
  assign fft_split_auto_mem_in_w_valid = axi4buf_10_auto_out_w_valid; // @[LazyModule.scala 167:31]
  assign fft_split_auto_mem_in_w_bits_data = axi4buf_10_auto_out_w_bits_data; // @[LazyModule.scala 167:31]
  assign fft_split_auto_mem_in_w_bits_strb = axi4buf_10_auto_out_w_bits_strb; // @[LazyModule.scala 167:31]
  assign fft_split_auto_mem_in_b_ready = axi4buf_10_auto_out_b_ready; // @[LazyModule.scala 167:31]
  assign fft_split_auto_mem_in_ar_valid = axi4buf_10_auto_out_ar_valid; // @[LazyModule.scala 167:31]
  assign fft_split_auto_mem_in_ar_bits_id = axi4buf_10_auto_out_ar_bits_id; // @[LazyModule.scala 167:31]
  assign fft_split_auto_mem_in_ar_bits_addr = axi4buf_10_auto_out_ar_bits_addr; // @[LazyModule.scala 167:31]
  assign fft_split_auto_mem_in_ar_bits_size = axi4buf_10_auto_out_ar_bits_size; // @[LazyModule.scala 167:31]
  assign fft_split_auto_mem_in_r_ready = axi4buf_10_auto_out_r_ready; // @[LazyModule.scala 167:31]
  assign fft_split_auto_stream_in_valid = fft_auto_stream_out_valid; // @[LazyModule.scala 167:57]
  assign fft_split_auto_stream_in_bits_data = fft_auto_stream_out_bits_data; // @[LazyModule.scala 167:57]
  assign fft_split_auto_stream_in_bits_last = fft_auto_stream_out_bits_last; // @[LazyModule.scala 167:57]
  assign fft_split_auto_stream_out_1_ready = fft_mux_0_auto_stream_in_0_ready; // @[LazyModule.scala 167:57]
  assign fft_split_auto_stream_out_0_ready = fft_mux_1_auto_stream_in_ready; // @[LazyModule.scala 167:57]
  assign fft_mux_0_clock = clock;
  assign fft_mux_0_reset = reset;
  assign fft_mux_0_auto_register_in_aw_valid = axi4buf_11_auto_out_aw_valid; // @[LazyModule.scala 167:31]
  assign fft_mux_0_auto_register_in_aw_bits_id = axi4buf_11_auto_out_aw_bits_id; // @[LazyModule.scala 167:31]
  assign fft_mux_0_auto_register_in_aw_bits_addr = axi4buf_11_auto_out_aw_bits_addr; // @[LazyModule.scala 167:31]
  assign fft_mux_0_auto_register_in_w_valid = axi4buf_11_auto_out_w_valid; // @[LazyModule.scala 167:31]
  assign fft_mux_0_auto_register_in_w_bits_data = axi4buf_11_auto_out_w_bits_data; // @[LazyModule.scala 167:31]
  assign fft_mux_0_auto_register_in_w_bits_strb = axi4buf_11_auto_out_w_bits_strb; // @[LazyModule.scala 167:31]
  assign fft_mux_0_auto_register_in_b_ready = axi4buf_11_auto_out_b_ready; // @[LazyModule.scala 167:31]
  assign fft_mux_0_auto_register_in_ar_valid = axi4buf_11_auto_out_ar_valid; // @[LazyModule.scala 167:31]
  assign fft_mux_0_auto_register_in_ar_bits_id = axi4buf_11_auto_out_ar_bits_id; // @[LazyModule.scala 167:31]
  assign fft_mux_0_auto_register_in_ar_bits_addr = axi4buf_11_auto_out_ar_bits_addr; // @[LazyModule.scala 167:31]
  assign fft_mux_0_auto_register_in_ar_bits_size = axi4buf_11_auto_out_ar_bits_size; // @[LazyModule.scala 167:31]
  assign fft_mux_0_auto_register_in_r_ready = axi4buf_11_auto_out_r_ready; // @[LazyModule.scala 167:31]
  assign fft_mux_0_auto_stream_in_2_valid = uRx_split_auto_stream_out_2_valid; // @[LazyModule.scala 167:31]
  assign fft_mux_0_auto_stream_in_2_bits_data = uRx_split_auto_stream_out_2_bits_data; // @[LazyModule.scala 167:31]
  assign fft_mux_0_auto_stream_in_2_bits_last = uRx_split_auto_stream_out_2_bits_last; // @[LazyModule.scala 167:31]
  assign fft_mux_0_auto_stream_in_1_valid = in_split_auto_stream_out_2_valid; // @[LazyModule.scala 167:57]
  assign fft_mux_0_auto_stream_in_1_bits_data = in_split_auto_stream_out_2_bits_data; // @[LazyModule.scala 167:57]
  assign fft_mux_0_auto_stream_in_1_bits_last = in_split_auto_stream_out_2_bits_last; // @[LazyModule.scala 167:57]
  assign fft_mux_0_auto_stream_in_0_valid = fft_split_auto_stream_out_1_valid; // @[LazyModule.scala 167:57]
  assign fft_mux_0_auto_stream_in_0_bits_data = fft_split_auto_stream_out_1_bits_data; // @[LazyModule.scala 167:57]
  assign fft_mux_0_auto_stream_in_0_bits_last = fft_split_auto_stream_out_1_bits_last; // @[LazyModule.scala 167:57]
  assign fft_mux_0_auto_stream_out_0_ready = buffer_1_auto_in_ready; // @[LazyModule.scala 167:57]
  assign fft_mux_1_clock = clock;
  assign fft_mux_1_reset = reset;
  assign fft_mux_1_auto_register_in_aw_valid = axi4buf_12_auto_out_aw_valid; // @[LazyModule.scala 167:31]
  assign fft_mux_1_auto_register_in_aw_bits_id = axi4buf_12_auto_out_aw_bits_id; // @[LazyModule.scala 167:31]
  assign fft_mux_1_auto_register_in_aw_bits_addr = axi4buf_12_auto_out_aw_bits_addr; // @[LazyModule.scala 167:31]
  assign fft_mux_1_auto_register_in_w_valid = axi4buf_12_auto_out_w_valid; // @[LazyModule.scala 167:31]
  assign fft_mux_1_auto_register_in_w_bits_data = axi4buf_12_auto_out_w_bits_data; // @[LazyModule.scala 167:31]
  assign fft_mux_1_auto_register_in_w_bits_strb = axi4buf_12_auto_out_w_bits_strb; // @[LazyModule.scala 167:31]
  assign fft_mux_1_auto_register_in_b_ready = axi4buf_12_auto_out_b_ready; // @[LazyModule.scala 167:31]
  assign fft_mux_1_auto_register_in_ar_valid = axi4buf_12_auto_out_ar_valid; // @[LazyModule.scala 167:31]
  assign fft_mux_1_auto_register_in_ar_bits_id = axi4buf_12_auto_out_ar_bits_id; // @[LazyModule.scala 167:31]
  assign fft_mux_1_auto_register_in_ar_bits_addr = axi4buf_12_auto_out_ar_bits_addr; // @[LazyModule.scala 167:31]
  assign fft_mux_1_auto_register_in_ar_bits_size = axi4buf_12_auto_out_ar_bits_size; // @[LazyModule.scala 167:31]
  assign fft_mux_1_auto_register_in_r_ready = axi4buf_12_auto_out_r_ready; // @[LazyModule.scala 167:31]
  assign fft_mux_1_auto_stream_in_valid = fft_split_auto_stream_out_0_valid; // @[LazyModule.scala 167:57]
  assign fft_mux_1_auto_stream_in_bits_data = fft_split_auto_stream_out_0_bits_data; // @[LazyModule.scala 167:57]
  assign fft_mux_1_auto_stream_in_bits_last = fft_split_auto_stream_out_0_bits_last; // @[LazyModule.scala 167:57]
  assign fft_mux_1_auto_stream_out_1_ready = buffer_4_auto_in_ready; // @[LazyModule.scala 167:57]
  assign mag_clock = clock;
  assign mag_reset = reset;
  assign mag_auto_mem_in_aw_valid = axi4buf_13_auto_out_aw_valid; // @[LazyModule.scala 167:31]
  assign mag_auto_mem_in_aw_bits_id = axi4buf_13_auto_out_aw_bits_id; // @[LazyModule.scala 167:31]
  assign mag_auto_mem_in_aw_bits_addr = axi4buf_13_auto_out_aw_bits_addr; // @[LazyModule.scala 167:31]
  assign mag_auto_mem_in_w_valid = axi4buf_13_auto_out_w_valid; // @[LazyModule.scala 167:31]
  assign mag_auto_mem_in_w_bits_data = axi4buf_13_auto_out_w_bits_data; // @[LazyModule.scala 167:31]
  assign mag_auto_mem_in_w_bits_strb = axi4buf_13_auto_out_w_bits_strb; // @[LazyModule.scala 167:31]
  assign mag_auto_mem_in_b_ready = axi4buf_13_auto_out_b_ready; // @[LazyModule.scala 167:31]
  assign mag_auto_mem_in_ar_valid = axi4buf_13_auto_out_ar_valid; // @[LazyModule.scala 167:31]
  assign mag_auto_mem_in_ar_bits_id = axi4buf_13_auto_out_ar_bits_id; // @[LazyModule.scala 167:31]
  assign mag_auto_mem_in_ar_bits_addr = axi4buf_13_auto_out_ar_bits_addr; // @[LazyModule.scala 167:31]
  assign mag_auto_mem_in_ar_bits_size = axi4buf_13_auto_out_ar_bits_size; // @[LazyModule.scala 167:31]
  assign mag_auto_mem_in_r_ready = axi4buf_13_auto_out_r_ready; // @[LazyModule.scala 167:31]
  assign mag_auto_stream_in_valid = buffer_1_auto_out_valid; // @[LazyModule.scala 167:31]
  assign mag_auto_stream_in_bits_data = buffer_1_auto_out_bits_data; // @[LazyModule.scala 167:31]
  assign mag_auto_stream_in_bits_last = buffer_1_auto_out_bits_last; // @[LazyModule.scala 167:31]
  assign mag_auto_stream_out_ready = mag_split_auto_stream_in_ready; // @[LazyModule.scala 167:57]
  assign mag_split_clock = clock;
  assign mag_split_reset = reset;
  assign mag_split_auto_mem_in_aw_valid = axi4buf_14_auto_out_aw_valid; // @[LazyModule.scala 167:31]
  assign mag_split_auto_mem_in_aw_bits_id = axi4buf_14_auto_out_aw_bits_id; // @[LazyModule.scala 167:31]
  assign mag_split_auto_mem_in_aw_bits_addr = axi4buf_14_auto_out_aw_bits_addr; // @[LazyModule.scala 167:31]
  assign mag_split_auto_mem_in_w_valid = axi4buf_14_auto_out_w_valid; // @[LazyModule.scala 167:31]
  assign mag_split_auto_mem_in_w_bits_data = axi4buf_14_auto_out_w_bits_data; // @[LazyModule.scala 167:31]
  assign mag_split_auto_mem_in_w_bits_strb = axi4buf_14_auto_out_w_bits_strb; // @[LazyModule.scala 167:31]
  assign mag_split_auto_mem_in_b_ready = axi4buf_14_auto_out_b_ready; // @[LazyModule.scala 167:31]
  assign mag_split_auto_mem_in_ar_valid = axi4buf_14_auto_out_ar_valid; // @[LazyModule.scala 167:31]
  assign mag_split_auto_mem_in_ar_bits_id = axi4buf_14_auto_out_ar_bits_id; // @[LazyModule.scala 167:31]
  assign mag_split_auto_mem_in_ar_bits_addr = axi4buf_14_auto_out_ar_bits_addr; // @[LazyModule.scala 167:31]
  assign mag_split_auto_mem_in_ar_bits_size = axi4buf_14_auto_out_ar_bits_size; // @[LazyModule.scala 167:31]
  assign mag_split_auto_mem_in_r_ready = axi4buf_14_auto_out_r_ready; // @[LazyModule.scala 167:31]
  assign mag_split_auto_stream_in_valid = mag_auto_stream_out_valid; // @[LazyModule.scala 167:57]
  assign mag_split_auto_stream_in_bits_data = mag_auto_stream_out_bits_data; // @[LazyModule.scala 167:57]
  assign mag_split_auto_stream_in_bits_last = mag_auto_stream_out_bits_last; // @[LazyModule.scala 167:57]
  assign mag_split_auto_stream_out_1_ready = mag_mux_0_auto_stream_in_0_ready; // @[LazyModule.scala 167:57]
  assign mag_split_auto_stream_out_0_ready = mag_mux_1_auto_stream_in_ready; // @[LazyModule.scala 167:57]
  assign mag_mux_0_clock = clock;
  assign mag_mux_0_reset = reset;
  assign mag_mux_0_auto_register_in_aw_valid = axi4buf_15_auto_out_aw_valid; // @[LazyModule.scala 167:31]
  assign mag_mux_0_auto_register_in_aw_bits_id = axi4buf_15_auto_out_aw_bits_id; // @[LazyModule.scala 167:31]
  assign mag_mux_0_auto_register_in_aw_bits_addr = axi4buf_15_auto_out_aw_bits_addr; // @[LazyModule.scala 167:31]
  assign mag_mux_0_auto_register_in_w_valid = axi4buf_15_auto_out_w_valid; // @[LazyModule.scala 167:31]
  assign mag_mux_0_auto_register_in_w_bits_data = axi4buf_15_auto_out_w_bits_data; // @[LazyModule.scala 167:31]
  assign mag_mux_0_auto_register_in_w_bits_strb = axi4buf_15_auto_out_w_bits_strb; // @[LazyModule.scala 167:31]
  assign mag_mux_0_auto_register_in_b_ready = axi4buf_15_auto_out_b_ready; // @[LazyModule.scala 167:31]
  assign mag_mux_0_auto_register_in_ar_valid = axi4buf_15_auto_out_ar_valid; // @[LazyModule.scala 167:31]
  assign mag_mux_0_auto_register_in_ar_bits_id = axi4buf_15_auto_out_ar_bits_id; // @[LazyModule.scala 167:31]
  assign mag_mux_0_auto_register_in_ar_bits_addr = axi4buf_15_auto_out_ar_bits_addr; // @[LazyModule.scala 167:31]
  assign mag_mux_0_auto_register_in_ar_bits_size = axi4buf_15_auto_out_ar_bits_size; // @[LazyModule.scala 167:31]
  assign mag_mux_0_auto_register_in_r_ready = axi4buf_15_auto_out_r_ready; // @[LazyModule.scala 167:31]
  assign mag_mux_0_auto_stream_in_2_valid = uRx_split_auto_stream_out_3_valid; // @[LazyModule.scala 167:31]
  assign mag_mux_0_auto_stream_in_2_bits_data = uRx_split_auto_stream_out_3_bits_data; // @[LazyModule.scala 167:31]
  assign mag_mux_0_auto_stream_in_2_bits_last = uRx_split_auto_stream_out_3_bits_last; // @[LazyModule.scala 167:31]
  assign mag_mux_0_auto_stream_in_1_valid = in_split_auto_stream_out_3_valid; // @[LazyModule.scala 167:57]
  assign mag_mux_0_auto_stream_in_1_bits_data = in_split_auto_stream_out_3_bits_data; // @[LazyModule.scala 167:57]
  assign mag_mux_0_auto_stream_in_1_bits_last = in_split_auto_stream_out_3_bits_last; // @[LazyModule.scala 167:57]
  assign mag_mux_0_auto_stream_in_0_valid = mag_split_auto_stream_out_1_valid; // @[LazyModule.scala 167:57]
  assign mag_mux_0_auto_stream_in_0_bits_data = mag_split_auto_stream_out_1_bits_data; // @[LazyModule.scala 167:57]
  assign mag_mux_0_auto_stream_in_0_bits_last = mag_split_auto_stream_out_1_bits_last; // @[LazyModule.scala 167:57]
  assign mag_mux_0_auto_stream_out_0_ready = buffer_2_auto_in_ready; // @[LazyModule.scala 167:57]
  assign mag_mux_1_clock = clock;
  assign mag_mux_1_reset = reset;
  assign mag_mux_1_auto_register_in_aw_valid = axi4buf_16_auto_out_aw_valid; // @[LazyModule.scala 167:31]
  assign mag_mux_1_auto_register_in_aw_bits_id = axi4buf_16_auto_out_aw_bits_id; // @[LazyModule.scala 167:31]
  assign mag_mux_1_auto_register_in_aw_bits_addr = axi4buf_16_auto_out_aw_bits_addr; // @[LazyModule.scala 167:31]
  assign mag_mux_1_auto_register_in_w_valid = axi4buf_16_auto_out_w_valid; // @[LazyModule.scala 167:31]
  assign mag_mux_1_auto_register_in_w_bits_data = axi4buf_16_auto_out_w_bits_data; // @[LazyModule.scala 167:31]
  assign mag_mux_1_auto_register_in_w_bits_strb = axi4buf_16_auto_out_w_bits_strb; // @[LazyModule.scala 167:31]
  assign mag_mux_1_auto_register_in_b_ready = axi4buf_16_auto_out_b_ready; // @[LazyModule.scala 167:31]
  assign mag_mux_1_auto_register_in_ar_valid = axi4buf_16_auto_out_ar_valid; // @[LazyModule.scala 167:31]
  assign mag_mux_1_auto_register_in_ar_bits_id = axi4buf_16_auto_out_ar_bits_id; // @[LazyModule.scala 167:31]
  assign mag_mux_1_auto_register_in_ar_bits_addr = axi4buf_16_auto_out_ar_bits_addr; // @[LazyModule.scala 167:31]
  assign mag_mux_1_auto_register_in_ar_bits_size = axi4buf_16_auto_out_ar_bits_size; // @[LazyModule.scala 167:31]
  assign mag_mux_1_auto_register_in_r_ready = axi4buf_16_auto_out_r_ready; // @[LazyModule.scala 167:31]
  assign mag_mux_1_auto_stream_in_valid = mag_split_auto_stream_out_0_valid; // @[LazyModule.scala 167:57]
  assign mag_mux_1_auto_stream_in_bits_data = mag_split_auto_stream_out_0_bits_data; // @[LazyModule.scala 167:57]
  assign mag_mux_1_auto_stream_in_bits_last = mag_split_auto_stream_out_0_bits_last; // @[LazyModule.scala 167:57]
  assign mag_mux_1_auto_stream_out_1_ready = buffer_3_auto_in_ready; // @[LazyModule.scala 167:57]
  assign acc_clock = clock;
  assign acc_reset = reset;
  assign acc_auto_bus_in_aw_valid = bus_auto_out_20_aw_valid; // @[LazyModule.scala 167:31]
  assign acc_auto_bus_in_aw_bits_id = bus_auto_out_20_aw_bits_id; // @[LazyModule.scala 167:31]
  assign acc_auto_bus_in_aw_bits_addr = bus_auto_out_20_aw_bits_addr; // @[LazyModule.scala 167:31]
  assign acc_auto_bus_in_aw_bits_size = bus_auto_out_20_aw_bits_size; // @[LazyModule.scala 167:31]
  assign acc_auto_bus_in_w_valid = bus_auto_out_20_w_valid; // @[LazyModule.scala 167:31]
  assign acc_auto_bus_in_w_bits_data = bus_auto_out_20_w_bits_data; // @[LazyModule.scala 167:31]
  assign acc_auto_bus_in_w_bits_strb = bus_auto_out_20_w_bits_strb; // @[LazyModule.scala 167:31]
  assign acc_auto_bus_in_w_bits_last = bus_auto_out_20_w_bits_last; // @[LazyModule.scala 167:31]
  assign acc_auto_bus_in_b_ready = bus_auto_out_20_b_ready; // @[LazyModule.scala 167:31]
  assign acc_auto_bus_in_ar_valid = bus_auto_out_20_ar_valid; // @[LazyModule.scala 167:31]
  assign acc_auto_bus_in_ar_bits_id = bus_auto_out_20_ar_bits_id; // @[LazyModule.scala 167:31]
  assign acc_auto_bus_in_ar_bits_addr = bus_auto_out_20_ar_bits_addr; // @[LazyModule.scala 167:31]
  assign acc_auto_bus_in_ar_bits_size = bus_auto_out_20_ar_bits_size; // @[LazyModule.scala 167:31]
  assign acc_auto_bus_in_r_ready = bus_auto_out_20_r_ready; // @[LazyModule.scala 167:31]
  assign acc_auto_dspQueue_stream_out_ready = widthAdapter_1_auto_in_ready; // @[LazyModule.scala 167:57]
  assign acc_auto_accumulator_slave_in_valid = buffer_2_auto_out_valid; // @[LazyModule.scala 167:31]
  assign acc_auto_accumulator_slave_in_bits_data = buffer_2_auto_out_bits_data; // @[LazyModule.scala 167:31]
  assign acc_auto_accumulator_slave_in_bits_last = buffer_2_auto_out_bits_last; // @[LazyModule.scala 167:31]
  assign widthAdapter_1_clock = clock;
  assign widthAdapter_1_reset = reset;
  assign widthAdapter_1_auto_in_valid = acc_auto_dspQueue_stream_out_valid; // @[LazyModule.scala 167:57]
  assign widthAdapter_1_auto_in_bits_data = acc_auto_dspQueue_stream_out_bits_data; // @[LazyModule.scala 167:57]
  assign widthAdapter_1_auto_in_bits_last = acc_auto_dspQueue_stream_out_bits_last; // @[LazyModule.scala 167:57]
  assign widthAdapter_1_auto_out_ready = acc_queue_auto_in_in_ready; // @[LazyModule.scala 167:57]
  assign acc_queue_clock = clock;
  assign acc_queue_reset = reset;
  assign acc_queue_auto_out_out_ready = out_mux_auto_stream_in_0_ready; // @[LazyModule.scala 167:57]
  assign acc_queue_auto_in_in_valid = widthAdapter_1_auto_out_valid; // @[LazyModule.scala 167:57]
  assign acc_queue_auto_in_in_bits_data = widthAdapter_1_auto_out_bits_data; // @[LazyModule.scala 167:57]
  assign acc_queue_auto_in_in_bits_last = widthAdapter_1_auto_out_bits_last; // @[LazyModule.scala 167:57]
  assign out_mux_clock = clock;
  assign out_mux_reset = reset;
  assign out_mux_auto_register_in_aw_valid = axi4buf_17_auto_out_aw_valid; // @[LazyModule.scala 167:31]
  assign out_mux_auto_register_in_aw_bits_id = axi4buf_17_auto_out_aw_bits_id; // @[LazyModule.scala 167:31]
  assign out_mux_auto_register_in_aw_bits_addr = axi4buf_17_auto_out_aw_bits_addr; // @[LazyModule.scala 167:31]
  assign out_mux_auto_register_in_w_valid = axi4buf_17_auto_out_w_valid; // @[LazyModule.scala 167:31]
  assign out_mux_auto_register_in_w_bits_data = axi4buf_17_auto_out_w_bits_data; // @[LazyModule.scala 167:31]
  assign out_mux_auto_register_in_w_bits_strb = axi4buf_17_auto_out_w_bits_strb; // @[LazyModule.scala 167:31]
  assign out_mux_auto_register_in_b_ready = axi4buf_17_auto_out_b_ready; // @[LazyModule.scala 167:31]
  assign out_mux_auto_register_in_ar_valid = axi4buf_17_auto_out_ar_valid; // @[LazyModule.scala 167:31]
  assign out_mux_auto_register_in_ar_bits_id = axi4buf_17_auto_out_ar_bits_id; // @[LazyModule.scala 167:31]
  assign out_mux_auto_register_in_ar_bits_addr = axi4buf_17_auto_out_ar_bits_addr; // @[LazyModule.scala 167:31]
  assign out_mux_auto_register_in_ar_bits_size = axi4buf_17_auto_out_ar_bits_size; // @[LazyModule.scala 167:31]
  assign out_mux_auto_register_in_r_ready = axi4buf_17_auto_out_r_ready; // @[LazyModule.scala 167:31]
  assign out_mux_auto_stream_in_6_valid = buffer_8_auto_out_valid; // @[LazyModule.scala 167:31]
  assign out_mux_auto_stream_in_6_bits_data = buffer_8_auto_out_bits_data; // @[LazyModule.scala 167:31]
  assign out_mux_auto_stream_in_6_bits_last = buffer_8_auto_out_bits_last; // @[LazyModule.scala 167:31]
  assign out_mux_auto_stream_in_5_valid = buffer_7_auto_out_valid; // @[LazyModule.scala 167:31]
  assign out_mux_auto_stream_in_5_bits_data = buffer_7_auto_out_bits_data; // @[LazyModule.scala 167:31]
  assign out_mux_auto_stream_in_5_bits_last = buffer_7_auto_out_bits_last; // @[LazyModule.scala 167:31]
  assign out_mux_auto_stream_in_4_valid = buffer_6_auto_out_valid; // @[LazyModule.scala 167:31]
  assign out_mux_auto_stream_in_4_bits_data = buffer_6_auto_out_bits_data; // @[LazyModule.scala 167:31]
  assign out_mux_auto_stream_in_4_bits_last = buffer_6_auto_out_bits_last; // @[LazyModule.scala 167:31]
  assign out_mux_auto_stream_in_3_valid = buffer_5_auto_out_valid; // @[LazyModule.scala 167:31]
  assign out_mux_auto_stream_in_3_bits_data = buffer_5_auto_out_bits_data; // @[LazyModule.scala 167:31]
  assign out_mux_auto_stream_in_3_bits_last = buffer_5_auto_out_bits_last; // @[LazyModule.scala 167:31]
  assign out_mux_auto_stream_in_2_valid = buffer_4_auto_out_valid; // @[LazyModule.scala 167:31]
  assign out_mux_auto_stream_in_2_bits_data = buffer_4_auto_out_bits_data; // @[LazyModule.scala 167:31]
  assign out_mux_auto_stream_in_2_bits_last = buffer_4_auto_out_bits_last; // @[LazyModule.scala 167:31]
  assign out_mux_auto_stream_in_1_valid = buffer_3_auto_out_valid; // @[LazyModule.scala 167:31]
  assign out_mux_auto_stream_in_1_bits_data = buffer_3_auto_out_bits_data; // @[LazyModule.scala 167:31]
  assign out_mux_auto_stream_in_1_bits_last = buffer_3_auto_out_bits_last; // @[LazyModule.scala 167:31]
  assign out_mux_auto_stream_in_0_valid = acc_queue_auto_out_out_valid; // @[LazyModule.scala 167:57]
  assign out_mux_auto_stream_in_0_bits_data = acc_queue_auto_out_out_bits_data; // @[LazyModule.scala 167:57]
  assign out_mux_auto_stream_in_0_bits_last = acc_queue_auto_out_out_bits_last; // @[LazyModule.scala 167:57]
  assign out_mux_auto_stream_out_1_ready = uTx_queue_auto_in_in_ready; // @[LazyModule.scala 167:57]
  assign out_mux_auto_stream_out_0_ready = buffer_9_auto_in_ready; // @[LazyModule.scala 167:57]
  assign out_queue_clock = clock;
  assign out_queue_reset = reset;
  assign out_queue_auto_out_out_ready = widthAdapter_2_auto_in_ready; // @[LazyModule.scala 167:57]
  assign out_queue_auto_in_in_valid = buffer_9_auto_out_valid; // @[LazyModule.scala 167:31]
  assign out_queue_auto_in_in_bits_data = buffer_9_auto_out_bits_data; // @[LazyModule.scala 167:31]
  assign out_queue_auto_in_in_bits_last = buffer_9_auto_out_bits_last; // @[LazyModule.scala 167:31]
  assign widthAdapter_2_clock = clock;
  assign widthAdapter_2_reset = reset;
  assign widthAdapter_2_auto_in_valid = out_queue_auto_out_out_valid; // @[LazyModule.scala 167:57]
  assign widthAdapter_2_auto_in_bits_data = out_queue_auto_out_out_bits_data; // @[LazyModule.scala 167:57]
  assign widthAdapter_2_auto_in_bits_last = out_queue_auto_out_out_bits_last; // @[LazyModule.scala 167:57]
  assign widthAdapter_2_auto_out_ready = converter_1_auto_in_ready; // @[LazyModule.scala 167:57]
  assign uTx_queue_clock = clock;
  assign uTx_queue_reset = reset;
  assign uTx_queue_auto_out_out_ready = widthAdapter_3_auto_in_ready; // @[LazyModule.scala 167:57]
  assign uTx_queue_auto_in_in_valid = out_mux_auto_stream_out_1_valid; // @[LazyModule.scala 167:57]
  assign uTx_queue_auto_in_in_bits_data = out_mux_auto_stream_out_1_bits_data; // @[LazyModule.scala 167:57]
  assign uTx_queue_auto_in_in_bits_last = out_mux_auto_stream_out_1_bits_last; // @[LazyModule.scala 167:57]
  assign widthAdapter_3_clock = clock;
  assign widthAdapter_3_reset = reset;
  assign widthAdapter_3_auto_in_valid = uTx_queue_auto_out_out_valid; // @[LazyModule.scala 167:57]
  assign widthAdapter_3_auto_in_bits_data = uTx_queue_auto_out_out_bits_data; // @[LazyModule.scala 167:57]
  assign widthAdapter_3_auto_in_bits_last = uTx_queue_auto_out_out_bits_last; // @[LazyModule.scala 167:57]
  assign widthAdapter_3_auto_out_ready = uart_auto_in_in_ready; // @[LazyModule.scala 167:57]
  assign widthAdapter_4_clock = clock;
  assign widthAdapter_4_reset = reset;
  assign widthAdapter_4_auto_in_valid = uart_auto_out_out_valid; // @[LazyModule.scala 167:31]
  assign widthAdapter_4_auto_in_bits_data = uart_auto_out_out_bits_data; // @[LazyModule.scala 167:31]
  assign widthAdapter_4_auto_in_bits_last = 1'h0; // @[LazyModule.scala 167:31]
  assign widthAdapter_4_auto_out_ready = uRx_split_auto_stream_in_ready; // @[LazyModule.scala 167:57]
  assign uRx_split_clock = clock;
  assign uRx_split_reset = reset;
  assign uRx_split_auto_mem_in_aw_valid = axi4buf_19_auto_out_aw_valid; // @[LazyModule.scala 167:31]
  assign uRx_split_auto_mem_in_aw_bits_id = axi4buf_19_auto_out_aw_bits_id; // @[LazyModule.scala 167:31]
  assign uRx_split_auto_mem_in_aw_bits_addr = axi4buf_19_auto_out_aw_bits_addr; // @[LazyModule.scala 167:31]
  assign uRx_split_auto_mem_in_w_valid = axi4buf_19_auto_out_w_valid; // @[LazyModule.scala 167:31]
  assign uRx_split_auto_mem_in_w_bits_data = axi4buf_19_auto_out_w_bits_data; // @[LazyModule.scala 167:31]
  assign uRx_split_auto_mem_in_w_bits_strb = axi4buf_19_auto_out_w_bits_strb; // @[LazyModule.scala 167:31]
  assign uRx_split_auto_mem_in_b_ready = axi4buf_19_auto_out_b_ready; // @[LazyModule.scala 167:31]
  assign uRx_split_auto_mem_in_ar_valid = axi4buf_19_auto_out_ar_valid; // @[LazyModule.scala 167:31]
  assign uRx_split_auto_mem_in_ar_bits_id = axi4buf_19_auto_out_ar_bits_id; // @[LazyModule.scala 167:31]
  assign uRx_split_auto_mem_in_ar_bits_addr = axi4buf_19_auto_out_ar_bits_addr; // @[LazyModule.scala 167:31]
  assign uRx_split_auto_mem_in_ar_bits_size = axi4buf_19_auto_out_ar_bits_size; // @[LazyModule.scala 167:31]
  assign uRx_split_auto_mem_in_r_ready = axi4buf_19_auto_out_r_ready; // @[LazyModule.scala 167:31]
  assign uRx_split_auto_stream_in_valid = widthAdapter_4_auto_out_valid; // @[LazyModule.scala 167:57]
  assign uRx_split_auto_stream_in_bits_data = widthAdapter_4_auto_out_bits_data; // @[LazyModule.scala 167:57]
  assign uRx_split_auto_stream_in_bits_last = widthAdapter_4_auto_out_bits_last; // @[LazyModule.scala 167:57]
  assign uRx_split_auto_stream_out_4_ready = buffer_8_auto_in_ready; // @[LazyModule.scala 167:57]
  assign uRx_split_auto_stream_out_3_ready = mag_mux_0_auto_stream_in_2_ready; // @[LazyModule.scala 167:31]
  assign uRx_split_auto_stream_out_2_ready = fft_mux_0_auto_stream_in_2_ready; // @[LazyModule.scala 167:31]
  assign uRx_split_auto_stream_out_1_ready = nco_mux_0_auto_stream_in_2_ready; // @[LazyModule.scala 167:31]
  assign uRx_split_auto_stream_out_0_ready = plfg_mux_0_auto_stream_in_2_ready; // @[LazyModule.scala 167:31]
  assign uart_clock = clock;
  assign uart_reset = reset;
  assign uart_auto_mem_in_aw_valid = axi4buf_18_auto_out_aw_valid; // @[LazyModule.scala 167:31]
  assign uart_auto_mem_in_aw_bits_id = axi4buf_18_auto_out_aw_bits_id; // @[LazyModule.scala 167:31]
  assign uart_auto_mem_in_aw_bits_addr = axi4buf_18_auto_out_aw_bits_addr; // @[LazyModule.scala 167:31]
  assign uart_auto_mem_in_w_valid = axi4buf_18_auto_out_w_valid; // @[LazyModule.scala 167:31]
  assign uart_auto_mem_in_w_bits_data = axi4buf_18_auto_out_w_bits_data; // @[LazyModule.scala 167:31]
  assign uart_auto_mem_in_w_bits_strb = axi4buf_18_auto_out_w_bits_strb; // @[LazyModule.scala 167:31]
  assign uart_auto_mem_in_b_ready = axi4buf_18_auto_out_b_ready; // @[LazyModule.scala 167:31]
  assign uart_auto_mem_in_ar_valid = axi4buf_18_auto_out_ar_valid; // @[LazyModule.scala 167:31]
  assign uart_auto_mem_in_ar_bits_id = axi4buf_18_auto_out_ar_bits_id; // @[LazyModule.scala 167:31]
  assign uart_auto_mem_in_ar_bits_addr = axi4buf_18_auto_out_ar_bits_addr; // @[LazyModule.scala 167:31]
  assign uart_auto_mem_in_ar_bits_size = axi4buf_18_auto_out_ar_bits_size; // @[LazyModule.scala 167:31]
  assign uart_auto_mem_in_r_ready = axi4buf_18_auto_out_r_ready; // @[LazyModule.scala 167:31]
  assign uart_auto_in_in_valid = widthAdapter_3_auto_out_valid; // @[LazyModule.scala 167:57]
  assign uart_auto_in_in_bits_data = widthAdapter_3_auto_out_bits_data; // @[LazyModule.scala 167:57]
  assign uart_auto_out_out_ready = widthAdapter_4_auto_in_ready; // @[LazyModule.scala 167:31]
  assign uart_io_rxd = uRx; // @[SpectrometerTest.scala 266:24]
  assign bus_clock = clock;
  assign bus_reset = reset;
  assign bus_auto_in_aw_valid = converter_auto_out_aw_valid; // @[LazyModule.scala 167:31]
  assign bus_auto_in_aw_bits_id = converter_auto_out_aw_bits_id; // @[LazyModule.scala 167:31]
  assign bus_auto_in_aw_bits_addr = converter_auto_out_aw_bits_addr; // @[LazyModule.scala 167:31]
  assign bus_auto_in_aw_bits_size = converter_auto_out_aw_bits_size; // @[LazyModule.scala 167:31]
  assign bus_auto_in_w_valid = converter_auto_out_w_valid; // @[LazyModule.scala 167:31]
  assign bus_auto_in_w_bits_data = converter_auto_out_w_bits_data; // @[LazyModule.scala 167:31]
  assign bus_auto_in_w_bits_strb = converter_auto_out_w_bits_strb; // @[LazyModule.scala 167:31]
  assign bus_auto_in_w_bits_last = converter_auto_out_w_bits_last; // @[LazyModule.scala 167:31]
  assign bus_auto_in_b_ready = converter_auto_out_b_ready; // @[LazyModule.scala 167:31]
  assign bus_auto_in_ar_valid = converter_auto_out_ar_valid; // @[LazyModule.scala 167:31]
  assign bus_auto_in_ar_bits_id = converter_auto_out_ar_bits_id; // @[LazyModule.scala 167:31]
  assign bus_auto_in_ar_bits_addr = converter_auto_out_ar_bits_addr; // @[LazyModule.scala 167:31]
  assign bus_auto_in_ar_bits_size = converter_auto_out_ar_bits_size; // @[LazyModule.scala 167:31]
  assign bus_auto_in_r_ready = converter_auto_out_r_ready; // @[LazyModule.scala 167:31]
  assign bus_auto_out_20_aw_ready = acc_auto_bus_in_aw_ready; // @[LazyModule.scala 167:31]
  assign bus_auto_out_20_w_ready = acc_auto_bus_in_w_ready; // @[LazyModule.scala 167:31]
  assign bus_auto_out_20_b_valid = acc_auto_bus_in_b_valid; // @[LazyModule.scala 167:31]
  assign bus_auto_out_20_b_bits_resp = acc_auto_bus_in_b_bits_resp; // @[LazyModule.scala 167:31]
  assign bus_auto_out_20_ar_ready = acc_auto_bus_in_ar_ready; // @[LazyModule.scala 167:31]
  assign bus_auto_out_20_r_valid = acc_auto_bus_in_r_valid; // @[LazyModule.scala 167:31]
  assign bus_auto_out_20_r_bits_data = acc_auto_bus_in_r_bits_data; // @[LazyModule.scala 167:31]
  assign bus_auto_out_20_r_bits_resp = acc_auto_bus_in_r_bits_resp; // @[LazyModule.scala 167:31]
  assign bus_auto_out_20_r_bits_last = acc_auto_bus_in_r_bits_last; // @[LazyModule.scala 167:31]
  assign bus_auto_out_19_aw_ready = axi4buf_19_auto_in_aw_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_19_w_ready = axi4buf_19_auto_in_w_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_19_b_valid = axi4buf_19_auto_in_b_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_19_b_bits_id = axi4buf_19_auto_in_b_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_19_b_bits_resp = axi4buf_19_auto_in_b_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_19_ar_ready = axi4buf_19_auto_in_ar_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_19_r_valid = axi4buf_19_auto_in_r_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_19_r_bits_id = axi4buf_19_auto_in_r_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_19_r_bits_data = axi4buf_19_auto_in_r_bits_data; // @[LazyModule.scala 167:57]
  assign bus_auto_out_19_r_bits_resp = axi4buf_19_auto_in_r_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_19_r_bits_last = axi4buf_19_auto_in_r_bits_last; // @[LazyModule.scala 167:57]
  assign bus_auto_out_18_aw_ready = axi4buf_18_auto_in_aw_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_18_w_ready = axi4buf_18_auto_in_w_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_18_b_valid = axi4buf_18_auto_in_b_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_18_b_bits_id = axi4buf_18_auto_in_b_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_18_b_bits_resp = axi4buf_18_auto_in_b_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_18_ar_ready = axi4buf_18_auto_in_ar_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_18_r_valid = axi4buf_18_auto_in_r_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_18_r_bits_id = axi4buf_18_auto_in_r_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_18_r_bits_data = axi4buf_18_auto_in_r_bits_data; // @[LazyModule.scala 167:57]
  assign bus_auto_out_18_r_bits_resp = axi4buf_18_auto_in_r_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_18_r_bits_last = axi4buf_18_auto_in_r_bits_last; // @[LazyModule.scala 167:57]
  assign bus_auto_out_17_aw_ready = axi4buf_17_auto_in_aw_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_17_w_ready = axi4buf_17_auto_in_w_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_17_b_valid = axi4buf_17_auto_in_b_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_17_b_bits_id = axi4buf_17_auto_in_b_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_17_b_bits_resp = axi4buf_17_auto_in_b_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_17_ar_ready = axi4buf_17_auto_in_ar_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_17_r_valid = axi4buf_17_auto_in_r_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_17_r_bits_id = axi4buf_17_auto_in_r_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_17_r_bits_data = axi4buf_17_auto_in_r_bits_data; // @[LazyModule.scala 167:57]
  assign bus_auto_out_17_r_bits_resp = axi4buf_17_auto_in_r_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_17_r_bits_last = axi4buf_17_auto_in_r_bits_last; // @[LazyModule.scala 167:57]
  assign bus_auto_out_16_aw_ready = axi4buf_16_auto_in_aw_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_16_w_ready = axi4buf_16_auto_in_w_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_16_b_valid = axi4buf_16_auto_in_b_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_16_b_bits_id = axi4buf_16_auto_in_b_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_16_b_bits_resp = axi4buf_16_auto_in_b_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_16_ar_ready = axi4buf_16_auto_in_ar_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_16_r_valid = axi4buf_16_auto_in_r_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_16_r_bits_id = axi4buf_16_auto_in_r_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_16_r_bits_data = axi4buf_16_auto_in_r_bits_data; // @[LazyModule.scala 167:57]
  assign bus_auto_out_16_r_bits_resp = axi4buf_16_auto_in_r_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_16_r_bits_last = axi4buf_16_auto_in_r_bits_last; // @[LazyModule.scala 167:57]
  assign bus_auto_out_15_aw_ready = axi4buf_15_auto_in_aw_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_15_w_ready = axi4buf_15_auto_in_w_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_15_b_valid = axi4buf_15_auto_in_b_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_15_b_bits_id = axi4buf_15_auto_in_b_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_15_b_bits_resp = axi4buf_15_auto_in_b_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_15_ar_ready = axi4buf_15_auto_in_ar_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_15_r_valid = axi4buf_15_auto_in_r_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_15_r_bits_id = axi4buf_15_auto_in_r_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_15_r_bits_data = axi4buf_15_auto_in_r_bits_data; // @[LazyModule.scala 167:57]
  assign bus_auto_out_15_r_bits_resp = axi4buf_15_auto_in_r_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_15_r_bits_last = axi4buf_15_auto_in_r_bits_last; // @[LazyModule.scala 167:57]
  assign bus_auto_out_14_aw_ready = axi4buf_14_auto_in_aw_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_14_w_ready = axi4buf_14_auto_in_w_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_14_b_valid = axi4buf_14_auto_in_b_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_14_b_bits_id = axi4buf_14_auto_in_b_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_14_b_bits_resp = axi4buf_14_auto_in_b_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_14_ar_ready = axi4buf_14_auto_in_ar_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_14_r_valid = axi4buf_14_auto_in_r_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_14_r_bits_id = axi4buf_14_auto_in_r_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_14_r_bits_data = axi4buf_14_auto_in_r_bits_data; // @[LazyModule.scala 167:57]
  assign bus_auto_out_14_r_bits_resp = axi4buf_14_auto_in_r_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_14_r_bits_last = axi4buf_14_auto_in_r_bits_last; // @[LazyModule.scala 167:57]
  assign bus_auto_out_13_aw_ready = axi4buf_13_auto_in_aw_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_13_w_ready = axi4buf_13_auto_in_w_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_13_b_valid = axi4buf_13_auto_in_b_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_13_b_bits_id = axi4buf_13_auto_in_b_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_13_b_bits_resp = axi4buf_13_auto_in_b_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_13_ar_ready = axi4buf_13_auto_in_ar_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_13_r_valid = axi4buf_13_auto_in_r_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_13_r_bits_id = axi4buf_13_auto_in_r_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_13_r_bits_data = axi4buf_13_auto_in_r_bits_data; // @[LazyModule.scala 167:57]
  assign bus_auto_out_13_r_bits_resp = axi4buf_13_auto_in_r_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_13_r_bits_last = axi4buf_13_auto_in_r_bits_last; // @[LazyModule.scala 167:57]
  assign bus_auto_out_12_aw_ready = axi4buf_12_auto_in_aw_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_12_w_ready = axi4buf_12_auto_in_w_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_12_b_valid = axi4buf_12_auto_in_b_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_12_b_bits_id = axi4buf_12_auto_in_b_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_12_b_bits_resp = axi4buf_12_auto_in_b_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_12_ar_ready = axi4buf_12_auto_in_ar_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_12_r_valid = axi4buf_12_auto_in_r_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_12_r_bits_id = axi4buf_12_auto_in_r_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_12_r_bits_data = axi4buf_12_auto_in_r_bits_data; // @[LazyModule.scala 167:57]
  assign bus_auto_out_12_r_bits_resp = axi4buf_12_auto_in_r_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_12_r_bits_last = axi4buf_12_auto_in_r_bits_last; // @[LazyModule.scala 167:57]
  assign bus_auto_out_11_aw_ready = axi4buf_11_auto_in_aw_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_11_w_ready = axi4buf_11_auto_in_w_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_11_b_valid = axi4buf_11_auto_in_b_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_11_b_bits_id = axi4buf_11_auto_in_b_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_11_b_bits_resp = axi4buf_11_auto_in_b_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_11_ar_ready = axi4buf_11_auto_in_ar_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_11_r_valid = axi4buf_11_auto_in_r_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_11_r_bits_id = axi4buf_11_auto_in_r_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_11_r_bits_data = axi4buf_11_auto_in_r_bits_data; // @[LazyModule.scala 167:57]
  assign bus_auto_out_11_r_bits_resp = axi4buf_11_auto_in_r_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_11_r_bits_last = axi4buf_11_auto_in_r_bits_last; // @[LazyModule.scala 167:57]
  assign bus_auto_out_10_aw_ready = axi4buf_10_auto_in_aw_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_10_w_ready = axi4buf_10_auto_in_w_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_10_b_valid = axi4buf_10_auto_in_b_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_10_b_bits_id = axi4buf_10_auto_in_b_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_10_b_bits_resp = axi4buf_10_auto_in_b_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_10_ar_ready = axi4buf_10_auto_in_ar_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_10_r_valid = axi4buf_10_auto_in_r_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_10_r_bits_id = axi4buf_10_auto_in_r_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_10_r_bits_data = axi4buf_10_auto_in_r_bits_data; // @[LazyModule.scala 167:57]
  assign bus_auto_out_10_r_bits_resp = axi4buf_10_auto_in_r_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_10_r_bits_last = axi4buf_10_auto_in_r_bits_last; // @[LazyModule.scala 167:57]
  assign bus_auto_out_9_aw_ready = axi4buf_9_auto_in_aw_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_9_w_ready = axi4buf_9_auto_in_w_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_9_b_valid = axi4buf_9_auto_in_b_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_9_b_bits_id = axi4buf_9_auto_in_b_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_9_b_bits_resp = axi4buf_9_auto_in_b_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_9_ar_ready = axi4buf_9_auto_in_ar_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_9_r_valid = axi4buf_9_auto_in_r_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_9_r_bits_id = axi4buf_9_auto_in_r_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_9_r_bits_data = axi4buf_9_auto_in_r_bits_data; // @[LazyModule.scala 167:57]
  assign bus_auto_out_9_r_bits_resp = axi4buf_9_auto_in_r_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_9_r_bits_last = axi4buf_9_auto_in_r_bits_last; // @[LazyModule.scala 167:57]
  assign bus_auto_out_8_aw_ready = axi4buf_8_auto_in_aw_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_8_w_ready = axi4buf_8_auto_in_w_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_8_b_valid = axi4buf_8_auto_in_b_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_8_b_bits_id = axi4buf_8_auto_in_b_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_8_b_bits_resp = axi4buf_8_auto_in_b_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_8_ar_ready = axi4buf_8_auto_in_ar_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_8_r_valid = axi4buf_8_auto_in_r_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_8_r_bits_id = axi4buf_8_auto_in_r_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_8_r_bits_data = axi4buf_8_auto_in_r_bits_data; // @[LazyModule.scala 167:57]
  assign bus_auto_out_8_r_bits_resp = axi4buf_8_auto_in_r_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_8_r_bits_last = axi4buf_8_auto_in_r_bits_last; // @[LazyModule.scala 167:57]
  assign bus_auto_out_7_aw_ready = axi4buf_7_auto_in_aw_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_7_w_ready = axi4buf_7_auto_in_w_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_7_b_valid = axi4buf_7_auto_in_b_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_7_b_bits_id = axi4buf_7_auto_in_b_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_7_b_bits_resp = axi4buf_7_auto_in_b_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_7_ar_ready = axi4buf_7_auto_in_ar_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_7_r_valid = axi4buf_7_auto_in_r_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_7_r_bits_id = axi4buf_7_auto_in_r_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_7_r_bits_data = axi4buf_7_auto_in_r_bits_data; // @[LazyModule.scala 167:57]
  assign bus_auto_out_7_r_bits_resp = axi4buf_7_auto_in_r_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_7_r_bits_last = axi4buf_7_auto_in_r_bits_last; // @[LazyModule.scala 167:57]
  assign bus_auto_out_6_aw_ready = axi4buf_6_auto_in_aw_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_6_w_ready = axi4buf_6_auto_in_w_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_6_b_valid = axi4buf_6_auto_in_b_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_6_b_bits_id = axi4buf_6_auto_in_b_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_6_b_bits_resp = axi4buf_6_auto_in_b_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_6_ar_ready = axi4buf_6_auto_in_ar_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_6_r_valid = axi4buf_6_auto_in_r_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_6_r_bits_id = axi4buf_6_auto_in_r_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_6_r_bits_data = axi4buf_6_auto_in_r_bits_data; // @[LazyModule.scala 167:57]
  assign bus_auto_out_6_r_bits_resp = axi4buf_6_auto_in_r_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_6_r_bits_last = axi4buf_6_auto_in_r_bits_last; // @[LazyModule.scala 167:57]
  assign bus_auto_out_5_aw_ready = axi4buf_5_auto_in_aw_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_5_w_ready = axi4buf_5_auto_in_w_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_5_b_valid = axi4buf_5_auto_in_b_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_5_b_bits_id = axi4buf_5_auto_in_b_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_5_b_bits_resp = axi4buf_5_auto_in_b_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_5_ar_ready = axi4buf_5_auto_in_ar_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_5_r_valid = axi4buf_5_auto_in_r_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_5_r_bits_id = axi4buf_5_auto_in_r_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_5_r_bits_data = axi4buf_5_auto_in_r_bits_data; // @[LazyModule.scala 167:57]
  assign bus_auto_out_5_r_bits_resp = axi4buf_5_auto_in_r_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_5_r_bits_last = axi4buf_5_auto_in_r_bits_last; // @[LazyModule.scala 167:57]
  assign bus_auto_out_4_aw_ready = axi4buf_4_auto_in_aw_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_4_w_ready = axi4buf_4_auto_in_w_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_4_b_valid = axi4buf_4_auto_in_b_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_4_b_bits_id = axi4buf_4_auto_in_b_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_4_b_bits_resp = axi4buf_4_auto_in_b_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_4_ar_ready = axi4buf_4_auto_in_ar_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_4_r_valid = axi4buf_4_auto_in_r_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_4_r_bits_id = axi4buf_4_auto_in_r_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_4_r_bits_data = axi4buf_4_auto_in_r_bits_data; // @[LazyModule.scala 167:57]
  assign bus_auto_out_4_r_bits_resp = axi4buf_4_auto_in_r_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_4_r_bits_last = axi4buf_4_auto_in_r_bits_last; // @[LazyModule.scala 167:57]
  assign bus_auto_out_3_aw_ready = axi4buf_3_auto_in_aw_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_3_w_ready = axi4buf_3_auto_in_w_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_3_b_valid = axi4buf_3_auto_in_b_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_3_b_bits_id = axi4buf_3_auto_in_b_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_3_b_bits_resp = axi4buf_3_auto_in_b_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_3_ar_ready = axi4buf_3_auto_in_ar_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_3_r_valid = axi4buf_3_auto_in_r_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_3_r_bits_id = axi4buf_3_auto_in_r_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_3_r_bits_data = axi4buf_3_auto_in_r_bits_data; // @[LazyModule.scala 167:57]
  assign bus_auto_out_3_r_bits_resp = axi4buf_3_auto_in_r_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_3_r_bits_last = axi4buf_3_auto_in_r_bits_last; // @[LazyModule.scala 167:57]
  assign bus_auto_out_2_aw_ready = axi4buf_2_auto_in_aw_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_2_w_ready = axi4buf_2_auto_in_w_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_2_b_valid = axi4buf_2_auto_in_b_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_2_b_bits_id = axi4buf_2_auto_in_b_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_2_b_bits_resp = axi4buf_2_auto_in_b_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_2_ar_ready = axi4buf_2_auto_in_ar_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_2_r_valid = axi4buf_2_auto_in_r_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_2_r_bits_id = axi4buf_2_auto_in_r_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_2_r_bits_data = axi4buf_2_auto_in_r_bits_data; // @[LazyModule.scala 167:57]
  assign bus_auto_out_2_r_bits_resp = axi4buf_2_auto_in_r_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_2_r_bits_last = axi4buf_2_auto_in_r_bits_last; // @[LazyModule.scala 167:57]
  assign bus_auto_out_1_aw_ready = axi4buf_1_auto_in_aw_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_1_w_ready = axi4buf_1_auto_in_w_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_1_b_valid = axi4buf_1_auto_in_b_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_1_b_bits_id = axi4buf_1_auto_in_b_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_1_b_bits_resp = axi4buf_1_auto_in_b_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_1_ar_ready = axi4buf_1_auto_in_ar_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_1_r_valid = axi4buf_1_auto_in_r_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_1_r_bits_id = axi4buf_1_auto_in_r_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_1_r_bits_data = axi4buf_1_auto_in_r_bits_data; // @[LazyModule.scala 167:57]
  assign bus_auto_out_1_r_bits_resp = axi4buf_1_auto_in_r_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_1_r_bits_last = axi4buf_1_auto_in_r_bits_last; // @[LazyModule.scala 167:57]
  assign bus_auto_out_0_aw_ready = axi4buf_auto_in_aw_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_0_w_ready = axi4buf_auto_in_w_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_0_b_valid = axi4buf_auto_in_b_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_0_b_bits_id = axi4buf_auto_in_b_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_0_b_bits_resp = axi4buf_auto_in_b_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_0_ar_ready = axi4buf_auto_in_ar_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_0_r_valid = axi4buf_auto_in_r_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_0_r_bits_id = axi4buf_auto_in_r_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_0_r_bits_data = axi4buf_auto_in_r_bits_data; // @[LazyModule.scala 167:57]
  assign bus_auto_out_0_r_bits_resp = axi4buf_auto_in_r_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_0_r_bits_last = axi4buf_auto_in_r_bits_last; // @[LazyModule.scala 167:57]
  assign axi4buf_clock = clock;
  assign axi4buf_reset = reset;
  assign axi4buf_auto_in_aw_valid = bus_auto_out_0_aw_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_auto_in_aw_bits_id = bus_auto_out_0_aw_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_auto_in_aw_bits_addr = bus_auto_out_0_aw_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_auto_in_aw_bits_size = bus_auto_out_0_aw_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_auto_in_w_valid = bus_auto_out_0_w_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_auto_in_w_bits_data = bus_auto_out_0_w_bits_data; // @[LazyModule.scala 167:57]
  assign axi4buf_auto_in_w_bits_strb = bus_auto_out_0_w_bits_strb; // @[LazyModule.scala 167:57]
  assign axi4buf_auto_in_w_bits_last = bus_auto_out_0_w_bits_last; // @[LazyModule.scala 167:57]
  assign axi4buf_auto_in_b_ready = bus_auto_out_0_b_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_auto_in_ar_valid = bus_auto_out_0_ar_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_auto_in_ar_bits_id = bus_auto_out_0_ar_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_auto_in_ar_bits_addr = bus_auto_out_0_ar_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_auto_in_ar_bits_size = bus_auto_out_0_ar_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_auto_in_r_ready = bus_auto_out_0_r_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_auto_out_aw_ready = in_split_auto_mem_in_aw_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_auto_out_w_ready = in_split_auto_mem_in_w_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_auto_out_b_valid = in_split_auto_mem_in_b_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_auto_out_b_bits_id = in_split_auto_mem_in_b_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_auto_out_b_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_auto_out_ar_ready = in_split_auto_mem_in_ar_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_auto_out_r_valid = in_split_auto_mem_in_r_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_auto_out_r_bits_id = in_split_auto_mem_in_r_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_auto_out_r_bits_data = in_split_auto_mem_in_r_bits_data; // @[LazyModule.scala 167:31]
  assign axi4buf_auto_out_r_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_auto_out_r_bits_last = 1'h1; // @[LazyModule.scala 167:31]
  assign axi4buf_1_clock = clock;
  assign axi4buf_1_reset = reset;
  assign axi4buf_1_auto_in_aw_valid = bus_auto_out_1_aw_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_1_auto_in_aw_bits_id = bus_auto_out_1_aw_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_1_auto_in_aw_bits_addr = bus_auto_out_1_aw_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_1_auto_in_aw_bits_size = bus_auto_out_1_aw_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_1_auto_in_w_valid = bus_auto_out_1_w_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_1_auto_in_w_bits_data = bus_auto_out_1_w_bits_data; // @[LazyModule.scala 167:57]
  assign axi4buf_1_auto_in_w_bits_strb = bus_auto_out_1_w_bits_strb; // @[LazyModule.scala 167:57]
  assign axi4buf_1_auto_in_w_bits_last = bus_auto_out_1_w_bits_last; // @[LazyModule.scala 167:57]
  assign axi4buf_1_auto_in_b_ready = bus_auto_out_1_b_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_1_auto_in_ar_valid = bus_auto_out_1_ar_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_1_auto_in_ar_bits_id = bus_auto_out_1_ar_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_1_auto_in_ar_bits_addr = bus_auto_out_1_ar_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_1_auto_in_ar_bits_size = bus_auto_out_1_ar_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_1_auto_in_r_ready = bus_auto_out_1_r_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_1_auto_out_aw_ready = plfg_auto_mem_in_aw_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_1_auto_out_w_ready = plfg_auto_mem_in_w_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_1_auto_out_b_valid = plfg_auto_mem_in_b_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_1_auto_out_b_bits_id = 1'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_1_auto_out_b_bits_resp = plfg_auto_mem_in_b_bits_resp; // @[LazyModule.scala 167:31]
  assign axi4buf_1_auto_out_ar_ready = plfg_auto_mem_in_ar_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_1_auto_out_r_valid = plfg_auto_mem_in_r_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_1_auto_out_r_bits_id = 1'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_1_auto_out_r_bits_data = plfg_auto_mem_in_r_bits_data; // @[LazyModule.scala 167:31]
  assign axi4buf_1_auto_out_r_bits_resp = plfg_auto_mem_in_r_bits_resp; // @[LazyModule.scala 167:31]
  assign axi4buf_1_auto_out_r_bits_last = plfg_auto_mem_in_r_bits_last; // @[LazyModule.scala 167:31]
  assign axi4buf_2_clock = clock;
  assign axi4buf_2_reset = reset;
  assign axi4buf_2_auto_in_aw_valid = bus_auto_out_2_aw_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_2_auto_in_aw_bits_id = bus_auto_out_2_aw_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_2_auto_in_aw_bits_addr = bus_auto_out_2_aw_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_2_auto_in_aw_bits_size = bus_auto_out_2_aw_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_2_auto_in_w_valid = bus_auto_out_2_w_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_2_auto_in_w_bits_data = bus_auto_out_2_w_bits_data; // @[LazyModule.scala 167:57]
  assign axi4buf_2_auto_in_w_bits_strb = bus_auto_out_2_w_bits_strb; // @[LazyModule.scala 167:57]
  assign axi4buf_2_auto_in_w_bits_last = bus_auto_out_2_w_bits_last; // @[LazyModule.scala 167:57]
  assign axi4buf_2_auto_in_b_ready = bus_auto_out_2_b_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_2_auto_in_ar_valid = bus_auto_out_2_ar_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_2_auto_in_ar_bits_id = bus_auto_out_2_ar_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_2_auto_in_ar_bits_addr = bus_auto_out_2_ar_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_2_auto_in_ar_bits_size = bus_auto_out_2_ar_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_2_auto_in_r_ready = bus_auto_out_2_r_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_2_auto_out_aw_ready = plfg_split_auto_mem_in_aw_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_2_auto_out_w_ready = plfg_split_auto_mem_in_w_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_2_auto_out_b_valid = plfg_split_auto_mem_in_b_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_2_auto_out_b_bits_id = plfg_split_auto_mem_in_b_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_2_auto_out_b_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_2_auto_out_ar_ready = plfg_split_auto_mem_in_ar_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_2_auto_out_r_valid = plfg_split_auto_mem_in_r_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_2_auto_out_r_bits_id = plfg_split_auto_mem_in_r_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_2_auto_out_r_bits_data = plfg_split_auto_mem_in_r_bits_data; // @[LazyModule.scala 167:31]
  assign axi4buf_2_auto_out_r_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_2_auto_out_r_bits_last = 1'h1; // @[LazyModule.scala 167:31]
  assign axi4buf_3_clock = clock;
  assign axi4buf_3_reset = reset;
  assign axi4buf_3_auto_in_aw_valid = bus_auto_out_3_aw_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_3_auto_in_aw_bits_id = bus_auto_out_3_aw_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_3_auto_in_aw_bits_addr = bus_auto_out_3_aw_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_3_auto_in_aw_bits_size = bus_auto_out_3_aw_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_3_auto_in_w_valid = bus_auto_out_3_w_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_3_auto_in_w_bits_data = bus_auto_out_3_w_bits_data; // @[LazyModule.scala 167:57]
  assign axi4buf_3_auto_in_w_bits_strb = bus_auto_out_3_w_bits_strb; // @[LazyModule.scala 167:57]
  assign axi4buf_3_auto_in_w_bits_last = bus_auto_out_3_w_bits_last; // @[LazyModule.scala 167:57]
  assign axi4buf_3_auto_in_b_ready = bus_auto_out_3_b_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_3_auto_in_ar_valid = bus_auto_out_3_ar_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_3_auto_in_ar_bits_id = bus_auto_out_3_ar_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_3_auto_in_ar_bits_addr = bus_auto_out_3_ar_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_3_auto_in_ar_bits_size = bus_auto_out_3_ar_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_3_auto_in_r_ready = bus_auto_out_3_r_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_3_auto_out_aw_ready = plfg_mux_0_auto_register_in_aw_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_3_auto_out_w_ready = plfg_mux_0_auto_register_in_w_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_3_auto_out_b_valid = plfg_mux_0_auto_register_in_b_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_3_auto_out_b_bits_id = plfg_mux_0_auto_register_in_b_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_3_auto_out_b_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_3_auto_out_ar_ready = plfg_mux_0_auto_register_in_ar_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_3_auto_out_r_valid = plfg_mux_0_auto_register_in_r_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_3_auto_out_r_bits_id = plfg_mux_0_auto_register_in_r_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_3_auto_out_r_bits_data = plfg_mux_0_auto_register_in_r_bits_data; // @[LazyModule.scala 167:31]
  assign axi4buf_3_auto_out_r_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_3_auto_out_r_bits_last = 1'h1; // @[LazyModule.scala 167:31]
  assign axi4buf_4_clock = clock;
  assign axi4buf_4_reset = reset;
  assign axi4buf_4_auto_in_aw_valid = bus_auto_out_4_aw_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_4_auto_in_aw_bits_id = bus_auto_out_4_aw_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_4_auto_in_aw_bits_addr = bus_auto_out_4_aw_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_4_auto_in_aw_bits_size = bus_auto_out_4_aw_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_4_auto_in_w_valid = bus_auto_out_4_w_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_4_auto_in_w_bits_data = bus_auto_out_4_w_bits_data; // @[LazyModule.scala 167:57]
  assign axi4buf_4_auto_in_w_bits_strb = bus_auto_out_4_w_bits_strb; // @[LazyModule.scala 167:57]
  assign axi4buf_4_auto_in_w_bits_last = bus_auto_out_4_w_bits_last; // @[LazyModule.scala 167:57]
  assign axi4buf_4_auto_in_b_ready = bus_auto_out_4_b_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_4_auto_in_ar_valid = bus_auto_out_4_ar_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_4_auto_in_ar_bits_id = bus_auto_out_4_ar_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_4_auto_in_ar_bits_addr = bus_auto_out_4_ar_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_4_auto_in_ar_bits_size = bus_auto_out_4_ar_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_4_auto_in_r_ready = bus_auto_out_4_r_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_4_auto_out_aw_ready = plfg_mux_1_auto_register_in_aw_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_4_auto_out_w_ready = plfg_mux_1_auto_register_in_w_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_4_auto_out_b_valid = plfg_mux_1_auto_register_in_b_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_4_auto_out_b_bits_id = plfg_mux_1_auto_register_in_b_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_4_auto_out_b_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_4_auto_out_ar_ready = plfg_mux_1_auto_register_in_ar_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_4_auto_out_r_valid = plfg_mux_1_auto_register_in_r_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_4_auto_out_r_bits_id = plfg_mux_1_auto_register_in_r_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_4_auto_out_r_bits_data = plfg_mux_1_auto_register_in_r_bits_data; // @[LazyModule.scala 167:31]
  assign axi4buf_4_auto_out_r_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_4_auto_out_r_bits_last = 1'h1; // @[LazyModule.scala 167:31]
  assign axi4buf_5_clock = clock;
  assign axi4buf_5_reset = reset;
  assign axi4buf_5_auto_in_aw_valid = bus_auto_out_5_aw_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_5_auto_in_aw_bits_id = bus_auto_out_5_aw_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_5_auto_in_aw_bits_addr = bus_auto_out_5_aw_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_5_auto_in_aw_bits_size = bus_auto_out_5_aw_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_5_auto_in_w_valid = bus_auto_out_5_w_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_5_auto_in_w_bits_data = bus_auto_out_5_w_bits_data; // @[LazyModule.scala 167:57]
  assign axi4buf_5_auto_in_w_bits_strb = bus_auto_out_5_w_bits_strb; // @[LazyModule.scala 167:57]
  assign axi4buf_5_auto_in_w_bits_last = bus_auto_out_5_w_bits_last; // @[LazyModule.scala 167:57]
  assign axi4buf_5_auto_in_b_ready = bus_auto_out_5_b_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_5_auto_in_ar_valid = bus_auto_out_5_ar_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_5_auto_in_ar_bits_id = bus_auto_out_5_ar_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_5_auto_in_ar_bits_addr = bus_auto_out_5_ar_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_5_auto_in_ar_bits_size = bus_auto_out_5_ar_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_5_auto_in_r_ready = bus_auto_out_5_r_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_5_auto_out_aw_ready = 1'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_5_auto_out_w_ready = 1'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_5_auto_out_b_valid = 1'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_5_auto_out_b_bits_id = 1'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_5_auto_out_b_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_5_auto_out_ar_ready = 1'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_5_auto_out_r_valid = 1'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_5_auto_out_r_bits_id = 1'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_5_auto_out_r_bits_data = 32'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_5_auto_out_r_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_5_auto_out_r_bits_last = 1'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_6_clock = clock;
  assign axi4buf_6_reset = reset;
  assign axi4buf_6_auto_in_aw_valid = bus_auto_out_6_aw_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_6_auto_in_aw_bits_id = bus_auto_out_6_aw_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_6_auto_in_aw_bits_addr = bus_auto_out_6_aw_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_6_auto_in_aw_bits_size = bus_auto_out_6_aw_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_6_auto_in_w_valid = bus_auto_out_6_w_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_6_auto_in_w_bits_data = bus_auto_out_6_w_bits_data; // @[LazyModule.scala 167:57]
  assign axi4buf_6_auto_in_w_bits_strb = bus_auto_out_6_w_bits_strb; // @[LazyModule.scala 167:57]
  assign axi4buf_6_auto_in_w_bits_last = bus_auto_out_6_w_bits_last; // @[LazyModule.scala 167:57]
  assign axi4buf_6_auto_in_b_ready = bus_auto_out_6_b_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_6_auto_in_ar_valid = bus_auto_out_6_ar_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_6_auto_in_ar_bits_id = bus_auto_out_6_ar_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_6_auto_in_ar_bits_addr = bus_auto_out_6_ar_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_6_auto_in_ar_bits_size = bus_auto_out_6_ar_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_6_auto_in_r_ready = bus_auto_out_6_r_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_6_auto_out_aw_ready = nco_split_auto_mem_in_aw_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_6_auto_out_w_ready = nco_split_auto_mem_in_w_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_6_auto_out_b_valid = nco_split_auto_mem_in_b_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_6_auto_out_b_bits_id = nco_split_auto_mem_in_b_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_6_auto_out_b_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_6_auto_out_ar_ready = nco_split_auto_mem_in_ar_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_6_auto_out_r_valid = nco_split_auto_mem_in_r_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_6_auto_out_r_bits_id = nco_split_auto_mem_in_r_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_6_auto_out_r_bits_data = nco_split_auto_mem_in_r_bits_data; // @[LazyModule.scala 167:31]
  assign axi4buf_6_auto_out_r_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_6_auto_out_r_bits_last = 1'h1; // @[LazyModule.scala 167:31]
  assign axi4buf_7_clock = clock;
  assign axi4buf_7_reset = reset;
  assign axi4buf_7_auto_in_aw_valid = bus_auto_out_7_aw_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_7_auto_in_aw_bits_id = bus_auto_out_7_aw_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_7_auto_in_aw_bits_addr = bus_auto_out_7_aw_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_7_auto_in_aw_bits_size = bus_auto_out_7_aw_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_7_auto_in_w_valid = bus_auto_out_7_w_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_7_auto_in_w_bits_data = bus_auto_out_7_w_bits_data; // @[LazyModule.scala 167:57]
  assign axi4buf_7_auto_in_w_bits_strb = bus_auto_out_7_w_bits_strb; // @[LazyModule.scala 167:57]
  assign axi4buf_7_auto_in_w_bits_last = bus_auto_out_7_w_bits_last; // @[LazyModule.scala 167:57]
  assign axi4buf_7_auto_in_b_ready = bus_auto_out_7_b_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_7_auto_in_ar_valid = bus_auto_out_7_ar_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_7_auto_in_ar_bits_id = bus_auto_out_7_ar_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_7_auto_in_ar_bits_addr = bus_auto_out_7_ar_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_7_auto_in_ar_bits_size = bus_auto_out_7_ar_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_7_auto_in_r_ready = bus_auto_out_7_r_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_7_auto_out_aw_ready = nco_mux_0_auto_register_in_aw_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_7_auto_out_w_ready = nco_mux_0_auto_register_in_w_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_7_auto_out_b_valid = nco_mux_0_auto_register_in_b_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_7_auto_out_b_bits_id = nco_mux_0_auto_register_in_b_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_7_auto_out_b_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_7_auto_out_ar_ready = nco_mux_0_auto_register_in_ar_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_7_auto_out_r_valid = nco_mux_0_auto_register_in_r_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_7_auto_out_r_bits_id = nco_mux_0_auto_register_in_r_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_7_auto_out_r_bits_data = nco_mux_0_auto_register_in_r_bits_data; // @[LazyModule.scala 167:31]
  assign axi4buf_7_auto_out_r_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_7_auto_out_r_bits_last = 1'h1; // @[LazyModule.scala 167:31]
  assign axi4buf_8_clock = clock;
  assign axi4buf_8_reset = reset;
  assign axi4buf_8_auto_in_aw_valid = bus_auto_out_8_aw_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_8_auto_in_aw_bits_id = bus_auto_out_8_aw_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_8_auto_in_aw_bits_addr = bus_auto_out_8_aw_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_8_auto_in_aw_bits_size = bus_auto_out_8_aw_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_8_auto_in_w_valid = bus_auto_out_8_w_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_8_auto_in_w_bits_data = bus_auto_out_8_w_bits_data; // @[LazyModule.scala 167:57]
  assign axi4buf_8_auto_in_w_bits_strb = bus_auto_out_8_w_bits_strb; // @[LazyModule.scala 167:57]
  assign axi4buf_8_auto_in_w_bits_last = bus_auto_out_8_w_bits_last; // @[LazyModule.scala 167:57]
  assign axi4buf_8_auto_in_b_ready = bus_auto_out_8_b_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_8_auto_in_ar_valid = bus_auto_out_8_ar_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_8_auto_in_ar_bits_id = bus_auto_out_8_ar_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_8_auto_in_ar_bits_addr = bus_auto_out_8_ar_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_8_auto_in_ar_bits_size = bus_auto_out_8_ar_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_8_auto_in_r_ready = bus_auto_out_8_r_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_8_auto_out_aw_ready = nco_mux_1_auto_register_in_aw_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_8_auto_out_w_ready = nco_mux_1_auto_register_in_w_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_8_auto_out_b_valid = nco_mux_1_auto_register_in_b_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_8_auto_out_b_bits_id = nco_mux_1_auto_register_in_b_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_8_auto_out_b_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_8_auto_out_ar_ready = nco_mux_1_auto_register_in_ar_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_8_auto_out_r_valid = nco_mux_1_auto_register_in_r_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_8_auto_out_r_bits_id = nco_mux_1_auto_register_in_r_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_8_auto_out_r_bits_data = nco_mux_1_auto_register_in_r_bits_data; // @[LazyModule.scala 167:31]
  assign axi4buf_8_auto_out_r_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_8_auto_out_r_bits_last = 1'h1; // @[LazyModule.scala 167:31]
  assign axi4buf_9_clock = clock;
  assign axi4buf_9_reset = reset;
  assign axi4buf_9_auto_in_aw_valid = bus_auto_out_9_aw_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_9_auto_in_aw_bits_id = bus_auto_out_9_aw_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_9_auto_in_aw_bits_addr = bus_auto_out_9_aw_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_9_auto_in_aw_bits_size = bus_auto_out_9_aw_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_9_auto_in_w_valid = bus_auto_out_9_w_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_9_auto_in_w_bits_data = bus_auto_out_9_w_bits_data; // @[LazyModule.scala 167:57]
  assign axi4buf_9_auto_in_w_bits_strb = bus_auto_out_9_w_bits_strb; // @[LazyModule.scala 167:57]
  assign axi4buf_9_auto_in_w_bits_last = bus_auto_out_9_w_bits_last; // @[LazyModule.scala 167:57]
  assign axi4buf_9_auto_in_b_ready = bus_auto_out_9_b_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_9_auto_in_ar_valid = bus_auto_out_9_ar_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_9_auto_in_ar_bits_id = bus_auto_out_9_ar_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_9_auto_in_ar_bits_addr = bus_auto_out_9_ar_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_9_auto_in_ar_bits_size = bus_auto_out_9_ar_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_9_auto_in_r_ready = bus_auto_out_9_r_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_9_auto_out_aw_ready = fft_auto_mem_in_aw_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_9_auto_out_w_ready = fft_auto_mem_in_w_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_9_auto_out_b_valid = fft_auto_mem_in_b_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_9_auto_out_b_bits_id = fft_auto_mem_in_b_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_9_auto_out_b_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_9_auto_out_ar_ready = fft_auto_mem_in_ar_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_9_auto_out_r_valid = fft_auto_mem_in_r_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_9_auto_out_r_bits_id = fft_auto_mem_in_r_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_9_auto_out_r_bits_data = fft_auto_mem_in_r_bits_data; // @[LazyModule.scala 167:31]
  assign axi4buf_9_auto_out_r_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_9_auto_out_r_bits_last = 1'h1; // @[LazyModule.scala 167:31]
  assign axi4buf_10_clock = clock;
  assign axi4buf_10_reset = reset;
  assign axi4buf_10_auto_in_aw_valid = bus_auto_out_10_aw_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_10_auto_in_aw_bits_id = bus_auto_out_10_aw_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_10_auto_in_aw_bits_addr = bus_auto_out_10_aw_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_10_auto_in_aw_bits_size = bus_auto_out_10_aw_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_10_auto_in_w_valid = bus_auto_out_10_w_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_10_auto_in_w_bits_data = bus_auto_out_10_w_bits_data; // @[LazyModule.scala 167:57]
  assign axi4buf_10_auto_in_w_bits_strb = bus_auto_out_10_w_bits_strb; // @[LazyModule.scala 167:57]
  assign axi4buf_10_auto_in_w_bits_last = bus_auto_out_10_w_bits_last; // @[LazyModule.scala 167:57]
  assign axi4buf_10_auto_in_b_ready = bus_auto_out_10_b_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_10_auto_in_ar_valid = bus_auto_out_10_ar_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_10_auto_in_ar_bits_id = bus_auto_out_10_ar_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_10_auto_in_ar_bits_addr = bus_auto_out_10_ar_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_10_auto_in_ar_bits_size = bus_auto_out_10_ar_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_10_auto_in_r_ready = bus_auto_out_10_r_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_10_auto_out_aw_ready = fft_split_auto_mem_in_aw_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_10_auto_out_w_ready = fft_split_auto_mem_in_w_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_10_auto_out_b_valid = fft_split_auto_mem_in_b_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_10_auto_out_b_bits_id = fft_split_auto_mem_in_b_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_10_auto_out_b_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_10_auto_out_ar_ready = fft_split_auto_mem_in_ar_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_10_auto_out_r_valid = fft_split_auto_mem_in_r_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_10_auto_out_r_bits_id = fft_split_auto_mem_in_r_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_10_auto_out_r_bits_data = fft_split_auto_mem_in_r_bits_data; // @[LazyModule.scala 167:31]
  assign axi4buf_10_auto_out_r_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_10_auto_out_r_bits_last = 1'h1; // @[LazyModule.scala 167:31]
  assign axi4buf_11_clock = clock;
  assign axi4buf_11_reset = reset;
  assign axi4buf_11_auto_in_aw_valid = bus_auto_out_11_aw_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_11_auto_in_aw_bits_id = bus_auto_out_11_aw_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_11_auto_in_aw_bits_addr = bus_auto_out_11_aw_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_11_auto_in_aw_bits_size = bus_auto_out_11_aw_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_11_auto_in_w_valid = bus_auto_out_11_w_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_11_auto_in_w_bits_data = bus_auto_out_11_w_bits_data; // @[LazyModule.scala 167:57]
  assign axi4buf_11_auto_in_w_bits_strb = bus_auto_out_11_w_bits_strb; // @[LazyModule.scala 167:57]
  assign axi4buf_11_auto_in_w_bits_last = bus_auto_out_11_w_bits_last; // @[LazyModule.scala 167:57]
  assign axi4buf_11_auto_in_b_ready = bus_auto_out_11_b_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_11_auto_in_ar_valid = bus_auto_out_11_ar_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_11_auto_in_ar_bits_id = bus_auto_out_11_ar_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_11_auto_in_ar_bits_addr = bus_auto_out_11_ar_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_11_auto_in_ar_bits_size = bus_auto_out_11_ar_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_11_auto_in_r_ready = bus_auto_out_11_r_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_11_auto_out_aw_ready = fft_mux_0_auto_register_in_aw_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_11_auto_out_w_ready = fft_mux_0_auto_register_in_w_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_11_auto_out_b_valid = fft_mux_0_auto_register_in_b_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_11_auto_out_b_bits_id = fft_mux_0_auto_register_in_b_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_11_auto_out_b_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_11_auto_out_ar_ready = fft_mux_0_auto_register_in_ar_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_11_auto_out_r_valid = fft_mux_0_auto_register_in_r_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_11_auto_out_r_bits_id = fft_mux_0_auto_register_in_r_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_11_auto_out_r_bits_data = fft_mux_0_auto_register_in_r_bits_data; // @[LazyModule.scala 167:31]
  assign axi4buf_11_auto_out_r_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_11_auto_out_r_bits_last = 1'h1; // @[LazyModule.scala 167:31]
  assign axi4buf_12_clock = clock;
  assign axi4buf_12_reset = reset;
  assign axi4buf_12_auto_in_aw_valid = bus_auto_out_12_aw_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_12_auto_in_aw_bits_id = bus_auto_out_12_aw_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_12_auto_in_aw_bits_addr = bus_auto_out_12_aw_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_12_auto_in_aw_bits_size = bus_auto_out_12_aw_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_12_auto_in_w_valid = bus_auto_out_12_w_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_12_auto_in_w_bits_data = bus_auto_out_12_w_bits_data; // @[LazyModule.scala 167:57]
  assign axi4buf_12_auto_in_w_bits_strb = bus_auto_out_12_w_bits_strb; // @[LazyModule.scala 167:57]
  assign axi4buf_12_auto_in_w_bits_last = bus_auto_out_12_w_bits_last; // @[LazyModule.scala 167:57]
  assign axi4buf_12_auto_in_b_ready = bus_auto_out_12_b_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_12_auto_in_ar_valid = bus_auto_out_12_ar_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_12_auto_in_ar_bits_id = bus_auto_out_12_ar_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_12_auto_in_ar_bits_addr = bus_auto_out_12_ar_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_12_auto_in_ar_bits_size = bus_auto_out_12_ar_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_12_auto_in_r_ready = bus_auto_out_12_r_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_12_auto_out_aw_ready = fft_mux_1_auto_register_in_aw_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_12_auto_out_w_ready = fft_mux_1_auto_register_in_w_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_12_auto_out_b_valid = fft_mux_1_auto_register_in_b_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_12_auto_out_b_bits_id = fft_mux_1_auto_register_in_b_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_12_auto_out_b_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_12_auto_out_ar_ready = fft_mux_1_auto_register_in_ar_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_12_auto_out_r_valid = fft_mux_1_auto_register_in_r_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_12_auto_out_r_bits_id = fft_mux_1_auto_register_in_r_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_12_auto_out_r_bits_data = fft_mux_1_auto_register_in_r_bits_data; // @[LazyModule.scala 167:31]
  assign axi4buf_12_auto_out_r_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_12_auto_out_r_bits_last = 1'h1; // @[LazyModule.scala 167:31]
  assign axi4buf_13_clock = clock;
  assign axi4buf_13_reset = reset;
  assign axi4buf_13_auto_in_aw_valid = bus_auto_out_13_aw_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_13_auto_in_aw_bits_id = bus_auto_out_13_aw_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_13_auto_in_aw_bits_addr = bus_auto_out_13_aw_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_13_auto_in_aw_bits_size = bus_auto_out_13_aw_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_13_auto_in_w_valid = bus_auto_out_13_w_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_13_auto_in_w_bits_data = bus_auto_out_13_w_bits_data; // @[LazyModule.scala 167:57]
  assign axi4buf_13_auto_in_w_bits_strb = bus_auto_out_13_w_bits_strb; // @[LazyModule.scala 167:57]
  assign axi4buf_13_auto_in_w_bits_last = bus_auto_out_13_w_bits_last; // @[LazyModule.scala 167:57]
  assign axi4buf_13_auto_in_b_ready = bus_auto_out_13_b_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_13_auto_in_ar_valid = bus_auto_out_13_ar_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_13_auto_in_ar_bits_id = bus_auto_out_13_ar_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_13_auto_in_ar_bits_addr = bus_auto_out_13_ar_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_13_auto_in_ar_bits_size = bus_auto_out_13_ar_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_13_auto_in_r_ready = bus_auto_out_13_r_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_13_auto_out_aw_ready = mag_auto_mem_in_aw_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_13_auto_out_w_ready = mag_auto_mem_in_w_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_13_auto_out_b_valid = mag_auto_mem_in_b_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_13_auto_out_b_bits_id = mag_auto_mem_in_b_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_13_auto_out_b_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_13_auto_out_ar_ready = mag_auto_mem_in_ar_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_13_auto_out_r_valid = mag_auto_mem_in_r_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_13_auto_out_r_bits_id = mag_auto_mem_in_r_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_13_auto_out_r_bits_data = mag_auto_mem_in_r_bits_data; // @[LazyModule.scala 167:31]
  assign axi4buf_13_auto_out_r_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_13_auto_out_r_bits_last = 1'h1; // @[LazyModule.scala 167:31]
  assign axi4buf_14_clock = clock;
  assign axi4buf_14_reset = reset;
  assign axi4buf_14_auto_in_aw_valid = bus_auto_out_14_aw_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_14_auto_in_aw_bits_id = bus_auto_out_14_aw_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_14_auto_in_aw_bits_addr = bus_auto_out_14_aw_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_14_auto_in_aw_bits_size = bus_auto_out_14_aw_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_14_auto_in_w_valid = bus_auto_out_14_w_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_14_auto_in_w_bits_data = bus_auto_out_14_w_bits_data; // @[LazyModule.scala 167:57]
  assign axi4buf_14_auto_in_w_bits_strb = bus_auto_out_14_w_bits_strb; // @[LazyModule.scala 167:57]
  assign axi4buf_14_auto_in_w_bits_last = bus_auto_out_14_w_bits_last; // @[LazyModule.scala 167:57]
  assign axi4buf_14_auto_in_b_ready = bus_auto_out_14_b_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_14_auto_in_ar_valid = bus_auto_out_14_ar_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_14_auto_in_ar_bits_id = bus_auto_out_14_ar_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_14_auto_in_ar_bits_addr = bus_auto_out_14_ar_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_14_auto_in_ar_bits_size = bus_auto_out_14_ar_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_14_auto_in_r_ready = bus_auto_out_14_r_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_14_auto_out_aw_ready = mag_split_auto_mem_in_aw_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_14_auto_out_w_ready = mag_split_auto_mem_in_w_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_14_auto_out_b_valid = mag_split_auto_mem_in_b_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_14_auto_out_b_bits_id = mag_split_auto_mem_in_b_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_14_auto_out_b_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_14_auto_out_ar_ready = mag_split_auto_mem_in_ar_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_14_auto_out_r_valid = mag_split_auto_mem_in_r_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_14_auto_out_r_bits_id = mag_split_auto_mem_in_r_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_14_auto_out_r_bits_data = mag_split_auto_mem_in_r_bits_data; // @[LazyModule.scala 167:31]
  assign axi4buf_14_auto_out_r_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_14_auto_out_r_bits_last = 1'h1; // @[LazyModule.scala 167:31]
  assign axi4buf_15_clock = clock;
  assign axi4buf_15_reset = reset;
  assign axi4buf_15_auto_in_aw_valid = bus_auto_out_15_aw_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_15_auto_in_aw_bits_id = bus_auto_out_15_aw_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_15_auto_in_aw_bits_addr = bus_auto_out_15_aw_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_15_auto_in_aw_bits_size = bus_auto_out_15_aw_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_15_auto_in_w_valid = bus_auto_out_15_w_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_15_auto_in_w_bits_data = bus_auto_out_15_w_bits_data; // @[LazyModule.scala 167:57]
  assign axi4buf_15_auto_in_w_bits_strb = bus_auto_out_15_w_bits_strb; // @[LazyModule.scala 167:57]
  assign axi4buf_15_auto_in_w_bits_last = bus_auto_out_15_w_bits_last; // @[LazyModule.scala 167:57]
  assign axi4buf_15_auto_in_b_ready = bus_auto_out_15_b_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_15_auto_in_ar_valid = bus_auto_out_15_ar_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_15_auto_in_ar_bits_id = bus_auto_out_15_ar_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_15_auto_in_ar_bits_addr = bus_auto_out_15_ar_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_15_auto_in_ar_bits_size = bus_auto_out_15_ar_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_15_auto_in_r_ready = bus_auto_out_15_r_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_15_auto_out_aw_ready = mag_mux_0_auto_register_in_aw_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_15_auto_out_w_ready = mag_mux_0_auto_register_in_w_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_15_auto_out_b_valid = mag_mux_0_auto_register_in_b_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_15_auto_out_b_bits_id = mag_mux_0_auto_register_in_b_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_15_auto_out_b_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_15_auto_out_ar_ready = mag_mux_0_auto_register_in_ar_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_15_auto_out_r_valid = mag_mux_0_auto_register_in_r_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_15_auto_out_r_bits_id = mag_mux_0_auto_register_in_r_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_15_auto_out_r_bits_data = mag_mux_0_auto_register_in_r_bits_data; // @[LazyModule.scala 167:31]
  assign axi4buf_15_auto_out_r_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_15_auto_out_r_bits_last = 1'h1; // @[LazyModule.scala 167:31]
  assign axi4buf_16_clock = clock;
  assign axi4buf_16_reset = reset;
  assign axi4buf_16_auto_in_aw_valid = bus_auto_out_16_aw_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_16_auto_in_aw_bits_id = bus_auto_out_16_aw_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_16_auto_in_aw_bits_addr = bus_auto_out_16_aw_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_16_auto_in_aw_bits_size = bus_auto_out_16_aw_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_16_auto_in_w_valid = bus_auto_out_16_w_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_16_auto_in_w_bits_data = bus_auto_out_16_w_bits_data; // @[LazyModule.scala 167:57]
  assign axi4buf_16_auto_in_w_bits_strb = bus_auto_out_16_w_bits_strb; // @[LazyModule.scala 167:57]
  assign axi4buf_16_auto_in_w_bits_last = bus_auto_out_16_w_bits_last; // @[LazyModule.scala 167:57]
  assign axi4buf_16_auto_in_b_ready = bus_auto_out_16_b_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_16_auto_in_ar_valid = bus_auto_out_16_ar_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_16_auto_in_ar_bits_id = bus_auto_out_16_ar_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_16_auto_in_ar_bits_addr = bus_auto_out_16_ar_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_16_auto_in_ar_bits_size = bus_auto_out_16_ar_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_16_auto_in_r_ready = bus_auto_out_16_r_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_16_auto_out_aw_ready = mag_mux_1_auto_register_in_aw_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_16_auto_out_w_ready = mag_mux_1_auto_register_in_w_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_16_auto_out_b_valid = mag_mux_1_auto_register_in_b_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_16_auto_out_b_bits_id = mag_mux_1_auto_register_in_b_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_16_auto_out_b_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_16_auto_out_ar_ready = mag_mux_1_auto_register_in_ar_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_16_auto_out_r_valid = mag_mux_1_auto_register_in_r_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_16_auto_out_r_bits_id = mag_mux_1_auto_register_in_r_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_16_auto_out_r_bits_data = mag_mux_1_auto_register_in_r_bits_data; // @[LazyModule.scala 167:31]
  assign axi4buf_16_auto_out_r_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_16_auto_out_r_bits_last = 1'h1; // @[LazyModule.scala 167:31]
  assign axi4buf_17_clock = clock;
  assign axi4buf_17_reset = reset;
  assign axi4buf_17_auto_in_aw_valid = bus_auto_out_17_aw_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_17_auto_in_aw_bits_id = bus_auto_out_17_aw_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_17_auto_in_aw_bits_addr = bus_auto_out_17_aw_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_17_auto_in_aw_bits_size = bus_auto_out_17_aw_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_17_auto_in_w_valid = bus_auto_out_17_w_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_17_auto_in_w_bits_data = bus_auto_out_17_w_bits_data; // @[LazyModule.scala 167:57]
  assign axi4buf_17_auto_in_w_bits_strb = bus_auto_out_17_w_bits_strb; // @[LazyModule.scala 167:57]
  assign axi4buf_17_auto_in_w_bits_last = bus_auto_out_17_w_bits_last; // @[LazyModule.scala 167:57]
  assign axi4buf_17_auto_in_b_ready = bus_auto_out_17_b_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_17_auto_in_ar_valid = bus_auto_out_17_ar_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_17_auto_in_ar_bits_id = bus_auto_out_17_ar_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_17_auto_in_ar_bits_addr = bus_auto_out_17_ar_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_17_auto_in_ar_bits_size = bus_auto_out_17_ar_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_17_auto_in_r_ready = bus_auto_out_17_r_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_17_auto_out_aw_ready = out_mux_auto_register_in_aw_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_17_auto_out_w_ready = out_mux_auto_register_in_w_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_17_auto_out_b_valid = out_mux_auto_register_in_b_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_17_auto_out_b_bits_id = out_mux_auto_register_in_b_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_17_auto_out_b_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_17_auto_out_ar_ready = out_mux_auto_register_in_ar_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_17_auto_out_r_valid = out_mux_auto_register_in_r_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_17_auto_out_r_bits_id = out_mux_auto_register_in_r_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_17_auto_out_r_bits_data = out_mux_auto_register_in_r_bits_data; // @[LazyModule.scala 167:31]
  assign axi4buf_17_auto_out_r_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_17_auto_out_r_bits_last = 1'h1; // @[LazyModule.scala 167:31]
  assign axi4buf_18_clock = clock;
  assign axi4buf_18_reset = reset;
  assign axi4buf_18_auto_in_aw_valid = bus_auto_out_18_aw_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_18_auto_in_aw_bits_id = bus_auto_out_18_aw_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_18_auto_in_aw_bits_addr = bus_auto_out_18_aw_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_18_auto_in_aw_bits_size = bus_auto_out_18_aw_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_18_auto_in_w_valid = bus_auto_out_18_w_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_18_auto_in_w_bits_data = bus_auto_out_18_w_bits_data; // @[LazyModule.scala 167:57]
  assign axi4buf_18_auto_in_w_bits_strb = bus_auto_out_18_w_bits_strb; // @[LazyModule.scala 167:57]
  assign axi4buf_18_auto_in_w_bits_last = bus_auto_out_18_w_bits_last; // @[LazyModule.scala 167:57]
  assign axi4buf_18_auto_in_b_ready = bus_auto_out_18_b_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_18_auto_in_ar_valid = bus_auto_out_18_ar_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_18_auto_in_ar_bits_id = bus_auto_out_18_ar_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_18_auto_in_ar_bits_addr = bus_auto_out_18_ar_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_18_auto_in_ar_bits_size = bus_auto_out_18_ar_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_18_auto_in_r_ready = bus_auto_out_18_r_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_18_auto_out_aw_ready = uart_auto_mem_in_aw_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_18_auto_out_w_ready = uart_auto_mem_in_w_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_18_auto_out_b_valid = uart_auto_mem_in_b_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_18_auto_out_b_bits_id = uart_auto_mem_in_b_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_18_auto_out_b_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_18_auto_out_ar_ready = uart_auto_mem_in_ar_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_18_auto_out_r_valid = uart_auto_mem_in_r_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_18_auto_out_r_bits_id = uart_auto_mem_in_r_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_18_auto_out_r_bits_data = uart_auto_mem_in_r_bits_data; // @[LazyModule.scala 167:31]
  assign axi4buf_18_auto_out_r_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_18_auto_out_r_bits_last = 1'h1; // @[LazyModule.scala 167:31]
  assign axi4buf_19_clock = clock;
  assign axi4buf_19_reset = reset;
  assign axi4buf_19_auto_in_aw_valid = bus_auto_out_19_aw_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_19_auto_in_aw_bits_id = bus_auto_out_19_aw_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_19_auto_in_aw_bits_addr = bus_auto_out_19_aw_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_19_auto_in_aw_bits_size = bus_auto_out_19_aw_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_19_auto_in_w_valid = bus_auto_out_19_w_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_19_auto_in_w_bits_data = bus_auto_out_19_w_bits_data; // @[LazyModule.scala 167:57]
  assign axi4buf_19_auto_in_w_bits_strb = bus_auto_out_19_w_bits_strb; // @[LazyModule.scala 167:57]
  assign axi4buf_19_auto_in_w_bits_last = bus_auto_out_19_w_bits_last; // @[LazyModule.scala 167:57]
  assign axi4buf_19_auto_in_b_ready = bus_auto_out_19_b_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_19_auto_in_ar_valid = bus_auto_out_19_ar_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_19_auto_in_ar_bits_id = bus_auto_out_19_ar_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_19_auto_in_ar_bits_addr = bus_auto_out_19_ar_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_19_auto_in_ar_bits_size = bus_auto_out_19_ar_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_19_auto_in_r_ready = bus_auto_out_19_r_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_19_auto_out_aw_ready = uRx_split_auto_mem_in_aw_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_19_auto_out_w_ready = uRx_split_auto_mem_in_w_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_19_auto_out_b_valid = uRx_split_auto_mem_in_b_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_19_auto_out_b_bits_id = uRx_split_auto_mem_in_b_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_19_auto_out_b_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_19_auto_out_ar_ready = uRx_split_auto_mem_in_ar_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_19_auto_out_r_valid = uRx_split_auto_mem_in_r_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_19_auto_out_r_bits_id = uRx_split_auto_mem_in_r_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_19_auto_out_r_bits_data = uRx_split_auto_mem_in_r_bits_data; // @[LazyModule.scala 167:31]
  assign axi4buf_19_auto_out_r_bits_resp = 2'h0; // @[LazyModule.scala 167:31]
  assign axi4buf_19_auto_out_r_bits_last = 1'h1; // @[LazyModule.scala 167:31]
  assign buffer_clock = clock;
  assign buffer_reset = reset;
  assign buffer_auto_in_valid = nco_mux_0_auto_stream_out_0_valid; // @[LazyModule.scala 167:57]
  assign buffer_auto_in_bits_data = nco_mux_0_auto_stream_out_0_bits_data; // @[LazyModule.scala 167:57]
  assign buffer_auto_in_bits_last = nco_mux_0_auto_stream_out_0_bits_last; // @[LazyModule.scala 167:57]
  assign buffer_auto_out_ready = fft_auto_stream_in_ready; // @[LazyModule.scala 167:31]
  assign buffer_1_clock = clock;
  assign buffer_1_reset = reset;
  assign buffer_1_auto_in_valid = fft_mux_0_auto_stream_out_0_valid; // @[LazyModule.scala 167:57]
  assign buffer_1_auto_in_bits_data = fft_mux_0_auto_stream_out_0_bits_data; // @[LazyModule.scala 167:57]
  assign buffer_1_auto_in_bits_last = fft_mux_0_auto_stream_out_0_bits_last; // @[LazyModule.scala 167:57]
  assign buffer_1_auto_out_ready = mag_auto_stream_in_ready; // @[LazyModule.scala 167:31]
  assign buffer_2_clock = clock;
  assign buffer_2_reset = reset;
  assign buffer_2_auto_in_valid = mag_mux_0_auto_stream_out_0_valid; // @[LazyModule.scala 167:57]
  assign buffer_2_auto_in_bits_data = mag_mux_0_auto_stream_out_0_bits_data; // @[LazyModule.scala 167:57]
  assign buffer_2_auto_in_bits_last = mag_mux_0_auto_stream_out_0_bits_last; // @[LazyModule.scala 167:57]
  assign buffer_2_auto_out_ready = acc_auto_accumulator_slave_in_ready; // @[LazyModule.scala 167:31]
  assign buffer_3_clock = clock;
  assign buffer_3_reset = reset;
  assign buffer_3_auto_in_valid = mag_mux_1_auto_stream_out_1_valid; // @[LazyModule.scala 167:57]
  assign buffer_3_auto_in_bits_data = mag_mux_1_auto_stream_out_1_bits_data; // @[LazyModule.scala 167:57]
  assign buffer_3_auto_in_bits_last = mag_mux_1_auto_stream_out_1_bits_last; // @[LazyModule.scala 167:57]
  assign buffer_3_auto_out_ready = out_mux_auto_stream_in_1_ready; // @[LazyModule.scala 167:31]
  assign buffer_4_clock = clock;
  assign buffer_4_reset = reset;
  assign buffer_4_auto_in_valid = fft_mux_1_auto_stream_out_1_valid; // @[LazyModule.scala 167:57]
  assign buffer_4_auto_in_bits_data = fft_mux_1_auto_stream_out_1_bits_data; // @[LazyModule.scala 167:57]
  assign buffer_4_auto_in_bits_last = fft_mux_1_auto_stream_out_1_bits_last; // @[LazyModule.scala 167:57]
  assign buffer_4_auto_out_ready = out_mux_auto_stream_in_2_ready; // @[LazyModule.scala 167:31]
  assign buffer_5_clock = clock;
  assign buffer_5_reset = reset;
  assign buffer_5_auto_in_valid = nco_mux_1_auto_stream_out_1_valid; // @[LazyModule.scala 167:57]
  assign buffer_5_auto_in_bits_data = nco_mux_1_auto_stream_out_1_bits_data; // @[LazyModule.scala 167:57]
  assign buffer_5_auto_in_bits_last = nco_mux_1_auto_stream_out_1_bits_last; // @[LazyModule.scala 167:57]
  assign buffer_5_auto_out_ready = out_mux_auto_stream_in_3_ready; // @[LazyModule.scala 167:31]
  assign buffer_6_clock = clock;
  assign buffer_6_reset = reset;
  assign buffer_6_auto_in_valid = plfg_mux_1_auto_stream_out_1_valid; // @[LazyModule.scala 167:57]
  assign buffer_6_auto_in_bits_data = plfg_mux_1_auto_stream_out_1_bits_data; // @[LazyModule.scala 167:57]
  assign buffer_6_auto_in_bits_last = plfg_mux_1_auto_stream_out_1_bits_last; // @[LazyModule.scala 167:57]
  assign buffer_6_auto_out_ready = out_mux_auto_stream_in_4_ready; // @[LazyModule.scala 167:31]
  assign buffer_7_clock = clock;
  assign buffer_7_reset = reset;
  assign buffer_7_auto_in_valid = in_split_auto_stream_out_4_valid; // @[LazyModule.scala 167:57]
  assign buffer_7_auto_in_bits_data = in_split_auto_stream_out_4_bits_data; // @[LazyModule.scala 167:57]
  assign buffer_7_auto_in_bits_last = in_split_auto_stream_out_4_bits_last; // @[LazyModule.scala 167:57]
  assign buffer_7_auto_out_ready = out_mux_auto_stream_in_5_ready; // @[LazyModule.scala 167:31]
  assign buffer_8_clock = clock;
  assign buffer_8_reset = reset;
  assign buffer_8_auto_in_valid = uRx_split_auto_stream_out_4_valid; // @[LazyModule.scala 167:57]
  assign buffer_8_auto_in_bits_data = uRx_split_auto_stream_out_4_bits_data; // @[LazyModule.scala 167:57]
  assign buffer_8_auto_in_bits_last = uRx_split_auto_stream_out_4_bits_last; // @[LazyModule.scala 167:57]
  assign buffer_8_auto_out_ready = out_mux_auto_stream_in_6_ready; // @[LazyModule.scala 167:31]
  assign buffer_9_clock = clock;
  assign buffer_9_reset = reset;
  assign buffer_9_auto_in_valid = out_mux_auto_stream_out_0_valid; // @[LazyModule.scala 167:57]
  assign buffer_9_auto_in_bits_data = out_mux_auto_stream_out_0_bits_data; // @[LazyModule.scala 167:57]
  assign buffer_9_auto_in_bits_last = out_mux_auto_stream_out_0_bits_last; // @[LazyModule.scala 167:57]
  assign buffer_9_auto_out_ready = out_queue_auto_in_in_ready; // @[LazyModule.scala 167:31]
  assign converter_auto_in_aw_valid = ioMem_0_aw_valid; // @[LazyModule.scala 167:57]
  assign converter_auto_in_aw_bits_id = ioMem_0_aw_bits_id; // @[LazyModule.scala 167:57]
  assign converter_auto_in_aw_bits_addr = ioMem_0_aw_bits_addr; // @[LazyModule.scala 167:57]
  assign converter_auto_in_aw_bits_size = ioMem_0_aw_bits_size; // @[LazyModule.scala 167:57]
  assign converter_auto_in_w_valid = ioMem_0_w_valid; // @[LazyModule.scala 167:57]
  assign converter_auto_in_w_bits_data = ioMem_0_w_bits_data; // @[LazyModule.scala 167:57]
  assign converter_auto_in_w_bits_strb = ioMem_0_w_bits_strb; // @[LazyModule.scala 167:57]
  assign converter_auto_in_w_bits_last = ioMem_0_w_bits_last; // @[LazyModule.scala 167:57]
  assign converter_auto_in_b_ready = ioMem_0_b_ready; // @[LazyModule.scala 167:57]
  assign converter_auto_in_ar_valid = ioMem_0_ar_valid; // @[LazyModule.scala 167:57]
  assign converter_auto_in_ar_bits_id = ioMem_0_ar_bits_id; // @[LazyModule.scala 167:57]
  assign converter_auto_in_ar_bits_addr = ioMem_0_ar_bits_addr; // @[LazyModule.scala 167:57]
  assign converter_auto_in_ar_bits_size = ioMem_0_ar_bits_size; // @[LazyModule.scala 167:57]
  assign converter_auto_in_r_ready = ioMem_0_r_ready; // @[LazyModule.scala 167:57]
  assign converter_auto_out_aw_ready = bus_auto_in_aw_ready; // @[LazyModule.scala 167:31]
  assign converter_auto_out_w_ready = bus_auto_in_w_ready; // @[LazyModule.scala 167:31]
  assign converter_auto_out_b_valid = bus_auto_in_b_valid; // @[LazyModule.scala 167:31]
  assign converter_auto_out_b_bits_resp = bus_auto_in_b_bits_resp; // @[LazyModule.scala 167:31]
  assign converter_auto_out_ar_ready = bus_auto_in_ar_ready; // @[LazyModule.scala 167:31]
  assign converter_auto_out_r_valid = bus_auto_in_r_valid; // @[LazyModule.scala 167:31]
  assign converter_auto_out_r_bits_data = bus_auto_in_r_bits_data; // @[LazyModule.scala 167:31]
  assign converter_auto_out_r_bits_resp = bus_auto_in_r_bits_resp; // @[LazyModule.scala 167:31]
  assign converter_auto_out_r_bits_last = bus_auto_in_r_bits_last; // @[LazyModule.scala 167:31]
  assign converter_1_auto_in_valid = widthAdapter_2_auto_out_valid; // @[LazyModule.scala 167:57]
  assign converter_1_auto_in_bits_data = widthAdapter_2_auto_out_bits_data; // @[LazyModule.scala 167:57]
  assign converter_1_auto_in_bits_last = widthAdapter_2_auto_out_bits_last; // @[LazyModule.scala 167:57]
  assign converter_1_auto_out_ready = outStream_0_ready; // @[LazyModule.scala 167:31]
  assign converter_2_auto_in_valid = inStream_0_valid; // @[LazyModule.scala 167:57]
  assign converter_2_auto_in_bits_data = inStream_0_bits_data; // @[LazyModule.scala 167:57]
  assign converter_2_auto_in_bits_last = inStream_0_bits_last; // @[LazyModule.scala 167:57]
  assign converter_2_auto_out_ready = in_queue_auto_in_in_ready; // @[LazyModule.scala 167:31]
endmodule
